* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre=0.0
* statistics {
*   process {
*   }
*   mismatch {
*     vary sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre dist=gauss std = 1.0
*   }
* }
.subckt sky130_fd_pr__pfet_g5v0d10v5 d g s b
.param l=1 w=1 ad=0 as=0 pd=0 ps=0 nrd=0 nrs=0 sa=0 sb=0 sd=0 mult=1 nf=1.0
msky130_fd_pr__pfet_g5v0d10v5 d g s b sky130_fd_pr__pfet_g5v0d10v5__model l={l} w={w} ad={ad} as={as} pd={pd} ps={ps} nrd={nrd} nrs={nrs} sa={sa} sb={sb} sd={sd} nf={nf}
.model sky130_fd_pr__pfet_g5v0d10v5__model.0 pmos
* DC IV MOS Parameters
+  lmin=2.0e-05 lmax=1.0e-04 wmin=2.0e-05 wmax=1.0e-4
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.057134+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+  k1=0.59521
+  k2=0.0294389
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=200000.0
+  ua=2.7344678e-9
+  ub=-4.4406e-19
+  uc=-3.9972e-11
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0207994
+  a0=0.911307
+  keta=-0.0079259
+  a1=0.0
+  a2=0.5
+  ags=0.1271299
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.093204657+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.69967+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.08353125
+  pdiblc1=0.39
+  pdiblc2=0.0029407877
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=333712830.0
+  pscbe2=1.5000958e-8
+  pvag=0.0
+  delta=0.01
+  alpha0=5.0667189e-5
+  alpha1=0.0
+  beta0=38.266046
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=7.3657e-9
+  bgidl=1704700000.0
+  cgidl=700.0
+  egidl=0.69350825
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.57573
+  kt2=-0.019032
+  at=430000.0
+  ute=-1.3864
+  ua1=7.0656e-10
+  ub1=-3.145e-18
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.1 pmos
* DC IV MOS Parameters
+  lmin=8e-06 lmax=2.0e-05 wmin=2.0e-05 wmax=1.0e-4
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.057134+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+  k1=0.59521
+  k2=0.0294389
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=200000.0
+  ua=2.7344678e-9
+  ub=-4.4406e-19
+  uc=-3.9972e-11
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0207994
+  a0=0.911307
+  keta=-0.0079259
+  a1=0.0
+  a2=0.5
+  ags=0.1271299
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.093204657+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.69967+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.08353125
+  pdiblc1=0.39
+  pdiblc2=0.0029407877
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=333712830.0
+  pscbe2=1.5000958e-8
+  pvag=0.0
+  delta=0.01
+  alpha0=5.0667189e-5
+  alpha1=0.0
+  beta0=38.266046
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=7.3657e-9
+  bgidl=1704700000.0
+  cgidl=700.0
+  egidl=0.69350825
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.57573
+  kt2=-0.019032
+  at=430000.0
+  ute=-1.3864
+  ua1=7.0656e-10
+  ub1=-3.145e-18
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.2 pmos
* DC IV MOS Parameters
+  lmin=4e-06 lmax=8e-06 wmin=2.0e-05 wmax=1.0e-4
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.06129678645+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=3.30687592801532e-8
+  k1=0.60423167125 lk1=-7.16672542428745e-8
+  k2=0.0278592694525 lk2=1.25484271062852e-8
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=298587.64025 lvsat=-0.783170355381975
+  ua=2.4949572179375e-09 lua=1.90264811284629e-15
+  ub=-2.008594065e-19 lub=-1.93196119470465e-24
+  uc=-5.1678481175e-11 luc=9.29951158060825e-17
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0199748291075 lu0=6.55030871293077e-9
+  a0=0.933098033475 la0=-1.73105790822051e-7
+  keta=-0.0049304093525 lketa=-2.37958781546752e-8
+  a1=0.0
+  a2=0.5
+  ags=0.104081156815 lags=1.83096910987322e-7
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.09479041045225+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=1.25970668493288e-8
+  nfactor={1.7321085775+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-2.57688815802249e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-0.6548060915245 lpclm=5.86527800733647e-06 wpclm=-1.6940658945086e-21 ppclm=-3.23117426778526e-27
+  pdiblc1=0.39
+  pdiblc2=0.0045684231025075 lpdiblc2=-1.29297728739793e-8
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=564147837.55925 lpscbe1=-1830.55265654993
+  pscbe2=-1.558611817795e-08 lpscbe2=2.42980674450017e-13
+  pvag=0.0
+  delta=0.01
+  alpha0=7.83968484975e-05 lalpha0=-2.2028164208219e-10
+  alpha1=0.0
+  beta0=39.148037118575 lbeta0=-7.00644924684799e-6
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=6.5314665525e-09 lagidl=6.62706708359525e-15
+  bgidl=1476348190.0 lbgidl=1814.003943459
+  cgidl=934.66205 lcgidl=-0.001864131858995
+  egidl=1.21389074000325 legidl=-4.13386646233682e-6
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.58532353675 lkt1=7.62100965883249e-8
+  kt2=-0.019032
+  at=675202.12275 lat=-1.94786114291372
+  ute=-1.2190800425 lute=-1.32917301038425e-6
+  ua1=1.3814243924e-09 lua1=-5.36105524678636e-15
+  ub1=-2.605671675e-18 lub1=-4.2843702809675e-24
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.3 pmos
* DC IV MOS Parameters
+  lmin=2e-06 lmax=4e-06 wmin=2.0e-05 wmax=1.0e-4
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.0381655746+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-5.81584271350592e-8
+  k1=0.602894174 lk1=-6.63922988386e-8
+  k2=0.0297949601 lk2=4.91425676161001e-9
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=84264.41 lvsat=0.062099032401
+  ua=3.28797678225e-09 lua=-1.22494174684578e-15
+  ub=-1.7328156315e-18 lub=4.10992096107285e-24 wub=-5.87747175411144e-39 pub=-1.12103877145985e-44
+  uc=-5.540982305e-11 luc=1.07711155026895e-16
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.02086513804 lu0=3.039019314044e-9
+  a0=0.8222697474 la0=2.63989886629141e-7
+  keta=-0.0049806758 lketa=-2.359763231238e-8
+  a1=0.0
+  a2=0.5
+  ags=0.101458501175 lags=1.93440402565918e-7
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.06358776784865+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=-1.10463035315009e-7
+  nfactor={2.07037515335+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.59177836429707e-6
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.01798959 leta0=2.44562855999e-7
+  etab=-0.1233522794 letab=2.1041605472566e-7
+  dsub=0.8193648575 ldsub=-1.02290906149425e-6
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=1.0526929389875 lpclm=-8.68927419099802e-7
+  pdiblc1=0.58503867943 lpdiblc1=-7.69213047803977e-7
+  pdiblc2=-0.0011773222896 lpdiblc2=9.73087237795344e-09 ppdiblc2=2.52435489670724e-29
+  pdiblcb=0.16939 lpdiblcb=-7.66654721e-07 wpdiblcb=-2.11758236813575e-22 ppdiblcb=4.03896783473158e-28
+  drout=0.132342 ldrout=1.6866403862e-6
+  pscbe1=-160819458.431 lpscbe1=1028.64586210602
+  pscbe2=7.662008170125e-08 lpscbe2=-1.2067135725356e-13
+  pvag=0.0
+  delta=0.01
+  alpha0=4.445374715855e-05 lalpha0=-8.64134447115054e-11
+  alpha1=-9.7195e-11 lalpha1=3.833273605e-16
+  beta0=70.77889717255 lbeta0=-0.00013175539821372
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=9.21504679e-09 lagidl=-3.956705015081e-15
+  bgidl=2632410590 lbgidl=-2745.390555901
+  cgidl=455.6337275 lcgidl=2.51079421127497e-5
+  egidl=-1.617101386419 legidl=7.0312833850599e-06 wegidl=1.6940658945086e-21 pegidl=3.23117426778526e-27
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.56697195 lkt1=3.83327360500023e-9
+  kt2=-0.019032
+  at=210964.1945 lat=-0.11695317768855
+  ute=-1.707821395 lute=5.98374009740501e-7
+  ua1=-4.933329728e-10 lua1=2.03280032582592e-15 wua1=7.88860905221012e-31 pua1=-1.50463276905253e-36
+  ub1=-3.720478135e-18 lub1=1.12314916626499e-25
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.4 pmos
* DC IV MOS Parameters
+  lmin=1e-06 lmax=2e-06 wmin=2.0e-05 wmax=1.0e-4
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.0877095688+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=3.81501431903203e-8
+  k1=0.558687465 lk1=1.95411227864998e-8
+  k2=0.0276516389 lk2=9.08065884229002e-9
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=180698.1919 lvsat=-0.12535859623441
+  ua=3.54875561152e-09 lua=-1.73186971306373e-15
+  ub=-5.0176592e-20 lub=8.390389321888e-25
+  uc=5.52615694e-13 luc=-1.0742296475666e-18
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.02533542883 lu0=-5.650778952637e-9
+  a0=1.0672917251 la0=-2.1230833582189e-7
+  keta=0.0466423328 lketa=-1.2394759872992e-07 pketa=1.0097419586829e-28
+  a1=0.0
+  a2=0.5
+  ags=-0.2686976498 lags=9.1298694444622e-7
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.1606776136623+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=7.8269915962145e-8
+  nfactor={0.9875336553+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=5.1315722376233e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.47195e-05 lcit=-9.17423605e-12
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.2795057857601 leta0=-2.63798476939058e-7
+  etab=-0.0293684412 letab=2.772087164868e-8
+  dsub=0.056221661 ldsub=4.605649981821e-7
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.041796294998 lpclm=1.09615456715139e-6
+  pdiblc1=-0.00906932782000003 lpdiblc1=3.85673507489298e-7
+  pdiblc2=0.00602058784087 lpdiblc2=-4.26114512466719e-9
+  pdiblcb=-0.41378 lpdiblcb=3.66969442e-7
+  drout=1.556250265901 ldrout=-1.08129489188495e-6
+  pscbe1=433349461.692 lpscbe1=-126.359101721079
+  pscbe2=1.45323618864e-08 lpscbe2=2.09612945270377e-17
+  pvag=0.0
+  delta=0.01
+  alpha0=-6.40086482779e-05 lalpha0=1.2442660577741e-10 walpha0=-9.59846506427666e-26 palpha0=-4.10095184369112e-32
+  alpha1=1.9439e-10 lalpha1=-1.83484721e-16
+  beta0=-41.5076459075 lbeta0=8.65184128795893e-05 wbeta0=-2.71050543121376e-20 pbeta0=7.75481824268463e-26
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=3.71510944e-09 lagidl=6.734623199584e-15
+  bgidl=841407320.0 lbgidl=736.140700652
+  cgidl=438.411273 lcgidl=5.85866714152999e-5
+  egidl=3.152521570876 legidl=-2.24038668162586e-6
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.49779432 lkt1=-1.30641121352e-7
+  kt2=-0.019032
+  at=265011.9 lat=-0.22201651241 wat=-8.88178419700125e-16 pat=-8.470329472543e-22
+  ute=-1.20470709 lute=-3.79629887749e-7
+  ua1=6.77542262e-10 lua1=-2.432640431018e-16 wua1=-3.15544362088405e-30
+  ub1=-3.52706157e-18 lub1=-2.63667544077e-25
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=2.81e-6
+  sbref=2.81e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.5 pmos
* DC IV MOS Parameters
+  lmin=8.0e-07 lmax=1e-06 wmin=2.0e-05 wmax=1.0e-4
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.1149757415+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=6.38866836018495e-8
+  k1=0.59077167 lk1=-1.07431583129997e-8
+  k2=0.032577991 lk2=4.43067509510002e-9
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=7814.73505000002 lvsat=0.037826098686305
+  ua=-8.493986931e-10 lua=2.41954813506709e-15
+  ub=4.763137255e-18 lub=-3.7042480079945e-24 wub=-1.17549435082229e-38
+  uc=6.40846463e-12 luc=-6.601565458257e-18 puc=-1.17549435082229e-38
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.01791493275 lu0=1.353427297275e-9
+  a0=0.838106172500001 la0=4.01990727724933e-9
+  keta=-0.157135299 lketa=6.83981079261e-8
+  a1=0.0
+  a2=0.5
+  ags=0.614610324 lags=7.92325479764003e-8
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.096109477214+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=1.73240519685945e-8
+  nfactor={1.600506602+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-6.54279406278e-8
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-1.35975e-05 lcit=1.755418025e-11
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=-7.65650575e-05 leta0=9.930399767425e-11
+  etab=0.000791398015 letab=-7.470005863585e-10
+  dsub=1.54597013 ldsub=-9.45608581707e-7
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=2.061904095825 lpclm=-8.10625186049218e-7
+  pdiblc1=0.185912130255 lpdiblc1=2.01630509212305e-7
+  pdiblc2=-0.03533450056535 lpdiblc2=3.47739228219639e-8
+  pdiblcb=-0.025
+  drout=0.33218586617 ldrout=7.40994950211371e-8
+  pscbe1=-74402724.1499999 lpscbe1=352.908186495185
+  pscbe2=1.8463592403e-08 lpscbe2=-3.6897271900917e-15
+  pvag=0.0
+  delta=0.01
+  alpha0=0.000255919397305 lalpha0=-1.7755347644829e-10
+  alpha1=0.0
+  beta0=68.0295673025 lbeta0=-1.68737626693297e-5
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=8.953055e-09 lagidl=1.7905263855e-15
+  bgidl=929473000.000002 lbgidl=653.0155053
+  cgidl=427.87536 lcgidl=6.85315196959999e-5
+  egidl=1.887175135705 legidl=-1.04602618146795e-6
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.60904765 lkt1=-2.56291031649999e-8
+  kt2=-0.019032
+  at=47653.6 lat=-0.01685201304
+  ute=-2.07964845 lute=4.46227261955e-7
+  ua1=-7.33113099999995e-11 lua1=4.65466643509e-16
+  ub1=-4.60795225e-18 lub1=7.56585168775001e-25
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=2.41e-6
+  sbref=2.41e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.6 pmos
* DC IV MOS Parameters
+  lmin=6e-07 lmax=8.0e-07 wmin=2.0e-05 wmax=1.0e-4
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.961308743+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-5.04261965823001e-8
+  k1=0.595611255000001 lk1=-1.43433255945002e-8
+  k2=0.035286917 lk2=2.41550504370001e-9
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=61668.41945 lvsat=-0.00223565713885501
+  ua=-2.2348497994e-09 lua=3.45018521304366e-15
+  ub=2.5967598753e-18 lub=-2.09267987523567e-24 wub=-5.87747175411144e-39 pub=-5.60519385729927e-45
+  uc=3.1396334e-12 luc=-4.16988190626e-18
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.00582160995000001 lu0=1.0349650128195e-8
+  a0=0.945572835 la0=-7.59245429565004e-8
+  keta=0.0210589425 lketa=-6.416058832575e-8
+  a1=0.0
+  a2=0.5
+  ags=-0.717169159999999 lags=1.069943306124e-6
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={0.0170483782754999+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=-6.68540767300445e-8
+  nfactor={2.020420625+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-3.778019823375e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=-0.064270328243 leta0=4.78530444313677e-08 weta0=-8.43724224804088e-23 peta0=-5.99534287967969e-29
+  etab=-0.000791398015 letab=4.304413803585e-10
+  dsub=0.18350229023 ldsub=6.79312442979029e-8
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.170632713425 lpclm=5.96291595318143e-7
+  pdiblc1=0.157259843575 lpdiblc1=2.22944945273558e-7
+  pdiblc2=0.0277574173458 lpdiblc2=-1.21601549121406e-8
+  pdiblcb=-0.025
+  drout=-0.81794092163 ldrout=9.29678812465557e-7
+  pscbe1=434417012.98 lpscbe1=-25.6028159558219
+  pscbe2=1.03443636915e-08 lpscbe2=2.35016704839315e-15
+  pvag=0.0
+  delta=0.01
+  alpha0=-0.0001310877634225 lalpha0=1.10341150416898e-10 walpha0=-2.06795153138257e-25 palpha0=1.97215226305253e-31
+  alpha1=0.0
+  beta0=25.181273087 lbeta0=1.50010833975807e-5
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=2.451938855e-08 lagidl=-9.78926914234501e-15
+  bgidl=2079521950.0 lbgidl=-202.505908605
+  cgidl=1308.655 lcgidl=-0.0005866804545
+  egidl=-0.2962646614 legidl=5.7823468359846e-7
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.71154189 lkt1=5.0616361971e-8
+  kt2=-0.019032
+  at=44036.5 lat=-0.01416125235
+  ute=-1.62257375 lute=1.06209392624999e-7
+  ua1=5.534878e-10 lua1=-8.0921441999993e-19
+  ub1=-4.38417815e-18 lub1=5.90119615785e-25
+  uc1=-2.93321028e-10 luc1=1.369676327292e-16
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=2.02e-6
+  sbref=2.01e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.7 pmos
* DC IV MOS Parameters
+  lmin=5e-07 lmax=6e-07 wmin=2.0e-05 wmax=1.0e-4
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.950578983000001+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-5.62621130463e-8
+  k1=0.4413968 lk1=6.95339164800002e-8
+  k2=0.055242305 lk2=-8.4382304895e-9
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=39884.1215 lvsat=0.00961282251615
+  ua=1.24951991657e-08 lua=-4.56148841907423e-15
+  ub=-1.07262765756e-17 lub=5.15371965040884e-24
+  uc=-1.17777450000001e-12 luc=-1.82164374945e-18
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.04045856741 lu0=-8.489391034299e-9
+  a0=0.12388326 la0=3.70992416886e-7
+  keta=-0.145889365 lketa=2.66425961235e-8
+  a1=0.0
+  a2=0.5
+  ags=1.25
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.12509291583+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=1.0456573133937e-8
+  nfactor={1.486344874+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-8.73181813685997e-8
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=3.2195e-05 lcit=-1.20718605e-11
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=-0.226400016 leta0=1.360353816024e-07 weta0=4.2351647362715e-22 peta0=-2.01948391736579e-28
+  etab=0.0170914817 letab=-9.29605689663e-9
+  dsub=0.43592626954 ldsub=-6.9362158048806e-8
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.9578198815 lpclm=1.6814049460215e-7
+  pdiblc1=1.77958506268 lpdiblc1=-6.59437741397652e-7
+  pdiblc2=0.00805992596100001 lpdiblc2=-1.4466893479479e-9
+  pdiblcb=-0.025
+  drout=0.854662854460001 ldrout=1.9949618650206e-8
+  pscbe1=497007191.6 lpscbe1=-59.6456141072401
+  pscbe2=1.5458070132e-08 lpscbe2=-4.31177884594793e-16
+  pvag=0.0
+  delta=0.01
+  alpha0=-4.0758659736e-05 lalpha0=6.12111509218104e-11
+  alpha1=0.0
+  beta0=44.227233967 lbeta0=4.6419852749487e-6
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-2.61805691e-08 lagidl=1.778643782349e-14
+  bgidl=2118695300.0 lbgidl=-223.812293669999
+  cgidl=-2637.594 lcgidl=0.0015596843766 wcgidl=3.46944695195361e-18 pcgidl=-1.65436122510606e-24
+  egidl=1.2178352726 legidl=-2.4528427050414e-7
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.640674999999999 lkt1=1.20718605e-8
+  kt2=-0.019032
+  at=18000.0
+  ute=-1.6710011 lute=1.3254902829e-7
+  ua1=5.52e-10
+  ub1=-8.3561088e-18 lub1=2.75045269632e-24
+  uc1=-4.1496e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=1.81e-6
+  sbref=1.81e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.8 pmos
* DC IV MOS Parameters
+  lmin=2.0e-05 lmax=1.0e-04 wmin=1.5e-05 wmax=2.0e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.057134+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+  k1=0.59521
+  k2=0.0294389
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=200000.0
+  ua=2.7344678e-9
+  ub=-4.4406e-19
+  uc=-3.9972e-11
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0207994
+  a0=0.911307
+  keta=-0.0079259
+  a1=0.0
+  a2=0.5
+  ags=0.1271299
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.093204657+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.69967+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.08353125
+  pdiblc1=0.39
+  pdiblc2=0.0029407877
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=333712830.0
+  pscbe2=1.5000958e-8
+  pvag=0.0
+  delta=0.01
+  alpha0=5.0667189e-5
+  alpha1=0.0
+  beta0=38.266046
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=7.3657e-9
+  bgidl=1704700000.0
+  cgidl=700.0
+  egidl=0.69350825
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.57573
+  kt2=-0.019032
+  at=430000.0
+  ute=-1.3864
+  ua1=7.0656e-10
+  ub1=-3.145e-18
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.9 pmos
* DC IV MOS Parameters
+  lmin=8e-06 lmax=2.0e-05 wmin=1.5e-05 wmax=2.0e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.057134+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+  k1=0.59521
+  k2=0.0294389
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=200000.0
+  ua=2.7344678e-9
+  ub=-4.4406e-19
+  uc=-3.9972e-11
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0207994
+  a0=0.911307
+  keta=-0.0079259
+  a1=0.0
+  a2=0.5
+  ags=0.1271299
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.093204657+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.69967+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.08353125
+  pdiblc1=0.39
+  pdiblc2=0.0029407877
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=333712830.0
+  pscbe2=1.5000958e-8
+  pvag=0.0
+  delta=0.01
+  alpha0=5.0667189e-5
+  alpha1=0.0
+  beta0=38.266046
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=7.3657e-9
+  bgidl=1704700000.0
+  cgidl=700.0
+  egidl=0.69350825
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.57573
+  kt2=-0.019032
+  at=430000.0
+  ute=-1.3864
+  ua1=7.0656e-10
+  ub1=-3.145e-18
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.10 pmos
* DC IV MOS Parameters
+  lmin=4e-06 lmax=8e-06 wmin=1.5e-05 wmax=2.0e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.06129678645+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=3.30687592801549e-8
+  k1=0.60423167125 lk1=-7.16672542428762e-8
+  k2=0.0278592694525001 lk2=1.25484271062854e-8
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=298587.64025 lvsat=-0.783170355381975
+  ua=2.4949572179375e-09 lua=1.9026481128463e-15
+  ub=-2.00859406500001e-19 lub=-1.93196119470465e-24
+  uc=-5.16784811750001e-11 luc=9.29951158060826e-17
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0199748291075 lu0=6.55030871293071e-9
+  a0=0.933098033475001 la0=-1.73105790822052e-7
+  keta=-0.0049304093525 lketa=-2.37958781546752e-8
+  a1=0.0
+  a2=0.5
+  ags=0.104081156815 lags=1.83096910987321e-7
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.0947904104522501+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=1.25970668493291e-8
+  nfactor={1.7321085775+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-2.57688815802243e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-0.6548060915245 lpclm=5.86527800733648e-06 wpclm=1.6940658945086e-21 ppclm=6.46234853557053e-27
+  pdiblc1=0.39
+  pdiblc2=0.0045684231025075 lpdiblc2=-1.29297728739793e-8
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=564147837.55925 lpscbe1=-1830.55265654993
+  pscbe2=-1.558611817795e-08 lpscbe2=2.42980674450017e-13 ppscbe2=-1.54074395550979e-33
+  pvag=0.0
+  delta=0.01
+  alpha0=7.83968484975e-05 lalpha0=-2.2028164208219e-10
+  alpha1=0.0
+  beta0=39.148037118575 lbeta0=-7.00644924684778e-6
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=6.53146655250001e-09 lagidl=6.6270670835952e-15
+  bgidl=1476348190 lbgidl=1814.003943459
+  cgidl=934.66205 lcgidl=-0.00186413185899499
+  egidl=1.21389074000325 legidl=-4.13386646233682e-6
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.58532353675 lkt1=7.62100965883241e-8
+  kt2=-0.019032
+  at=675202.12275 lat=-1.94786114291372
+  ute=-1.2190800425 lute=-1.32917301038425e-6
+  ua1=1.3814243924e-09 lua1=-5.36105524678636e-15
+  ub1=-2.605671675e-18 lub1=-4.28437028096751e-24
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.11 pmos
* DC IV MOS Parameters
+  lmin=2e-06 lmax=4e-06 wmin=1.5e-05 wmax=2.0e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.0381655746+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-5.81584271350634e-8
+  k1=0.602894174 lk1=-6.63922988386004e-8
+  k2=0.0297949601 lk2=4.91425676161003e-9
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=84264.41 lvsat=0.062099032401
+  ua=3.28797678225e-09 lua=-1.22494174684578e-15
+  ub=-1.7328156315e-18 lub=4.10992096107285e-24 pub=-2.24207754291971e-44
+  uc=-5.540982305e-11 luc=1.07711155026895e-16
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.02086513804 lu0=3.03901931404397e-9
+  a0=0.8222697474 la0=2.63989886629138e-7
+  keta=-0.00498067579999999 lketa=-2.359763231238e-8
+  a1=0.0
+  a2=0.5
+  ags=0.101458501175 lags=1.93440402565917e-7
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.0635877678486498+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=-1.10463035315009e-7
+  nfactor={2.07037515335+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.59177836429707e-6
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.0179895899999999 leta0=2.44562855999e-7
+  etab=-0.1233522794 letab=2.1041605472566e-7
+  dsub=0.8193648575 ldsub=-1.02290906149425e-6
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=1.0526929389875 lpclm=-8.689274190998e-7
+  pdiblc1=0.585038679429999 lpdiblc1=-7.69213047803978e-7
+  pdiblc2=-0.0011773222896 lpdiblc2=9.73087237795343e-9
+  pdiblcb=0.16939 lpdiblcb=-7.66654721e-07 wpdiblcb=8.470329472543e-22 ppdiblcb=8.07793566946316e-28
+  drout=0.132342 ldrout=1.6866403862e-6
+  pscbe1=-160819458.431 lpscbe1=1028.64586210602 ppscbe1=-3.46944695195361e-18
+  pscbe2=7.662008170125e-08 lpscbe2=-1.2067135725356e-13
+  pvag=0.0
+  delta=0.01
+  alpha0=4.445374715855e-05 lalpha0=-8.64134447115054e-11
+  alpha1=-9.7195e-11 lalpha1=3.833273605e-16
+  beta0=70.77889717255 lbeta0=-0.00013175539821372
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=9.21504679e-09 lagidl=-3.956705015081e-15
+  bgidl=2632410590.0 lbgidl=-2745.39055590099
+  cgidl=455.6337275 lcgidl=2.51079421127497e-5
+  egidl=-1.617101386419 legidl=7.0312833850599e-06 pegidl=-1.29246970711411e-26
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.56697195 lkt1=3.83327360499981e-9
+  kt2=-0.019032
+  at=210964.1945 lat=-0.11695317768855
+  ute=-1.707821395 lute=5.98374009740499e-7
+  ua1=-4.933329728e-10 lua1=2.03280032582592e-15 wua1=-1.97215226305253e-30 pua1=1.20370621524202e-35
+  ub1=-3.720478135e-18 lub1=1.12314916626508e-25
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.12 pmos
* DC IV MOS Parameters
+  lmin=1e-06 lmax=2e-06 wmin=1.5e-05 wmax=2.0e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.0707046569979+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=5.09429513822171e-09 wvth0=-3.38586431363115e-07 pvth0=6.58178163926759e-13
+  k1=0.558687465 lk1=1.95411227865009e-8
+  k2=0.0276910477338404 lk2=9.00405201018782e-09 wk2=-7.84673073842475e-10 pk2=1.52532598824255e-15
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=180698.1919 lvsat=-0.12535859623441
+  ua=3.53798292529808e-09 lua=-1.71092868831694e-15 wua=2.14495989542561e-16 pua=-4.16958754071732e-22
+  ub=-1.6817586113233e-18 lub=4.01067121955137e-24 wub=3.24865862186201e-23 pub=-6.31506749503757e-29
+  uc=5.52615694e-13 luc=-1.0742296475666e-18
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0213390915869213 lu0=2.11770101418372e-09 wu0=7.95714544953161e-08 pu0=-1.54678950393445e-13
+  a0=1.08865243900813 la0=-2.53831427587913e-07 wa0=-4.25315225253395e-07 pa0=8.26770266370079e-13
+  keta=0.0466423328 lketa=-1.2394759872992e-7
+  a1=0.0
+  a2=0.5
+  ags=-0.20668221991885 lags=7.92435150300254e-07 wags=-1.23479517784484e-06 pags=2.40031834621257e-12
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.1606776136623+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=7.82699159621451e-8
+  nfactor={1.21627378657603+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=6.85092825748608e-08 wnfactor=-4.55446671288959e-06 pnfactor=8.85342784318611e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.47195e-05 lcit=-9.17423605e-12
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.279543725207421 leta0=-2.63872227430706e-07 weta0=-7.55415977804464e-10 peta0=1.46845311925236e-15
+  etab=-0.0293684412 letab=2.772087164868e-8
+  dsub=0.0562216610000004 ldsub=4.605649981821e-7
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.041796294998 lpclm=1.09615456715139e-6
+  pdiblc1=-0.00906932782000003 lpdiblc1=3.85673507489298e-7
+  pdiblc2=0.00602058784087 lpdiblc2=-4.26114512466719e-09 wpdiblc2=-5.29395592033938e-23
+  pdiblcb=-0.41378 lpdiblcb=3.66969442e-7
+  drout=1.556250265901 ldrout=-1.08129489188495e-06 pdrout=1.29246970711411e-26
+  pscbe1=433349461.692 lpscbe1=-126.359101721078
+  pscbe2=1.45323618864e-08 lpscbe2=2.09612945270314e-17
+  pvag=0.0
+  delta=0.01
+  alpha0=-6.40086482779e-05 lalpha0=1.2442660577741e-10 walpha0=3.01906534758944e-25 palpha0=-1.14761350561174e-31
+  alpha1=1.9439e-10 lalpha1=-1.83484721e-16
+  beta0=-41.5076459075 lbeta0=8.65184128795893e-05 wbeta0=2.16840434497101e-19 pbeta0=-2.06795153138257e-25
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-3.33231601733033e-09 lagidl=2.04341135460885e-14 wagidl=1.40321964833749e-13 pagidl=-2.72771867440324e-19
+  bgidl=1031695689.11469 lbgidl=366.239139929958 wbgidl=-3788.84998512597 pbgidl=0.00736514548608638
+  cgidl=65.4911082024591 lcgidl=0.000783506179765242 wcgidl=0.00742524920161967 pcgidl=-1.44339419230285e-8
+  egidl=3.152521570876 legidl=-2.24038668162586e-6
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.5118689035144 lkt1=-1.03281538458358e-07 wkt1=2.80240383515248e-07 pkt1=-5.44759281515263e-13
+  kt2=-0.019032
+  at=270641.73340576 lat=-0.232960345567457 wat=-0.112096153406096 pat=2.17903712606106e-7
+  ute=-1.20470709 lute=-3.79629887748999e-7
+  ua1=6.77542262e-10 lua1=-2.432640431018e-16
+  ub1=-3.52706157e-18 lub1=-2.63667544076999e-25
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=2.81e-6
+  sbref=2.81e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.13 pmos
* DC IV MOS Parameters
+  lmin=8.0e-07 lmax=1e-06 wmin=1.5e-05 wmax=2.0e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.20000030051049+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=1.27136453049752e-07 wvth0=1.69293215681552e-06 pvth0=-1.25937223145506e-12
+  k1=0.590771670000001 lk1=-1.07431583129997e-8
+  k2=0.0323809468307983 lk2=4.57725625256903e-09 wk2=3.92336536921322e-09 pk2=-2.91859149815825e-15
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=7814.73505000002 lvsat=0.0378260986863049
+  ua=-7.95535261990397e-10 lua=2.37947912866466e-15 wua=-1.07247994771281e-15 pua=7.97817833103526e-22
+  ub=1.29210473516165e-17 lub=-9.77291732886754e-24 wub=-1.62432931093101e-22 pub=1.20833857440158e-28
+  uc=6.40846463e-12 luc=-6.601565458257e-18
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0378966189653937 lu0=-1.35109490783564e-08 wu0=-3.97857272476581e-07 pu0=2.95966024995328e-13
+  a0=0.73130260295933 la0=8.34710826585546e-08 wa0=2.126576126267e-06 pa0=-1.58195998033004e-12
+  keta=-0.157135299 lketa=6.83981079260999e-8
+  a1=0.0
+  a2=0.5
+  ags=0.304533174594255 lags=3.09898939419337e-07 wags=6.17397588922416e-06 pags=-4.59282066399386e-12
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.0961094772139999+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=1.73240519685944e-8
+  nfactor={0.456805945619859+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=7.85370977653392e-07 wnfactor=2.2772333564448e-05 pnfactor=-1.69403389385929e-11
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-1.35975e-05 lcit=1.755418025e-11
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=-0.000266262294107083 leta0=2.40419771986259e-10 weta0=3.77707988901835e-09 peta0=-2.80976972944075e-15
+  etab=0.000791398015 letab=-7.470005863585e-10
+  dsub=1.54597013 ldsub=-9.45608581707e-7
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=2.061904095825 lpclm=-8.10625186049219e-7
+  pdiblc1=0.185912130255001 lpdiblc1=2.01630509212305e-7
+  pdiblc2=-0.03533450056535 lpdiblc2=3.47739228219639e-08 wpdiblc2=-1.58818677610181e-22
+  pdiblcb=-0.025
+  drout=0.33218586617 ldrout=7.40994950211363e-8
+  pscbe1=-74402724.1499996 lpscbe1=352.908186495184
+  pscbe2=1.8463592403e-08 lpscbe2=-3.68972719009171e-15
+  pvag=0.0
+  delta=0.01
+  alpha0=0.000255919397305 lalpha0=-1.7755347644829e-10 palpha0=-1.57772181044202e-30
+  alpha1=0.0
+  beta0=68.0295673025 lbeta0=-1.68737626693297e-5
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=4.41901822866519e-08 lagidl=-2.44223726030403e-14 wagidl=-7.01609824168745e-13 pagidl=5.2192754819913e-19
+  bgidl=-21968845.5734406 lbgidl=1360.79309422208 wbgidl=18944.2499256299 pbgidl=-0.0140926275196761
+  cgidl=2292.47618398771 lcgidl=-0.00131854503326846 wcgidl=-0.0371262460080985 pcgidl=2.76182144054245e-8
+  egidl=1.887175135705 legidl=-1.04602618146795e-6
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.538674732428001 lkt1=-7.79795165468112e-08 wkt1=-1.40120191757619e-06 pkt1=1.04235410648493e-12
+  kt2=-0.019032
+  at=19504.4329712 lat=0.0040881523127243 wat=0.560480767030471 pat=-4.16941642593968e-7
+  ute=-2.07964845 lute=4.46227261954998e-7
+  ua1=-7.33113099999999e-11 lua1=4.65466643509001e-16
+  ub1=-4.60795225e-18 lub1=7.56585168775004e-25
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=2.41e-6
+  sbref=2.41e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.14 pmos
* DC IV MOS Parameters
+  lmin=6e-07 lmax=8.0e-07 wmin=1.5e-05 wmax=2.0e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.961308742999998+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-5.04261965823014e-8
+  k1=0.595611254999999 lk1=-1.43433255944998e-8
+  k2=0.035286917 lk2=2.41550504370001e-9
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=61668.4194499998 lvsat=-0.00223565713885499
+  ua=-2.23484979940001e-09 lua=3.45018521304366e-15
+  ub=2.5967598753e-18 lub=-2.09267987523567e-24 wub=5.87747175411144e-39
+  uc=3.13963340000001e-12 luc=-4.16988190626e-18
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.00582160994999997 lu0=1.0349650128195e-8
+  a0=0.945572835 la0=-7.59245429564991e-8
+  keta=0.0210589425000003 lketa=-6.41605883257501e-8
+  a1=0.0
+  a2=0.5
+  ags=-0.717169160000003 lags=1.069943306124e-6
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={0.0170483782755002+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=-6.68540767300445e-8
+  nfactor={2.020420625+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-3.778019823375e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=-0.0642703282430001 leta0=4.78530444313677e-08 weta0=-3.70576914423756e-22 peta0=-1.96426365400032e-28
+  etab=-0.000791398015 letab=4.304413803585e-10
+  dsub=0.18350229023 ldsub=6.79312442979028e-8
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.170632713424999 lpclm=5.96291595318144e-7
+  pdiblc1=0.157259843575 lpdiblc1=2.22944945273558e-7
+  pdiblc2=0.0277574173458 lpdiblc2=-1.21601549121406e-8
+  pdiblcb=-0.025
+  drout=-0.817940921630003 ldrout=9.29678812465559e-7
+  pscbe1=434417012.98 lpscbe1=-25.6028159558223
+  pscbe2=1.03443636915e-08 lpscbe2=2.35016704839316e-15
+  pvag=0.0
+  delta=0.01
+  alpha0=-0.0001310877634225 lalpha0=1.10341150416898e-10 walpha0=8.27180612553028e-25 palpha0=3.94430452610506e-31
+  alpha1=0.0
+  beta0=25.1812730869999 lbeta0=1.50010833975807e-5
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=2.451938855e-08 lagidl=-9.78926914234502e-15
+  bgidl=2079521950 lbgidl=-202.505908605001
+  cgidl=1308.655 lcgidl=-0.0005866804545
+  egidl=-0.296264661400001 legidl=5.78234683598461e-7
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.711541889999998 lkt1=5.06163619709991e-8
+  kt2=-0.019032
+  at=44036.5 lat=-0.01416125235
+  ute=-1.62257375 lute=1.06209392624998e-7
+  ua1=5.53487799999998e-10 lua1=-8.09214420000522e-19
+  ub1=-4.38417814999999e-18 lub1=5.90119615784998e-25
+  uc1=-2.93321028e-10 luc1=1.369676327292e-16 puc1=-1.50463276905253e-36
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=2.02e-6
+  sbref=2.01e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.15 pmos
* DC IV MOS Parameters
+  lmin=5e-07 lmax=6e-07 wmin=1.5e-05 wmax=2.0e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.07757179837928+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=1.28092792384893e-08 wvth0=2.5285661383271e-06 pvth0=-1.37528712263609e-12
+  k1=0.441396800000001 lk1=6.95339164800006e-8
+  k2=0.024199028437464 lk2=8.44620763286337e-09 wk2=6.18105659791205e-07 pk2=-3.36187668360436e-13
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=40338.1873362879 lvsat=0.00936585610779295 wvsat=-0.00904094845664716 pvsat=4.91737186557213e-9
+  ua=1.25025065809079e-08 lua=-4.56546292220581e-15 wua=-1.45498645716295e-16 pua=7.91367134051825e-23
+  ub=-1.27324400496595e-17 lub=6.2448719639498e-24 wub=3.99449135236923e-23 pub=-2.17260384655362e-29
+  uc=-1.17777449999999e-12 luc=-1.82164374945e-18
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0291981318121924 lu0=-2.36484011265145e-09 wu0=2.24207614189764e-07 pu0=-1.21946521357813e-13
+  a0=0.123883260000003 la0=3.70992416885998e-7
+  keta=-0.145889365 lketa=2.66425961235001e-8
+  a1=0.0
+  a2=0.5
+  ags=1.25
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.12509291583+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=1.04565731339369e-8
+  nfactor={8.07972500674621+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-3.67345763556926e-06 wnfactor=-0.000131281424787602 pnfactor=7.14039669419769e-11
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=3.2195e-05 lcit=-1.20718605e-11 wcit=-4.13590306276514e-25
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=-0.374772316090791 leta0=2.16735075621781e-07 weta0=2.95425511084854e-06 peta0=-1.60681935479052e-12
+  etab=0.0170914817 letab=-9.29605689663001e-9
+  dsub=0.43592626954 ldsub=-6.93621580488059e-8
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.957819881500004 lpclm=1.68140494602149e-7
+  pdiblc1=1.77958506268 lpdiblc1=-6.59437741397652e-7
+  pdiblc2=0.00805992596100001 lpdiblc2=-1.4466893479479e-9
+  pdiblcb=-0.025
+  drout=0.854662854460003 ldrout=1.99496186502068e-8
+  pscbe1=497007191.599999 lpscbe1=-59.6456141072404
+  pscbe2=1.5458070132e-08 lpscbe2=-4.31177884594831e-16
+  pvag=0.0
+  delta=0.01
+  alpha0=-4.07586597359999e-05 lalpha0=6.12111509218105e-11
+  alpha1=0.0
+  beta0=44.2272339669998 lbeta0=4.64198527494876e-6
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-2.9092944726336e-08 lagidl=1.93704789266542e-14 wagidl=5.79885906840361e-14 pagidl=-3.15399944730474e-20
+  bgidl=2184885655.144 lbgidl=-259.813227832823 wbgidl=-1317.9225155462 pbgidl=0.000716818056205631
+  cgidl=-10041.9118878284 lcgidl=0.00558689287578988 wcgidl=0.147428084279069 pcgidl=-8.01861350393857e-8
+  egidl=1.2178352726 legidl=-2.4528427050414e-7
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.508294289712001 lkt1=-5.9930007825643e-08 wkt1=-2.63584503109256e-06 pkt1=1.43363611241125e-12
+  kt2=-0.019032
+  at=18000.0
+  ute=-1.6710011 lute=1.32549028290001e-7
+  ua1=5.52e-10
+  ub1=-8.35610879999999e-18 lub1=2.75045269632e-24
+  uc1=-4.1496e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=1.81e-6
+  sbref=1.81e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.16 pmos
* DC IV MOS Parameters
+  lmin=2.0e-05 lmax=1.0e-04 wmin=1.0e-05 wmax=1.5e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.057134+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+  k1=0.59521
+  k2=0.0294389
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=200000.0
+  ua=2.7344678e-9
+  ub=-4.4406e-19
+  uc=-3.9972e-11
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0207994
+  a0=0.911307
+  keta=-0.0079259
+  a1=0.0
+  a2=0.5
+  ags=0.1271299
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.093204657+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.69967+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.08353125
+  pdiblc1=0.39
+  pdiblc2=0.0029407877
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=333712830.0
+  pscbe2=1.5000958e-8
+  pvag=0.0
+  delta=0.01
+  alpha0=5.0667189e-5
+  alpha1=0.0
+  beta0=38.266046
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=7.3657e-9
+  bgidl=1704700000.0
+  cgidl=700.0
+  egidl=0.69350825
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.57573
+  kt2=-0.019032
+  at=430000.0
+  ute=-1.3864
+  ua1=7.0656e-10
+  ub1=-3.145e-18
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.17 pmos
* DC IV MOS Parameters
+  lmin=8e-06 lmax=2.0e-05 wmin=1.0e-05 wmax=1.5e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.057134+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+  k1=0.59521
+  k2=0.0294389
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=200000.0
+  ua=2.7344678e-9
+  ub=-4.4406e-19
+  uc=-3.9972e-11
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0207994
+  a0=0.911307
+  keta=-0.0079259
+  a1=0.0
+  a2=0.5
+  ags=0.1271299
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.093204657+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.69967+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.08353125
+  pdiblc1=0.39
+  pdiblc2=0.0029407877
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=333712830.0
+  pscbe2=1.5000958e-8
+  pvag=0.0
+  delta=0.01
+  alpha0=5.0667189e-5
+  alpha1=0.0
+  beta0=38.266046
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=7.3657e-9
+  bgidl=1704700000.0
+  cgidl=700.0
+  egidl=0.69350825
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.57573
+  kt2=-0.019032
+  at=430000.0
+  ute=-1.3864
+  ua1=7.0656e-10
+  ub1=-3.145e-18
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.18 pmos
* DC IV MOS Parameters
+  lmin=4e-06 lmax=8e-06 wmin=1.0e-05 wmax=1.5e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.06129678645+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=3.30687592801515e-8
+  k1=0.60423167125 lk1=-7.16672542428745e-8
+  k2=0.0278592694525 lk2=1.25484271062853e-8
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=298587.64025 lvsat=-0.783170355381976
+  ua=2.4949572179375e-09 lua=1.9026481128463e-15
+  ub=-2.008594065e-19 lub=-1.93196119470465e-24
+  uc=-5.1678481175e-11 luc=9.29951158060826e-17
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0199748291075 lu0=6.55030871293082e-9
+  a0=0.933098033475 la0=-1.73105790822049e-7
+  keta=-0.0049304093525 lketa=-2.37958781546752e-8
+  a1=0.0
+  a2=0.5
+  ags=0.104081156815 lags=1.83096910987322e-7
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.09479041045225+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=1.25970668493291e-8
+  nfactor={1.7321085775+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-2.57688815802249e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-0.6548060915245 lpclm=5.86527800733648e-06 wpclm=8.470329472543e-22 ppclm=6.46234853557053e-27
+  pdiblc1=0.39
+  pdiblc2=0.0045684231025075 lpdiblc2=-1.29297728739793e-8
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=564147837.55925 lpscbe1=-1830.55265654993
+  pscbe2=-1.558611817795e-08 lpscbe2=2.42980674450017e-13
+  pvag=0.0
+  delta=0.01
+  alpha0=7.83968484975e-05 lalpha0=-2.2028164208219e-10
+  alpha1=0.0
+  beta0=39.148037118575 lbeta0=-7.00644924684789e-6
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=6.5314665525e-09 lagidl=6.62706708359527e-15
+  bgidl=1476348190 lbgidl=1814.00394345899
+  cgidl=934.66205 lcgidl=-0.001864131858995
+  egidl=1.21389074000325 legidl=-4.13386646233682e-6
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.58532353675 lkt1=7.62100965883275e-8
+  kt2=-0.019032
+  at=675202.12275 lat=-1.94786114291372
+  ute=-1.2190800425 lute=-1.32917301038425e-6
+  ua1=1.3814243924e-09 lua1=-5.36105524678636e-15
+  ub1=-2.605671675e-18 lub1=-4.28437028096751e-24
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.19 pmos
* DC IV MOS Parameters
+  lmin=2e-06 lmax=4e-06 wmin=1.0e-05 wmax=1.5e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.0381655746+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-5.815842713506e-8
+  k1=0.602894174 lk1=-6.63922988385996e-8
+  k2=0.0297949601 lk2=4.91425676161003e-9
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=84264.41 lvsat=0.0620990324010002
+  ua=3.28797678225e-09 lua=-1.22494174684578e-15
+  ub=-1.7328156315e-18 lub=4.10992096107285e-24
+  uc=-5.540982305e-11 luc=1.07711155026895e-16
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.02086513804 lu0=3.03901931404402e-9
+  a0=0.8222697474 la0=2.6398988662914e-7
+  keta=-0.00498067579999999 lketa=-2.359763231238e-8
+  a1=0.0
+  a2=0.5
+  ags=0.101458501175 lags=1.93440402565917e-7
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.0635877678486499+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=-1.10463035315009e-7
+  nfactor={2.07037515335+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.59177836429706e-6
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.01798959 leta0=2.44562855999e-7
+  etab=-0.1233522794 letab=2.1041605472566e-7
+  dsub=0.8193648575 ldsub=-1.02290906149425e-6
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=1.0526929389875 lpclm=-8.68927419099802e-7
+  pdiblc1=0.58503867943 lpdiblc1=-7.69213047803977e-7
+  pdiblc2=-0.0011773222896 lpdiblc2=9.73087237795344e-09 ppdiblc2=-2.52435489670724e-29
+  pdiblcb=0.16939 lpdiblcb=-7.66654721e-07 wpdiblcb=-2.11758236813575e-22 ppdiblcb=8.07793566946316e-28
+  drout=0.132342 ldrout=1.6866403862e-6
+  pscbe1=-160819458.431 lpscbe1=1028.64586210602
+  pscbe2=7.662008170125e-08 lpscbe2=-1.2067135725356e-13 ppscbe2=-7.70371977754894e-34
+  pvag=0.0
+  delta=0.01
+  alpha0=4.445374715855e-05 lalpha0=-8.64134447115054e-11
+  alpha1=-9.7195e-11 lalpha1=3.833273605e-16
+  beta0=70.77889717255 lbeta0=-0.00013175539821372
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=9.21504678999999e-09 lagidl=-3.956705015081e-15
+  bgidl=2632410590.0 lbgidl=-2745.390555901
+  cgidl=455.6337275 lcgidl=2.51079421127506e-5
+  egidl=-1.617101386419 legidl=7.0312833850599e-06 wegidl=1.6940658945086e-21
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.56697195 lkt1=3.83327360499981e-9
+  kt2=-0.019032
+  at=210964.1945 lat=-0.11695317768855
+  ute=-1.707821395 lute=5.98374009740499e-7
+  ua1=-4.933329728e-10 lua1=2.03280032582592e-15 wua1=-7.88860905221012e-31 pua1=-3.38542373036819e-36
+  ub1=-3.720478135e-18 lub1=1.12314916626502e-25
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.20 pmos
* DC IV MOS Parameters
+  lmin=1e-06 lmax=2e-06 wmin=1.0e-05 wmax=1.5e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.07950440154749+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=2.22001185681713e-08 wvth0=-2.0737259560867e-07 pvth0=4.03111588603706e-13
+  k1=0.558687465 lk1=1.95411227864996e-8
+  k2=0.0266411723973649 lk2=1.10449046767623e-08 wk2=1.48701188563737e-08 pk2=-2.89060240449047e-14
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=180698.1919 lvsat=-0.12535859623441
+  ua=3.54856039782964e-09 lua=-1.73149023717104e-15 wua=5.67742811870987e-17 pua=-1.10363525199607e-22
+  ub=1.10199481754436e-18 lub=-1.40066707082449e-24 wub=-9.02222839955481e-24 pub=1.75383097858946e-29
+  uc=5.52615694e-13 luc=-1.0742296475666e-18
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0276751678843488 lu0=-1.01989977003856e-08 wu0=-1.49063874389503e-08 pu0=2.89765265425757e-14
+  a0=1.0377004087159 la0=-1.54785775902831e-07 wa0=3.34435389829069e-07 pa0=-6.5010895428873e-13
+  keta=0.0466423328 lketa=-1.2394759872992e-7
+  a1=0.0
+  a2=0.5
+  ags=-0.326928012891223 lags=1.02618094725925e-06 wags=5.58201384762341e-07 pags=-1.08508767183951e-12
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.1606776136623+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=7.82699159621451e-8
+  nfactor={0.836552978195664+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=8.06648561985449e-07 wnfactor=1.10758671406762e-06 pnfactor=-2.15303781347603e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.47195e-05 lcit=-9.17423605000001e-12
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.2794930638759 leta0=-2.63773746868362e-7
+  etab=-0.0293684412 letab=2.772087164868e-8
+  dsub=0.0562216610000001 ldsub=4.605649981821e-7
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.0418196827067856 lpclm=1.09610910378428e-06 wpclm=-3.48736370930545e-10 ppclm=6.77908631455565e-16
+  pdiblc1=-0.00906932782000025 lpdiblc1=3.85673507489298e-7
+  pdiblc2=0.00602058784087 lpdiblc2=-4.26114512466719e-9
+  pdiblcb=-0.41378 lpdiblcb=3.66969442e-7
+  drout=1.556250265901 ldrout=-1.08129489188495e-6
+  pscbe1=433349461.692 lpscbe1=-126.359101721079
+  pscbe2=1.45323618864e-08 lpscbe2=2.0961294527044e-17
+  pvag=0.0
+  delta=0.01
+  alpha0=-6.40086482779e-05 lalpha0=1.2442660577741e-10 walpha0=1.41905821657492e-25 palpha0=3.39726519026063e-31
+  alpha1=1.9439e-10 lalpha1=-1.83484721e-16
+  beta0=-41.5076459075 lbeta0=8.65184128795893e-05 pbeta0=1.55096364853693e-25
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=6.07825748e-09 lagidl=2.14089972462801e-15
+  bgidl=777599680.0 lbgidl=860.176372048
+  cgidl=563.459145 lcgidl=-0.0001844938869655
+  egidl=3.152521570876 legidl=-2.24038668162586e-06 pegidl=1.29246970711411e-26
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.472119432927744 lkt1=-1.80550534331758e-07 wkt1=-3.12467788351572e-07 pkt1=6.07406133776612e-13
+  kt2=-0.019032
+  at=259756.269934816 lat=-0.211800093126289 wat=0.0502180374136447 pat=-9.76188429283846e-8
+  ute=-0.931351549709231 lute=-9.11005722520224e-07 wute=-4.07603070340751e-06 pute=7.92339608435386e-12
+  ua1=9.25601656467831e-10 lua1=-7.25466700007816e-16 wua1=-3.69883744461169e-15 pua1=7.19017010858067e-21
+  ub1=-3.12385747052936e-18 lub1=-1.04745599303798e-24 wub1=-6.01221503480029e-24 pub1=1.16871448061483e-29
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=2.81e-6
+  sbref=2.81e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.21 pmos
* DC IV MOS Parameters
+  lmin=8.0e-07 lmax=1e-06 wmin=1.0e-05 wmax=1.5e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.15600157776254+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=9.44058031975479e-08 wvth0=1.0368629780434e-06 pvth0=-7.71322369366479e-13
+  k1=0.590771670000001 lk1=-1.07431583130005e-8
+  k2=0.0376303235131751 lk2=6.72244938548987e-10 wk2=-7.43505942818686e-08 pk2=5.5309407086282e-14
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=7814.73505000002 lvsat=0.0378260986863049
+  ua=-8.48422624648193e-10 lua=2.41882203774579e-15 wua=-2.83871405935468e-16 pua=2.1117193887541e-22
+  ub=-9.9771979272181e-19 lub=5.81253549805755e-25 wub=4.51111419977739e-23 pub=-3.3558178532144e-29
+  uc=6.40846463e-12 luc=-6.601565458257e-18 puc=1.17549435082229e-38
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.00621623747825611 lu0=1.00560867099253e-08 wu0=7.45319371947515e-08 pu0=-5.54443080791753e-14
+  a0=0.986062754420518 la0=-1.06044994013424e-07 wa0=-1.67217694914534e-06 pa0=1.24393243246923e-12
+  keta=-0.157135299 lketa=6.83981079261001e-8
+  a1=0.0
+  a2=0.5
+  ags=0.905762139456115 lags=-1.37355287541405e-07 wags=-2.7910069238117e-06 pags=2.07623005062352e-12
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.0961094772140001+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=1.73240519685946e-8
+  nfactor={2.35540998752168+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-6.27000569117378e-07 wnfactor=-5.53793357033804e-06 pnfactor=4.11966878297445e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-1.35975e-05 lcit=1.755418025e-11
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=-1.29556365e-05 leta0=5.198494939235e-11
+  etab=0.000791398015 letab=-7.470005863585e-10
+  dsub=1.54597013 ldsub=-9.45608581707e-7
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=2.06178715728107 lpclm=-8.10538195466389e-07 wpclm=1.74368185463917e-09 ppclm=-1.29712493166547e-15
+  pdiblc1=0.185912130255 lpdiblc1=2.01630509212305e-7
+  pdiblc2=-0.03533450056535 lpdiblc2=3.47739228219639e-08 wpdiblc2=7.94093388050907e-23 ppdiblc2=-2.52435489670724e-29
+  pdiblcb=-0.025
+  drout=0.332185866170001 ldrout=7.40994950211371e-8
+  pscbe1=-74402724.1499987 lpscbe1=352.908186495184
+  pscbe2=1.8463592403e-08 lpscbe2=-3.68972719009171e-15
+  pvag=0.0
+  delta=0.01
+  alpha0=0.000255919397305 lalpha0=-1.77553476448289e-10 palpha0=7.88860905221012e-31
+  alpha1=0.0
+  beta0=68.0295673025001 lbeta0=-1.68737626693297e-5
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-2.86268519999999e-09 lagidl=1.058025552028e-14
+  bgidl=1248511200 lbgidl=415.682988320001
+  cgidl=-197.364 lcgidl=0.0005336470796
+  egidl=1.887175135705 legidl=-1.04602618146795e-6
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.737422085361279 lkt1=6.98686393002556e-08 wkt1=1.56233894175784e-06 pkt1=-1.16222393877366e-12
+  kt2=-0.019032
+  at=73931.75032592 lat=-0.0364003290674518 wat=-0.251090187068225 pat=1.86785990160052e-7
+  ute=-3.44642615145384 lute=1.46297319406651e-06 wute=2.03801535170375e-05 pute=-1.51607962013242e-11
+  ua1=-1.31360828233915e-09 lua1=1.38812356123209e-15 wua1=1.84941872230584e-14 pua1=-1.37578258752332e-20
+  ub1=-6.6239727473532e-18 lub1=2.25630281675605e-24 wub1=3.00610751740013e-23 pub1=-2.23624338219395e-29
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=2.41e-6
+  sbref=2.41e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.22 pmos
* DC IV MOS Parameters
+  lmin=6e-07 lmax=8.0e-07 wmin=1.0e-05 wmax=1.5e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.961308743+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-5.04261965822997e-8
+  k1=0.595611255 lk1=-1.43433255945002e-8
+  k2=0.035286917 lk2=2.41550504369998e-9
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=61668.41945 lvsat=-0.00223565713885499
+  ua=-2.2348497994e-09 lua=3.45018521304366e-15
+  ub=2.5967598753e-18 lub=-2.09267987523567e-24 wub=2.93873587705572e-39 pub=5.60519385729927e-45
+  uc=3.13963340000001e-12 luc=-4.16988190626e-18
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.00582160995 lu0=1.0349650128195e-8
+  a0=0.945572835000002 la0=-7.59245429565e-8
+  keta=0.0210589425000001 lketa=-6.41605883257499e-8
+  a1=0.0
+  a2=0.5
+  ags=-0.717169159999999 lags=1.069943306124e-6
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={0.0170483782755001+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=-6.68540767300444e-8
+  nfactor={2.020420625+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-3.778019823375e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=-0.064270328243 leta0=4.78530444313677e-08 weta0=4.46677530778635e-23 peta0=6.3897733322902e-29
+  etab=-0.000791398015 letab=4.304413803585e-10
+  dsub=0.18350229023 ldsub=6.7931244297903e-8
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.170632713424999 lpclm=5.96291595318143e-7
+  pdiblc1=0.157259843575 lpdiblc1=2.22944945273557e-7
+  pdiblc2=0.0277574173458 lpdiblc2=-1.21601549121406e-8
+  pdiblcb=-0.025
+  drout=-0.817940921629999 ldrout=9.29678812465557e-7
+  pscbe1=434417012.98 lpscbe1=-25.6028159558223
+  pscbe2=1.03443636915e-08 lpscbe2=2.35016704839314e-15
+  pvag=0.0
+  delta=0.01
+  alpha0=-0.0001310877634225 lalpha0=1.10341150416898e-10
+  alpha1=0.0
+  beta0=25.1812730870001 lbeta0=1.50010833975807e-5
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=2.451938855e-08 lagidl=-9.789269142345e-15
+  bgidl=2079521950.0 lbgidl=-202.505908605001
+  cgidl=1308.655 lcgidl=-0.000586680454500001
+  egidl=-0.2962646614 legidl=5.7823468359846e-7
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.711541889999999 lkt1=5.0616361971e-8
+  kt2=-0.019032
+  at=44036.5 lat=-0.01416125235
+  ute=-1.62257375 lute=1.06209392625001e-7
+  ua1=5.534878e-10 lua1=-8.09214420000127e-19
+  ub1=-4.38417815e-18 lub1=5.90119615784998e-25
+  uc1=-2.93321028e-10 luc1=1.369676327292e-16 puc1=-7.52316384526264e-37
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=2.02e-6
+  sbref=2.01e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.23 pmos
* DC IV MOS Parameters
+  lmin=5e-07 lmax=6e-07 wmin=1.0e-05 wmax=1.5e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.748626881526373+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-1.66103861037803e-07 wvth0=-2.37636309557857e-06 pvth0=1.29250388768518e-12
+  k1=0.441396799999998 lk1=6.95339164799997e-8
+  k2=0.0860832029288735 lk2=-2.52125948730143e-08 wk2=-3.04655206930955e-07 pk2=1.65701967049747e-13
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=68741.5210748505 lvsat=-0.00608271711261121 wvsat=-0.432565784552398 pvsat=2.35272530218048e-7
+  ua=1.25434050896128e-08 lua=-4.5877076210904e-15 wua=-7.55340235272042e-16 pua=4.10829553964425e-22
+  ub=-9.15935392822717e-18 lub=4.30147042250276e-24 wub=-1.33337166492529e-23 pub=7.25220848552868e-30
+  uc=-1.17777449999998e-12 luc=-1.82164374945e-18
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0443876170266114 lu0=-1.0626401120774e-08 wu0=-2.28425803301843e-09 pu0=1.24240794415867e-15
+  a0=0.123883259999998 la0=3.70992416886001e-7
+  keta=-0.145889365 lketa=2.66425961235001e-8
+  a1=0.0
+  a2=0.5
+  ags=1.25
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.12509291583+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=1.04565731339369e-8
+  nfactor={-3.64681182337477+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=2.70460574633354e-06 wnfactor=4.35740916338672e-05 pnfactor=-2.36999484396604e-11
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=3.2195e-05 lcit=-1.20718605e-11
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=-0.218909642151327 leta0=1.31961367266106e-07 weta0=6.30171816920492e-07 peta0=-3.42750451223055e-13
+  etab=-0.0133999391361006 letab=7.28822689612515e-09 wetab=4.54660503263497e-07 petab=-2.47289847725016e-13
+  dsub=0.435926269539999 ldsub=-6.93621580488063e-8
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.0171991885212819 lpclm=6.79744089513276e-07 wpclm=1.40256854525922e-05 ppclm=-7.62857031766493e-12
+  pdiblc1=1.77958506268 lpdiblc1=-6.59437741397653e-7
+  pdiblc2=0.00805992596099998 lpdiblc2=-1.4466893479479e-9
+  pdiblcb=-0.025
+  drout=0.854662854459999 ldrout=1.9949618650206e-8
+  pscbe1=497007191.599999 lpscbe1=-59.6456141072399
+  pscbe2=1.5458070132e-08 lpscbe2=-4.31177884594793e-16
+  pvag=0.0
+  delta=0.01
+  alpha0=-4.07586597360001e-05 lalpha0=6.12111509218104e-11
+  alpha1=0.0
+  beta0=44.2272339669998 lbeta0=4.6419852749487e-6
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-7.94766592056384e-08 lagidl=4.67741812319468e-14 wagidl=8.09264994121505e-13 pagidl=-4.40159230302687e-19
+  bgidl=1548318174.90576 lbgidl=86.4158246687584 wbgidl=8173.99629276426 pbgidl=-0.00444583658363444
+  cgidl=-614.08402770336 lcgidl=0.000459097302667858 wcgidl=0.00684883798526954 pcgidl=-3.72508298018811e-9
+  egidl=1.2178352726 legidl=-2.4528427050414e-7
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.685064999999998 lkt1=3.62155814999996e-8
+  kt2=-0.019032
+  at=18000.0
+  ute=-1.6710011 lute=1.32549028290001e-7
+  ua1=5.52e-10
+  ub1=-8.35610879999999e-18 lub1=2.75045269632e-24
+  uc1=-4.1496e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=1.81e-6
+  sbref=1.81e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.24 pmos
* DC IV MOS Parameters
+  lmin=2.0e-05 lmax=1.0e-04 wmin=7e-06 wmax=1.0e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.057134+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+  k1=0.59521
+  k2=0.0294389
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=200000.0
+  ua=2.7344678e-9
+  ub=-4.4406e-19
+  uc=-3.9972e-11
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0207994
+  a0=0.911307
+  keta=-0.0079259
+  a1=0.0
+  a2=0.5
+  ags=0.1271299
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.093204657+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.69967+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.08353125
+  pdiblc1=0.39
+  pdiblc2=0.0029407877
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=333712830.0
+  pscbe2=1.5000958e-8
+  pvag=0.0
+  delta=0.01
+  alpha0=5.0667189e-5
+  alpha1=0.0
+  beta0=38.266046
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=7.3657e-9
+  bgidl=1704700000.0
+  cgidl=700.0
+  egidl=0.69350825
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.57573
+  kt2=-0.019032
+  at=430000.0
+  ute=-1.3864
+  ua1=7.0656e-10
+  ub1=-3.145e-18
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.25 pmos
* DC IV MOS Parameters
+  lmin=8e-06 lmax=2.0e-05 wmin=7e-06 wmax=1.0e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.057134+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+  k1=0.59521
+  k2=0.0294389
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=200000.0
+  ua=2.7344678e-9
+  ub=-4.4406e-19
+  uc=-3.9972e-11
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0207994
+  a0=0.911307
+  keta=-0.0079259
+  a1=0.0
+  a2=0.5
+  ags=0.1271299
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.093204657+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.69967+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.08353125
+  pdiblc1=0.39
+  pdiblc2=0.0029407877
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=333712830.0
+  pscbe2=1.5000958e-8
+  pvag=0.0
+  delta=0.01
+  alpha0=5.0667189e-5
+  alpha1=0.0
+  beta0=38.266046
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=7.3657e-9
+  bgidl=1704700000.0
+  cgidl=700.0
+  egidl=0.69350825
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.57573
+  kt2=-0.019032
+  at=430000.0
+  ute=-1.3864
+  ua1=7.0656e-10
+  ub1=-3.145e-18
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.26 pmos
* DC IV MOS Parameters
+  lmin=4e-06 lmax=8e-06 wmin=7e-06 wmax=1.0e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.06129678645+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=3.30687592801549e-8
+  k1=0.60423167125 lk1=-7.16672542428762e-8
+  k2=0.0278592694525 lk2=1.25484271062852e-8
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=298587.64025 lvsat=-0.783170355381975
+  ua=2.4949572179375e-09 lua=1.90264811284629e-15
+  ub=-2.008594065e-19 lub=-1.93196119470465e-24
+  uc=-5.1678481175e-11 luc=9.29951158060824e-17
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0199748291075 lu0=6.55030871293082e-9
+  a0=0.933098033475 la0=-1.73105790822049e-7
+  keta=-0.00493040935250001 lketa=-2.37958781546752e-8
+  a1=0.0
+  a2=0.5
+  ags=0.104081156815 lags=1.83096910987321e-7
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.09479041045225+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=1.25970668493291e-8
+  nfactor={1.7321085775+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-2.57688815802249e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-0.6548060915245 lpclm=5.86527800733648e-06 wpclm=-4.2351647362715e-22 ppclm=9.69352280335579e-27
+  pdiblc1=0.39
+  pdiblc2=0.0045684231025075 lpdiblc2=-1.29297728739793e-8
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=564147837.55925 lpscbe1=-1830.55265654993 ppscbe1=6.93889390390723e-18
+  pscbe2=-1.558611817795e-08 lpscbe2=2.42980674450017e-13
+  pvag=0.0
+  delta=0.01
+  alpha0=7.83968484975e-05 lalpha0=-2.2028164208219e-10
+  alpha1=0.0
+  beta0=39.148037118575 lbeta0=-7.00644924684799e-6
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=6.5314665525e-09 lagidl=6.62706708359525e-15
+  bgidl=1476348190.0 lbgidl=1814.003943459
+  cgidl=934.662049999999 lcgidl=-0.001864131858995
+  egidl=1.21389074000325 legidl=-4.13386646233682e-6
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.58532353675 lkt1=7.62100965883258e-8
+  kt2=-0.019032
+  at=675202.12275 lat=-1.94786114291372
+  ute=-1.2190800425 lute=-1.32917301038424e-6
+  ua1=1.3814243924e-09 lua1=-5.36105524678636e-15
+  ub1=-2.605671675e-18 lub1=-4.2843702809675e-24
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.27 pmos
* DC IV MOS Parameters
+  lmin=2e-06 lmax=4e-06 wmin=7e-06 wmax=1.0e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.0381655746+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-5.815842713506e-8
+  k1=0.602894174 lk1=-6.63922988385996e-8
+  k2=0.0297949601 lk2=4.91425676160998e-9
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=84264.4099999999 lvsat=0.0620990324009998
+  ua=3.28797678225e-09 lua=-1.22494174684578e-15
+  ub=-1.7328156315e-18 lub=4.10992096107285e-24
+  uc=-5.540982305e-11 luc=1.07711155026895e-16
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.02086513804 lu0=3.03901931404402e-9
+  a0=0.8222697474 la0=2.63989886629138e-7
+  keta=-0.0049806758 lketa=-2.359763231238e-8
+  a1=0.0
+  a2=0.5
+  ags=0.101458501175 lags=1.93440402565918e-7
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.0635877678486498+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=-1.10463035315009e-7
+  nfactor={2.07037515335+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.59177836429707e-6
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.0179895899999999 leta0=2.44562855999e-7
+  etab=-0.1233522794 letab=2.1041605472566e-7
+  dsub=0.8193648575 ldsub=-1.02290906149425e-06 wdsub=-3.3881317890172e-21
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=1.0526929389875 lpclm=-8.68927419099803e-7
+  pdiblc1=0.58503867943 lpdiblc1=-7.69213047803977e-7
+  pdiblc2=-0.0011773222896 lpdiblc2=9.73087237795344e-09 ppdiblc2=-1.26217744835362e-29
+  pdiblcb=0.16939 lpdiblcb=-7.66654721e-07 wpdiblcb=2.11758236813575e-22 ppdiblcb=-1.61558713389263e-27
+  drout=0.132342 ldrout=1.6866403862e-6
+  pscbe1=-160819458.431 lpscbe1=1028.64586210602
+  pscbe2=7.662008170125e-08 lpscbe2=-1.2067135725356e-13
+  pvag=0.0
+  delta=0.01
+  alpha0=4.445374715855e-05 lalpha0=-8.64134447115054e-11
+  alpha1=-9.7195e-11 lalpha1=3.833273605e-16
+  beta0=70.77889717255 lbeta0=-0.00013175539821372
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=9.21504678999999e-09 lagidl=-3.95670501508101e-15
+  bgidl=2632410590 lbgidl=-2745.390555901
+  cgidl=455.6337275 lcgidl=2.51079421127506e-5
+  egidl=-1.617101386419 legidl=7.0312833850599e-06 wegidl=-1.6940658945086e-21
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.56697195 lkt1=3.83327360500066e-9
+  kt2=-0.019032
+  at=210964.1945 lat=-0.11695317768855
+  ute=-1.707821395 lute=5.98374009740503e-7
+  ua1=-4.933329728e-10 lua1=2.03280032582592e-15 pua1=-1.88079096131566e-36
+  ub1=-3.72047813499999e-18 lub1=1.12314916626502e-25
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.28 pmos
* DC IV MOS Parameters
+  lmin=1e-06 lmax=2e-06 wmin=7e-06 wmax=1.0e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.1004276774+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=6.28728744978609e-8
+  k1=0.558687465 lk1=1.95411227864996e-8
+  k2=0.028141523 lk2=8.12837314030003e-9
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=180698.1919 lvsat=-0.12535859623441
+  ua=3.55428875332e-09 lua=-1.74262558740875e-15
+  ub=1.91678905e-19 lub=3.68896031570501e-25
+  uc=5.52615694e-13 luc=-1.0742296475666e-18
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.02617115789 lu0=-7.27535267237097e-9
+  a0=1.0714439412 la0=-2.2037982869868e-7
+  keta=0.0466423328 lketa=-1.2394759872992e-07 wketa=-1.05879118406788e-22 pketa=2.01948391736579e-28
+  a1=0.0
+  a2=0.5
+  ags=-0.2706071595 lags=9.1669884035205e-07 pags=-1.61558713389263e-27
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.1606776136623+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=7.82699159621449e-8
+  nfactor={0.948305171299999+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=5.8941347380993e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.47195e-05 lcit=-9.17423605e-12
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.2794930638759 leta0=-2.63773746868362e-7
+  etab=-0.0293684412 letab=2.772087164868e-8
+  dsub=0.0562216610000001 ldsub=4.605649981821e-7
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.0417844962479998 lpclm=1.09617750274151e-6
+  pdiblc1=-0.00906932782000003 lpdiblc1=3.85673507489298e-7
+  pdiblc2=0.00602058784087 lpdiblc2=-4.2611451246672e-9
+  pdiblcb=-0.41378 lpdiblcb=3.66969442e-7
+  drout=1.556250265901 ldrout=-1.08129489188495e-6
+  pscbe1=433349461.692 lpscbe1=-126.359101721079
+  pscbe2=1.45323618864e-08 lpscbe2=2.0961294527044e-17
+  pvag=0.0
+  delta=0.01
+  alpha0=-6.40086482779e-05 lalpha0=1.2442660577741e-10 walpha0=9.33845650991582e-26 palpha0=-1.86169717147638e-31
+  alpha1=1.9439e-10 lalpha1=-1.83484721e-16
+  beta0=-41.5076459075 lbeta0=8.65184128795893e-05 wbeta0=-2.71050543121376e-20 pbeta0=-1.03397576569128e-25
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=6.07825748e-09 lagidl=2.140899724628e-15
+  bgidl=777599680.0 lbgidl=860.176372047999
+  cgidl=563.459145 lcgidl=-0.0001844938869655
+  egidl=3.152521570876 legidl=-2.24038668162586e-6
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.5036465 lkt1=-1.1926506865e-7
+  kt2=-0.019032
+  at=264823.12 lat=-0.221649542968
+  ute=-1.34261088 lute=-1.11558710368001e-7
+  ua1=5.524e-10
+  ub1=-3.73047202e-18 lub1=1.31742029678002e-25
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=2.81e-6
+  sbref=2.81e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.29 pmos
* DC IV MOS Parameters
+  lmin=8.0e-07 lmax=1e-06 wmin=7e-06 wmax=1.0e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.0513851985+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=1.65816786641499e-8
+  k1=0.590771669999999 lk1=-1.07431583129997e-8
+  k2=0.0301285705 lk2=6.25279900505005e-9
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=7814.73505000002 lvsat=0.0378260986863052
+  ua=-8.77064402099999e-10 lua=2.44012865599219e-15
+  ub=3.55385977e-18 lub=-2.804666486903e-24 wub=1.17549435082229e-38
+  uc=6.40846463e-12 luc=-6.601565458257e-18 wuc=-1.23259516440783e-32 puc=5.87747175411144e-39
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.01373628745 lu0=4.46192153594499e-9
+  a0=0.817345092000002 la0=1.94640750612005e-8
+  keta=-0.157135299 lketa=6.83981079261001e-8
+  a1=0.0
+  a2=0.5
+  ags=0.6241578725 lags=7.21301266472508e-8
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.0961094772140001+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=1.73240519685946e-8
+  nfactor={1.796649022+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-2.113382868658e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-1.35975e-05 lcit=1.755418025e-11
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=-1.29556365e-05 leta0=5.198494939235e-11
+  etab=0.000791398015 letab=-7.470005863585e-10
+  dsub=1.54597013 ldsub=-9.45608581707e-7
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=2.061963089575 lpclm=-8.10669071499842e-7
+  pdiblc1=0.185912130255 lpdiblc1=2.01630509212305e-7
+  pdiblc2=-0.03533450056535 lpdiblc2=3.47739228219639e-08 wpdiblc2=2.64697796016969e-23 ppdiblc2=-2.52435489670724e-29
+  pdiblcb=-0.025
+  drout=0.33218586617 ldrout=7.40994950211379e-8
+  pscbe1=-74402724.1500006 lpscbe1=352.908186495185
+  pscbe2=1.8463592403e-08 lpscbe2=-3.68972719009169e-15
+  pvag=0.0
+  delta=0.01
+  alpha0=0.000255919397305 lalpha0=-1.77553476448289e-10
+  alpha1=0.0
+  beta0=68.0295673024999 lbeta0=-1.68737626693297e-5
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-2.8626852e-09 lagidl=1.058025552028e-14
+  bgidl=1248511200.0 lbgidl=415.682988320001
+  cgidl=-197.364 lcgidl=0.0005336470796
+  egidl=1.887175135705 legidl=-1.04602618146795e-6
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.57978675 lkt1=-4.73962866749997e-8
+  kt2=-0.019032
+  at=48597.5 lat=-0.01755418025
+  ute=-1.3901295 lute=-6.6705884950002e-8
+  ua1=5.524e-10
+  ub1=-3.5909e-18
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=2.41e-6
+  sbref=2.41e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.30 pmos
* DC IV MOS Parameters
+  lmin=6e-07 lmax=8.0e-07 wmin=7e-06 wmax=1.0e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.961308742999998+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-5.04261965822997e-8
+  k1=0.595611254999999 lk1=-1.43433255944998e-8
+  k2=0.0352869169999999 lk2=2.41550504370001e-9
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=61668.4194499999 lvsat=-0.00223565713885499
+  ua=-2.23484979940001e-09 lua=3.45018521304366e-15
+  ub=2.5967598753e-18 lub=-2.09267987523567e-24 wub=-2.93873587705572e-39 pub=1.40129846432482e-45
+  uc=3.13963340000002e-12 luc=-4.16988190626e-18
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.00582160994999997 lu0=1.0349650128195e-8
+  a0=0.945572835 la0=-7.59245429565e-8
+  keta=0.0210589425000002 lketa=-6.416058832575e-8
+  a1=0.0
+  a2=0.5
+  ags=-0.717169159999999 lags=1.069943306124e-6
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={0.0170483782755002+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=-6.68540767300446e-8
+  nfactor={2.020420625+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-3.778019823375e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=-0.064270328243 leta0=4.78530444313677e-08 weta0=-4.46677530778635e-23 peta0=1.0097419586829e-28
+  etab=-0.000791398015 letab=4.304413803585e-10
+  dsub=0.18350229023 ldsub=6.7931244297903e-8
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.170632713424999 lpclm=5.96291595318145e-7
+  pdiblc1=0.157259843575 lpdiblc1=2.22944945273557e-7
+  pdiblc2=0.0277574173458 lpdiblc2=-1.21601549121406e-8
+  pdiblcb=-0.025
+  drout=-0.817940921630002 ldrout=9.29678812465558e-7
+  pscbe1=434417012.98 lpscbe1=-25.6028159558218
+  pscbe2=1.03443636915e-08 lpscbe2=2.35016704839314e-15
+  pvag=0.0
+  delta=0.01
+  alpha0=-0.0001310877634225 lalpha0=1.10341150416898e-10 walpha0=2.06795153138257e-25
+  alpha1=0.0
+  beta0=25.1812730869998 lbeta0=1.50010833975807e-5
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=2.451938855e-08 lagidl=-9.789269142345e-15
+  bgidl=2079521950 lbgidl=-202.505908605001
+  cgidl=1308.655 lcgidl=-0.0005866804545
+  egidl=-0.296264661400001 legidl=5.7823468359846e-7
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.711541889999998 lkt1=5.0616361971e-8
+  kt2=-0.019032
+  at=44036.4999999999 lat=-0.01416125235
+  ute=-1.62257375 lute=1.06209392624999e-7
+  ua1=5.53487799999998e-10 lua1=-8.09214420000522e-19
+  ub1=-4.38417815e-18 lub1=5.90119615784998e-25
+  uc1=-2.93321028e-10 luc1=1.369676327292e-16
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=2.02e-6
+  sbref=2.01e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.31 pmos
* DC IV MOS Parameters
+  lmin=5e-07 lmax=6e-07 wmin=7e-06 wmax=1.0e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.925688266085661+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-6.98001739760075e-08 wvth0=-6.21490715318524e-07 pvth0=3.38028800061769e-13
+  k1=0.441396799999998 lk1=6.95339164799989e-8
+  k2=0.0522663403672186 lk2=-6.81960332573027e-09 wk2=3.05069643364121e-08 pk2=-1.65927379025744e-14
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=-4417.69817220443 lvsat=0.0337085822358619 wvsat=0.292522260690212 pvsat=-1.59102857589407e-7
+  ua=1.23472820505605e-08 lua=-4.48103630014984e-15 wua=1.18845403258731e-15 pua=-6.46400148324212e-22
+  ub=-1.32945348469218e-17 lub=6.55059532418079e-24 wub=2.76504584132981e-23 pub=-1.50390843309929e-29
+  uc=-1.17777450000001e-12 luc=-1.82164374945e-18
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0425556298102994 lu0=-9.62998327382186e-09 wu0=1.58727431386233e-08 pu0=-8.63318499309724e-15
+  a0=0.123883259999998 la0=3.70992416886001e-7
+  keta=-0.145889365 lketa=2.66425961235001e-8
+  a1=0.0
+  a2=0.5
+  ags=1.25
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.12509291583+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=1.0456573133937e-8
+  nfactor={1.2773516544768+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=2.63532307300673e-08 wnfactor=-5.2297653148136e-06 pnfactor=2.84446935472711e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=3.2195e-05 lcit=-1.20718605e-11
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.00840319440352788 leta0=8.32591546392119e-09 weta0=-1.62274752820698e-06 peta0=8.82612380591777e-13
+  etab=0.0679105164268344 letab=-3.69365298845552e-08 wetab=-3.51215227624487e-07 petab=1.91025962304958e-13
+  dsub=0.435926269539999 ldsub=-6.93621580488059e-8
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=2.52584929486457 lpclm=-6.84710703326843e-07 wpclm=-1.08377865817864e-05 ppclm=5.89467212183362e-12
+  pdiblc1=1.77958506268 lpdiblc1=-6.59437741397653e-7
+  pdiblc2=0.00805992596099998 lpdiblc2=-1.4466893479479e-9
+  pdiblcb=-0.025
+  drout=0.854662854459997 ldrout=1.9949618650206e-8
+  pscbe1=497007191.6 lpscbe1=-59.6456141072399
+  pscbe2=1.5458070132e-08 lpscbe2=-4.31177884594831e-16
+  pvag=0.0
+  delta=0.01
+  alpha0=-4.07586597360001e-05 lalpha0=6.12111509218103e-11
+  alpha1=0.0
+  beta0=44.2272339669998 lbeta0=4.6419852749487e-6
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=2.97862825296e-08 lagidl=-1.26539327778494e-14 wagidl=-2.7365051065885e-13 pagidl=1.48838512747349e-19
+  bgidl=2373050000.0 lbgidl=-362.155815
+  cgidl=-848.31591114304 lcgidl=0.0005864960240707 wcgidl=0.00917033266830103 pcgidl=-4.98774393828893e-9
+  egidl=1.2178352726 legidl=-2.4528427050414e-7
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.685065 lkt1=3.62155814999996e-8
+  kt2=-0.019032
+  at=18000.0
+  ute=-1.67100109999999 lute=1.32549028289999e-7
+  ua1=5.52e-10
+  ub1=-8.35610879999999e-18 lub1=2.75045269632e-24
+  uc1=-4.1496e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=1.81e-6
+  sbref=1.81e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.32 pmos
* DC IV MOS Parameters
+  lmin=2.0e-05 lmax=1.0e-04 wmin=5.0e-06 wmax=7.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.078494812052+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} wvth0=1.47626622729329e-7
+  k1=0.59521
+  k2=0.0297438790616 wk2=-2.10773957270752e-9
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=200000.0
+  ua=2.778260043032e-09 wua=-3.02652395649487e-16
+  ub=-3.874596186e-19 wub=-3.91170669492014e-25
+  uc=-3.9972e-11
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0218710011472 wu0=-7.40593840200932e-9
+  a0=0.90251613816 wa0=6.07544900989777e-8
+  keta=-0.0079259
+  a1=0.0
+  a2=0.5
+  ags=0.12450860251 wags=1.81160385979492e-8
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.093204657+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.62236934896+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} wnfactor=5.34232220199943e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.08353125
+  pdiblc1=0.39
+  pdiblc2=0.0029407877
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=333712830.0
+  pscbe2=1.5000958e-8
+  pvag=0.0
+  delta=0.01
+  alpha0=5.0667189e-5
+  alpha1=0.0
+  beta0=38.266046
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-1.22794206644e-08 wagidl=1.35769314843252e-13
+  bgidl=1704700000.0
+  cgidl=-36.6643999999997 wcgidl=0.0050911583881824
+  egidl=0.69350825
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.57506700204 wkt1=-4.58204254936249e-9
+  kt2=-0.019032
+  at=383835.6976 wat=0.319045925659431
+  ute=-1.0188044644 wute=-2.54048803570302e-6
+  ua1=2.387294206272e-09 wua1=-1.16157154500296e-14
+  ub1=-1.8737628004e-18 wub1=-8.78564232520676e-24
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.33 pmos
* DC IV MOS Parameters
+  lmin=8e-06 lmax=2.0e-05 wmin=5.0e-06 wmax=7.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.078494812052+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} wvth0=1.47626622729325e-7
+  k1=0.59521
+  k2=0.0297438790616 wk2=-2.10773957270752e-9
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=200000.0
+  ua=2.778260043032e-09 wua=-3.02652395649487e-16
+  ub=-3.874596186e-19 wub=-3.91170669492016e-25
+  uc=-3.9972e-11
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0218710011472 wu0=-7.40593840200932e-9
+  a0=0.90251613816 wa0=6.07544900989777e-8
+  keta=-0.0079259
+  a1=0.0
+  a2=0.5
+  ags=0.12450860251 wags=1.81160385979492e-8
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.093204657+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.62236934896+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} wnfactor=5.34232220199943e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.08353125
+  pdiblc1=0.39
+  pdiblc2=0.0029407877
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=333712830.0
+  pscbe2=1.5000958e-8
+  pvag=0.0
+  delta=0.01
+  alpha0=5.0667189e-5
+  alpha1=0.0
+  beta0=38.266046
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-1.22794206644e-08 wagidl=1.35769314843252e-13
+  bgidl=1704700000.0
+  cgidl=-36.6643999999992 wcgidl=0.0050911583881824
+  egidl=0.69350825
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.57506700204 wkt1=-4.58204254936249e-9
+  kt2=-0.019032
+  at=383835.6976 wat=0.319045925659431
+  ute=-1.0188044644 wute=-2.54048803570302e-6
+  ua1=2.387294206272e-09 wua1=-1.16157154500296e-14
+  ub1=-1.8737628004e-18 wub1=-8.78564232520677e-24
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.34 pmos
* DC IV MOS Parameters
+  lmin=4e-06 lmax=8e-06 wmin=5.0e-06 wmax=7.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.08332340346031+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=3.8357847288455e-08 wvth0=1.52228064713471e-07 pvth0=-3.65533949778131e-14
+  k1=0.60423167125 lk1=-7.16672542428728e-8
+  k2=0.0267459628974581 lk2=2.3815146216327e-08 wk2=7.69416847932384e-09 pk2=-7.78653773745343e-14
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=358873.25283857 lvsat=-1.26207323322432 wvsat=-0.416639656018415 pvsat=3.30974376344469e-6
+  ua=2.57773899932799e-09 lua=1.59291911908029e-15 wua=-5.72112838240672e-16 pua=2.14056680990016e-21
+  ub=-9.54252577943193e-20 lub=-2.31989175880425e-24 wub=-7.28665523383239e-25 pub=2.68102536982648e-30
+  uc=-5.1678481175e-11 luc=9.29951158060826e-17
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0213599638623393 lu0=4.05962908720456e-09 wu0=-9.57279926363126e-09 pu0=1.7213325998638e-14
+  a0=0.928302001384846 la0=-2.04840318871846e-07 wa0=3.31458381941393e-08 pa0=2.19320369866775e-13
+  keta=-0.00493040935250001 lketa=-2.37958781546752e-8
+  a1=0.0
+  a2=0.5
+  ags=0.0908607286105325 lags=2.6729534546998e-07 wags=9.13676484821829e-08 pags=-5.81903463759359e-13
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.09479041045225+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=1.25970668493282e-8
+  nfactor={1.5537992615124+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=5.44713917674957e-07 wnfactor=1.23231280048461e-06 pnfactor=-5.54548232172338e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-0.6548060915245 lpclm=5.86527800733647e-06 ppclm=4.8467614016779e-27
+  pdiblc1=0.39
+  pdiblc2=0.0045684231025075 lpdiblc2=-1.29297728739793e-8
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=564147837.55925 lpscbe1=-1830.55265654993
+  pscbe2=-1.558611817795e-08 lpscbe2=2.42980674450017e-13 ppscbe2=-3.85185988877447e-34
+  pvag=0.0
+  delta=0.01
+  alpha0=7.83968484975e-05 lalpha0=-2.2028164208219e-10 palpha0=7.88860905221012e-31
+  alpha1=0.0
+  beta0=39.1480371185751 lbeta0=-7.00644924684778e-6
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-3.32478381620127e-08 lagidl=1.66571011759286e-13 wagidl=2.7491859369525e-13 pagidl=-1.10538795627238e-18
+  bgidl=1295975574.02215 lbgidl=3246.86596752545 wbgidl=1246.57246479406 pbgidl=-0.0099026470030775
+  cgidl=-48.9554618085976 lcgidl=9.76389659013317e-05 wcgidl=0.00679787505139036 pcgidl=-1.35579865008578e-8
+  egidl=1.21389074000325 legidl=-4.13386646233682e-6
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.608217928769389 lkt1=2.63347646845594e-07 wkt1=1.58225341107632e-07 pkt1=-1.2933255750328e-12
+  kt2=-0.019032
+  at=715205.087499687 lat=-2.63236529642412 wat=-0.2764643296697 pat=4.73067391730909e-6
+  ute=-0.489044498686791 lute=-4.20836019162916e-06 wute=-5.0453457267053e-06 pute=1.9898339011553e-11
+  ua1=4.71932050770103e-09 lua1=-1.85253837359221e-14 wua1=-2.30685204908725e-14 pua1=9.09799379639521e-20
+  ub1=-5.27963087719173e-19 lub1=-1.06908983375652e-23 wub1=-1.43592435067222e-23 pub1=4.42761304258405e-29
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.35 pmos
* DC IV MOS Parameters
+  lmin=2e-06 lmax=4e-06 wmin=5.0e-06 wmax=7.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.06740254912702+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-2.44324101165854e-08 wvth0=2.02059537705816e-07 pvth0=-2.3308374131231e-13
+  k1=0.602894174 lk1=-6.63922988386004e-8
+  k2=0.0322591734833372 lk2=2.07159498667843e-09 wk2=-1.70304152567282e-08 pk2=1.96459084220831e-14
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=-12440.11639114 lvsat=0.202349563680737 wvsat=0.668334265523702 pvsat=-9.69284885725264e-7
+  ua=3.14556735758786e-09 lua=-6.46539143060809e-16 wua=9.84205205144824e-16 pua=-3.99739592140789e-21
+  ub=-1.54800834740066e-18 lub=3.40895068829419e-24 wub=-1.27722088190982e-24 pub=4.84447284831951e-30
+  uc=-5.540982305e-11 luc=1.07711155026895e-16
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0213824654032186 lu0=3.97088526013084e-09 wu0=-3.57529907063061e-09 pu0=-6.44021501253672e-15
+  a0=0.723779673430536 la0=6.01775290347153e-07 wa0=6.80674356250064e-07 pa0=-2.33446735249393e-12
+  keta=-0.0049806758 lketa=-2.359763231238e-8
+  a1=0.0
+  a2=0.5
+  ags=0.10014304900978 lags=2.30686802047389e-07 wags=9.09121619724512e-09 pags=-2.57413442470797e-13
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.0635877678486502+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=-1.10463035315009e-7
+  nfactor={1.99700539229103+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.20324674150286e-06 wnfactor=5.07065462175618e-07 pnfactor=-2.68517934416656e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.01798959 leta0=2.44562855999e-7
+  etab=-0.1233522794 letab=2.1041605472566e-7
+  dsub=0.819364857500001 ldsub=-1.02290906149425e-6
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=1.0526929389875 lpclm=-8.689274190998e-7
+  pdiblc1=0.58503867943 lpdiblc1=-7.69213047803977e-7
+  pdiblc2=-0.0011773222896 lpdiblc2=9.73087237795344e-09 ppdiblc2=1.26217744835362e-29
+  pdiblcb=0.16939 lpdiblcb=-7.66654721e-07 wpdiblcb=1.05879118406788e-22 ppdiblcb=2.01948391736579e-28
+  drout=0.132342 ldrout=1.6866403862e-6
+  pscbe1=-160819458.431 lpscbe1=1028.64586210602
+  pscbe2=7.662008170125e-08 lpscbe2=-1.2067135725356e-13 ppscbe2=3.85185988877447e-34
+  pvag=0.0
+  delta=0.01
+  alpha0=4.445374715855e-05 lalpha0=-8.64134447115054e-11
+  alpha1=-9.7195e-11 lalpha1=3.833273605e-16
+  beta0=70.77889717255 lbeta0=-0.00013175539821372
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=1.67648326318183e-08 lagidl=-3.06739605845042e-14 wagidl=-5.21772947322467e-14 pagidl=1.84645518096819e-19
+  bgidl=2993155821.9557 lbgidl=-3446.64321229969 wbgidl=-2493.14492958811 pbgidl=0.00484642442862633
+  cgidl=-503.1254124628 lcgidl=0.00188883983428644 wcgidl=0.00662607645716035 pcgidl=-1.2880430025074e-8
+  egidl=-1.617101386419 legidl=7.0312833850599e-06 wegidl=-8.470329472543e-22 pegidl=-1.29246970711411e-26
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.54241647 lkt1=3.83327360500066e-09 wkt1=-1.6970527960608e-07 pkt1=6.46234853557053e-27
+  kt2=-0.019032
+  at=-162190.850332654 lat=0.827996542792846 wat=2.57891033772278 pat=-6.5306382334201e-6
+  ute=-1.82667755495428 lute=1.06713081898418e-06 wute=8.21426331635391e-07 pute=-3.23962330933681e-12
+  ua1=-4.933329728e-10 lua1=2.03280032582592e-15 wua1=-3.94430452610506e-31 pua1=-3.76158192263132e-37
+  ub1=-2.65524181732696e-18 lub1=-2.30112375586508e-24 wub1=-7.36195045412487e-24 pub1=1.66795063557019e-29
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.36 pmos
* DC IV MOS Parameters
+  lmin=1e-06 lmax=2e-06 wmin=5.0e-06 wmax=7.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.16826879607857+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=1.71641487332519e-07 wvth0=4.68856483934966e-07 pvth0=-7.51710325087159e-13
+  k1=0.558687465 lk1=1.95411227864996e-8
+  k2=0.0297529658161436 lk2=6.94341207093607e-09 wk2=-1.11368360008786e-08 pk2=8.18937970663712e-15
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=132964.794328 lvsat=-0.0803030422661992 wvsat=0.329890093026259 pvsat=-3.11383258807486e-7
+  ua=3.74672845161647e-09 lua=-1.81513619374303e-15 wua=-1.32996922913796e-15 pua=5.01127761394403e-22
+  ub=-1.67265680973944e-19 lub=7.24925019027302e-25 wub=2.48070049234618e-24 pub=-2.46055051109675e-30
+  uc=5.52615694e-13 luc=-1.0742296475666e-18
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0268496320149365 lu0=-6.65673991638746e-09 wu0=-4.68899981095172e-09 pu0=-4.2752921434267e-15
+  a0=1.78673210393568 la0=-1.46449793931181e-06 wa0=-4.94342516032994e-06 pa0=8.59821969778593e-12
+  keta=0.0466423328 lketa=-1.2394759872992e-07 pketa=-2.01948391736579e-28
+  a1=0.0
+  a2=0.5
+  ags=-0.399217885736026 lags=1.20139452309976e-06 wags=8.88841075646897e-07 pags=-1.96755919425498e-12
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.1606776136623+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=7.82699159621449e-8
+  nfactor={1.32407918772759+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.04854507548014e-07 wnfactor=-2.59701030183664e-06 pnfactor=3.34883353349686e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.47195e-05 lcit=-9.17423605e-12
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.280615734987127 leta0=-2.65956107241476e-07 weta0=-7.75888782611441e-09 peta0=1.50825020451841e-14
+  etab=-0.0293684412 letab=2.772087164868e-8
+  dsub=-0.512031344112724 ldsub=1.56519201482072e-06 wdsub=3.92725107062253e-06 pdsub=-7.63418335618313e-12
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.0417844962480007 lpclm=1.09617750274151e-6
+  pdiblc1=-0.00906932781999981 lpdiblc1=3.85673507489298e-7
+  pdiblc2=0.00602058784087 lpdiblc2=-4.26114512466719e-9
+  pdiblcb=-0.41378 lpdiblcb=3.66969442e-7
+  drout=1.556250265901 ldrout=-1.08129489188495e-6
+  pscbe1=433349461.692 lpscbe1=-126.359101721079
+  pscbe2=1.45323618864e-08 lpscbe2=2.09612945270314e-17
+  pvag=0.0
+  delta=0.01
+  alpha0=-6.40086482779e-05 lalpha0=1.2442660577741e-10 walpha0=4.5360685341566e-26 palpha0=-1.70934181886405e-31
+  alpha1=1.9439e-10 lalpha1=-1.83484721e-16
+  beta0=-41.5076459075 lbeta0=8.65184128795893e-05 wbeta0=1.35525271560688e-20 pbeta0=-5.16987882845642e-26
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-3.81344931588543e-09 lagidl=9.32816169363699e-15 wagidl=6.83625352702166e-14 pagidl=-4.96718574449701e-20
+  bgidl=487643931.174281 lbgidl=1423.82135219032 wbgidl=2003.91201588643 pbgidl=-0.00389540456768165
+  cgidl=563.459145 lcgidl=-0.0001844938869655
+  egidl=3.152521570876 legidl=-2.24038668162586e-6
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.455913102428 lkt1=-1.64320622618211e-07 wkt1=-3.29890093026258e-07 pkt1=3.11383258807485e-13
+  kt2=-0.019032
+  at=484396.7488312 lat=-0.42890509122177 wat=-1.51749442792079 pat=1.43236299051443e-6
+  ute=-1.10489856009144 lute=-3.35935369129691e-07 wute=-1.64285266327077e-06 pute=1.55068862886128e-12
+  ua1=5.524e-10
+  ub1=-4.07319781456696e-18 lub1=4.55240907169754e-25 wub1=2.36861086792855e-24 pub1=-2.23573179823776e-30
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=2.81e-6
+  sbref=2.81e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.37 pmos
* DC IV MOS Parameters
+  lmin=8.0e-07 lmax=1e-06 wmin=5.0e-06 wmax=7.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.761893802395491+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-2.11935869204932e-07 wvth0=-2.00070282965225e-06 pvth0=1.57930671100782e-12
+  k1=0.590771669999999 lk1=-1.07431583129997e-8
+  k2=0.032667510137854 lk2=4.19237368567356e-09 wk2=-1.75468555754145e-08 pk2=1.42397971830409e-14
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=8738.12288046454 lvsat=0.0369545129131293 wvsat=-0.00638162194157221 pvsat=6.02361295065062e-9
+  ua=-3.17634227606689e-10 lua=2.02121573917572e-15 wua=-3.86627564122e-15 pua=2.89514738375865e-21
+  ub=3.20612872144498e-18 lub=-2.45922195741592e-24 wub=2.40320265874442e-24 pub=-2.38740030596004e-30
+  uc=6.40846463e-12 luc=-6.601565458257e-18 wuc=-6.16297582203915e-33
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0145595834606626 lu0=4.94383691399157e-09 wu0=-5.6898777661066e-09 pu0=-3.33056344155617e-15
+  a0=-2.02744297703456 la0=2.13570191961601e-06 wa0=1.96606034447525e-05 pa0=-1.46255229025514e-11
+  keta=-0.157135299 lketa=6.83981079261002e-8
+  a1=0.0
+  a2=0.5
+  ags=1.44065796376763 lags=-5.35264291246741e-07 wags=-5.64291051475934e-06 pags=4.19776113192948e-12
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.0961094772140001+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=1.73240519685946e-8
+  nfactor={1.79811171336607+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-3.42584793402147e-07 wnfactor=-1.01088004492763e-08 pnfactor=9.07057206337322e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-1.35975e-05 lcit=1.755418025e-11
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.000352821377956578 leta0=-1.41594308577994e-09 weta0=-2.5279200615028e-09 peta0=1.0144991572167e-14
+  etab=-0.0021235300373519 letab=2.00440000225646e-09 wetab=2.0145347602897e-08 petab=-1.90151936023745e-14
+  dsub=4.38726721383548 ldsub=-3.05925589402658e-06 wdsub=-1.9636476910907e-05 pdsub=1.46076194855826e-11
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=2.061963089575 lpclm=-8.10669071499842e-7
+  pdiblc1=0.185912130255001 lpdiblc1=2.01630509212306e-7
+  pdiblc2=-0.03533450056535 lpdiblc2=3.47739228219639e-08 wpdiblc2=-2.64697796016969e-23 ppdiblc2=1.26217744835362e-29
+  pdiblcb=-0.025
+  drout=0.332185866169999 ldrout=7.40994950211371e-8
+  pscbe1=-74402724.1500006 lpscbe1=352.908186495185
+  pscbe2=1.8463592403e-08 lpscbe2=-3.68972719009169e-15
+  pvag=0.0
+  delta=0.01
+  alpha0=0.000255919397305 lalpha0=-1.77553476448289e-10
+  alpha1=0.0
+  beta0=68.0295673024999 lbeta0=-1.68737626693297e-5
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=3.52169284838196e-08 lagidl=-2.75126119115046e-14 wagidl=-2.63171865811791e-13 pagidl=2.63263463736337e-19
+  bgidl=2698289944.1286 lbgidl=-662.807419437268 wbgidl=-10019.5600794322 pbgidl=0.00745355074308961
+  cgidl=-197.364 lcgidl=0.000533647079599999
+  egidl=1.887175135705 legidl=-1.04602618146795e-6
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.552386517642001 lkt1=-7.32593659977181e-08 wkt1=-1.89365636248445e-07 pkt1=1.78742224054907e-13
+  kt2=-0.019032
+  at=48597.4999999999 lat=-0.01755418025
+  ute=-1.3901295 lute=-6.67058849499986e-8
+  ua1=5.524e-10
+  ub1=-3.5909e-18
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=2.41e-6
+  sbref=2.41e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.38 pmos
* DC IV MOS Parameters
+  lmin=6e-07 lmax=8.0e-07 wmin=5.0e-06 wmax=7.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.0271332345347+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-1.46242556365752e-08 wvth0=4.54919380147513e-07 pvth0=-2.4743065086224e-13
+  k1=0.595611255 lk1=-1.43433255945006e-8
+  k2=0.034428376386116 lk2=2.88246528359153e-09 wk2=5.93345660245138e-09 pk2=-3.22720704607327e-15
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=60745.0316195354 lvsat=-0.00173342649786534 wvsat=0.00638162194157266 pvsat=-3.4709641740214e-9
+  ua=-2.2486138494545e-09 lua=3.45767147986831e-15 wua=9.51246712754585e-17 pua=-5.1738308706721e-23
+  ub=3.030596887635e-18 lub=-2.32864382624468e-24 wub=-2.99828924060037e-24 pub=1.63076951796254e-30
+  uc=3.1396334e-12 luc=-4.16988190626e-18
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0112934363518926 lu0=7.37352374820563e-09 wu0=-3.78163175588142e-08 pu0=2.0568295120239e-14
+  a0=0.945572834999998 la0=-7.59245429564991e-8
+  keta=0.0210589425000002 lketa=-6.41605883257501e-8
+  a1=0.0
+  a2=0.5
+  ags=-0.717169160000001 lags=1.069943306124e-6
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={0.0170483782755001+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=-6.68540767300446e-8
+  nfactor={1.36962857285435+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-2.38361851754832e-08 wnfactor=4.49768634841556e-06 pnfactor=-2.44629160490322e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=-0.0702494608135902 leta0=5.11050946365117e-08 weta0=4.13223591920756e-08 peta0=-2.24752311645699e-14
+  etab=0.0021235300373519 letab=-1.1549879873157e-09 wetab=-2.0145347602897e-08 petab=1.09570545612157e-14
+  dsub=0.183470231958141 ldsub=6.79486807919671e-08 wdsub=2.21557794409088e-10 pdsub=-1.2050528437881e-16
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.170632713424999 lpclm=5.96291595318144e-7
+  pdiblc1=0.157259843574999 lpdiblc1=2.22944945273557e-7
+  pdiblc2=0.0277574173458 lpdiblc2=-1.21601549121406e-8
+  pdiblcb=-0.025
+  drout=-0.81794092163 ldrout=9.29678812465557e-7
+  pscbe1=434417012.98 lpscbe1=-25.6028159558223
+  pscbe2=1.03443636915e-08 lpscbe2=2.35016704839314e-15
+  pvag=0.0
+  delta=0.01
+  alpha0=-0.0001310877634225 lalpha0=1.10341150416898e-10
+  alpha1=0.0
+  beta0=25.181273087 lbeta0=1.50010833975807e-5
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-2.4307825511956e-08 lagidl=1.67678525859529e-14 wagidl=3.37449563794728e-13 pagidl=-1.83538817747952e-19
+  bgidl=2079521950.0 lbgidl=-202.505908604999
+  cgidl=1308.655 lcgidl=-0.0005866804545
+  egidl=-0.2962646614 legidl=5.7823468359846e-7
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.738942122357999 lkt1=6.55193483505157e-08 wkt1=1.89365636248445e-07 pkt1=-1.02995969555526e-13
+  kt2=-0.019032
+  at=44036.5 lat=-0.01416125235
+  ute=-1.62257375 lute=1.06209392624999e-7
+  ua1=5.53487799999999e-10 lua1=-8.09214420000522e-19
+  ub1=-4.38417814999999e-18 lub1=5.90119615784998e-25
+  uc1=-2.93321028e-10 luc1=1.369676327292e-16
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=2.02e-6
+  sbref=2.01e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.39 pmos
* DC IV MOS Parameters
+  lmin=5e-07 lmax=6e-07 wmin=5.0e-06 wmax=7.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.15137648365926+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=5.29516475622704e-08 wvth0=9.38262222401463e-07 pvth0=-5.10320822764163e-13
+  k1=0.314191727734757 lk1=1.38720755285064e-07 wk1=8.79126466112013e-07 pk1=-4.78156884918326e-13
+  k2=0.063100745589908 lk2=-1.2712436326351e-08 wk2=-4.43706502604944e-08 pk2=2.41331966766832e-14
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=108473.246047856 lvsat=-0.027692802325429 wvsat=-0.487677892345271 pvsat=2.65248005646593e-7
+  ua=1.92378105691265e-08 lua=-8.22879476139792e-15 wua=-4.64326500499605e-14 pua=2.52547183621735e-20
+  ub=-1.08092166002109e-17 lub=5.1988307297947e-24 wub=1.0474185419727e-23 pub=-5.6969094497895e-30
+  uc=-5.09501653292663e-11 luc=2.52495596225879e-17 wuc=3.43981771170579e-16 puc=-1.87091685339678e-22
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0695970451097486 lu0=-2.43378090551923e-08 wu0=-1.71013073971739e-07 pu0=9.3014010933229e-14
+  a0=-1.62897429535331 la0=1.32437164124267e-06 wa0=1.21141668393721e-05 pa0=-6.58889534393448e-12
+  keta=-0.034424149148728 lketa=-3.39833347780067e-08 wketa=-7.70346807408862e-07 pketa=4.18991628549679e-13
+  a1=0.0
+  a2=0.5
+  ags=1.25
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.467566684982424+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=1.96728056175941e-07 wvoff=2.36686909609425e-06 pvoff=-1.28734010136566e-12
+  nfactor={-1.48489212547227+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.52873762264437e-06 wnfactor=1.38603666238174e-05 pnfactor=-7.53865340669428e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=3.2195e-05 lcit=-1.20718605e-11
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=-0.659442270580415 leta0=3.71567063868688e-07 weta0=2.99279659346169e-06 peta0=-1.62778206718381e-12
+  etab=-0.0524374809785162 letab=2.8520745904215e-08 wetab=4.80521335851643e-07 petab=-2.61355554569709e-13
+  dsub=0.553855835700348 ldsub=-1.33504049083419e-07 wdsub=-8.15022552972508e-07 pdsub=4.43290766561747e-13
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-0.703946769493438 lpclm=1.07197537607748e-06 wpclm=1.1483644079414e-05 ppclm=-6.24595401479328e-12
+  pdiblc1=2.85501663826025 lpdiblc1=-1.24436497535575e-06 wpdiblc1=-7.43241086026637e-06 ppdiblc1=4.04248826689887e-12
+  pdiblc2=0.0425955558920985 lpdiblc2=-2.02306184674724e-08 wpdiblc2=-2.38679053874295e-07 ppdiblc2=1.29817537402229e-13
+  pdiblcb=-0.025
+  drout=-1.07400900603912 ldrout=1.06895424357567e-06 wdrout=1.3329236380408e-05 pdrout=-7.2497716673039e-12
+  pscbe1=5877345.72951794 lpscbe1=207.479909061715 wpscbe1=3394.2455132761 ppscbe1=-0.00184613013467087
+  pscbe2=1.51583479493027e-08 lpscbe2=-2.68158989425747e-16 wpscbe2=2.0714087779504e-15 ppscbe2=-1.12663923432726e-21
+  pvag=0.0
+  delta=0.01
+  alpha0=-0.000619055863127569 lalpha0=3.75746999846485e-10 walpha0=3.99666748917066e-09 palpha0=-2.17378744735992e-15
+  alpha1=0.0
+  beta0=-1.013647840614 lbeta0=2.92485008901098e-05 wbeta0=0.000312664077297074 pbeta0=-1.70057991641878e-10
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.82131753824793e-09 lagidl=3.80611680946946e-16 wagidl=-1.08026336966977e-13 pagidl=5.87555246763388e-20
+  bgidl=3622210349.75119 lbgidl=-1041.57412922968 wbgidl=-8633.06709652412 pbgidl=0.00469552519379945
+  cgidl=2942.02413127199 lcgidl=-0.00147506992499884 wcgidl=-0.0170250712374734 pcgidl=9.25993624606176e-9
+  egidl=1.3165878293526 legidl=-2.98995786121878e-07 wegidl=-6.82488399962662e-07 pegidl=3.71205440739691e-13
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.467061448559999 lkt1=-8.23565501282158e-08 wkt1=-1.50664347234277e-06 pkt1=8.19463384607236e-13
+  kt2=-0.019032
+  at=18000.0
+  ute=-1.67100109999999 lute=1.32549028289999e-7
+  ua1=5.52e-10
+  ub1=-1.6356839137848e-17 lub1=7.10204992707552e-24 wub1=5.52938154349799e-23 pub1=-3.00743062150856e-29
+  uc1=-4.1496e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=1.81e-6
+  sbref=1.81e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.40 pmos
* DC IV MOS Parameters
+  lmin=2.0e-05 lmax=1.0e-04 wmin=3.0e-06 wmax=5.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.067493945512+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} wvth0=9.36003110681999e-8
+  k1=0.59521
+  k2=0.0309593236852 wk2=-8.07690480189101e-9
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=200000.0
+  ua=2.691214109728e-09 wua=1.24838539216062e-16
+  ub=-3.275957242e-19 wub=-6.85168001824277e-25
+  uc=-3.9972e-11
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0214165256424 wu0=-5.17396556828806e-9
+  a0=0.92049813754 wa0=-2.7556835128144e-8
+  keta=-0.0079259
+  a1=0.0
+  a2=0.5
+  ags=0.1193262716044 wags=4.35669631791178e-8
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.093204657+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.76605404104+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} wnfactor=-1.71417096335381e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.08353125
+  pdiblc1=0.39
+  pdiblc2=0.0029407877
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=333712830.0
+  pscbe2=1.5000958e-8
+  pvag=0.0
+  delta=0.01
+  alpha0=5.0667189e-5
+  alpha1=0.0
+  beta0=38.266046
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=1.6226228868e-08 wagidl=-4.22466655271931e-15
+  bgidl=1601356092.0 wbgidl=507.531853203167
+  cgidl=1000.0
+  egidl=0.69350825
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.576
+  kt2=-0.019032
+  at=448800.0
+  ute=-1.5361
+  ua1=2.2096e-11
+  ub1=-3.6627e-18
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.41 pmos
* DC IV MOS Parameters
+  lmin=8e-06 lmax=2.0e-05 wmin=3.0e-06 wmax=5.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.067493945512+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} wvth0=9.36003110681999e-8
+  k1=0.59521
+  k2=0.0309593236852 wk2=-8.07690480189101e-9
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=200000.0
+  ua=2.691214109728e-09 wua=1.24838539216055e-16
+  ub=-3.275957242e-19 wub=-6.85168001824277e-25
+  uc=-3.9972e-11
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0214165256424 wu0=-5.17396556828806e-9
+  a0=0.92049813754 wa0=-2.7556835128144e-8
+  keta=-0.0079259
+  a1=0.0
+  a2=0.5
+  ags=0.1193262716044 wags=4.35669631791178e-8
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.093204657+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.76605404104+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} wnfactor=-1.71417096335378e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.08353125
+  pdiblc1=0.39
+  pdiblc2=0.0029407877
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=333712830.0
+  pscbe2=1.5000958e-8
+  pvag=0.0
+  delta=0.01
+  alpha0=5.0667189e-5
+  alpha1=0.0
+  beta0=38.266046
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=1.6226228868e-08 wagidl=-4.22466655271931e-15
+  bgidl=1601356092 wbgidl=507.531853203167
+  cgidl=1000.0
+  egidl=0.69350825
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.576
+  kt2=-0.019032
+  at=448800.0
+  ute=-1.5361
+  ua1=2.2096e-11
+  ub1=-3.6627e-18
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.42 pmos
* DC IV MOS Parameters
+  lmin=4e-06 lmax=8e-06 wmin=3.0e-06 wmax=5.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.06884109636262+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=1.07016316422427e-08 wvth0=8.1104064255246e-08 pvth0=9.92689350574326e-14
+  k1=0.60423167125 lk1=-7.16672542428762e-8
+  k2=0.0300897401552974 lk2=6.90788460319344e-09 wk2=-8.72744263654154e-09 pk2=5.16780750468094e-15
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=274036.86275 lvsat=-0.588141433999725
+  ua=2.40539279702907e-09 lua=2.27053592594906e-15 wua=2.74295906484747e-16 pua=-1.18727437984573e-21
+  ub=-1.84018288117508e-19 lub=-1.14056479449571e-24 wub=-2.93576646535144e-25 pub=-3.11076256728134e-30
+  uc=-5.1678481175e-11 luc=9.29951158060826e-17
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0201430880117847 lu0=1.01160611938452e-08 wu0=-3.59660514147549e-09 pu0=-1.25303934945565e-14
+  a0=0.940857490480744 la0=-1.61732663825988e-07 wa0=-2.85153740827762e-08 pa0=7.61453760170282e-15
+  keta=-0.00493040935249999 lketa=-2.37958781546752e-8
+  a1=0.0
+  a2=0.5
+  ags=0.0951173151486372 lags=1.92313529188934e-07 wags=7.04631433612426e-08 pags=-2.13660565748783e-13
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.0947904104522501+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=1.25970668493289e-8
+  nfactor={1.92167410284978+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.23623020901072e-06 wnfactor=-5.74355861308013e-07 pnfactor=3.20090525506613e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-0.6548060915245 lpclm=5.86527800733647e-06 wpclm=-2.11758236813575e-22 ppclm=-1.61558713389263e-27
+  pdiblc1=0.39
+  pdiblc2=0.0045684231025075 lpdiblc2=-1.29297728739793e-8
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=564147837.55925 lpscbe1=-1830.55265654993
+  pscbe2=-1.558611817795e-08 lpscbe2=2.42980674450017e-13 ppscbe2=-9.62964972193618e-35
+  pvag=0.0
+  delta=0.01
+  alpha0=7.83968484975e-05 lalpha0=-2.2028164208219e-10
+  alpha1=0.0
+  beta0=39.148037118575 lbeta0=-7.00644924684789e-6
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=2.65980677208335e-08 lagidl=-8.2392850663024e-14 wagidl=-1.89903953023725e-14 pagidl=1.1729747261437e-19
+  bgidl=1344564909.8097 lbgidl=2039.92347220152 wbgidl=1007.94557216516 pbgidl=-0.00397523654206218
+  cgidl=1335.2315 lcgidl=-0.00266304551285 wcgidl=-1.73472347597681e-18
+  egidl=1.21389074000325 legidl=-4.13386646233682e-6
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.576
+  kt2=-0.019032
+  at=650243.063506628 lat=-1.6002435521903 wat=0.0425704065145132 pat=-3.38175052310642e-7
+  ute=-1.5163805 lute=-1.5664973605e-7
+  ua1=2.2096e-11
+  ub1=-3.2752784729661e-18 lub1=-3.0776378686046e-24 wub1=-8.66913907497545e-25 pub1=6.8866773897697e-30
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.43 pmos
* DC IV MOS Parameters
+  lmin=2e-06 lmax=4e-06 wmin=3.0e-06 wmax=5.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.04482593828968+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-8.40117502816181e-08 wvth0=9.11836345289863e-08 pvth0=5.95161178548223e-14
+  k1=0.602894174 lk1=-6.63922988385996e-8
+  k2=0.0290042682041359 lk2=1.1188877431379e-08 wk2=-1.04526295966402e-09 pk2=-2.51299409229566e-14
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=137793.663786 lvsat=-0.0508118816056053 wvsat=-0.0694782513691294 pvsat=2.7401527557471e-7
+  ua=3.44586706484229e-09 lua=-1.83299053887953e-15 wua=-4.90595485953602e-16 pua=1.82938078279188e-21
+  ub=-1.6011320641667e-18 lub=4.4483902268647e-24 wub=-1.01632520899498e-24 pub=-2.60314511795978e-31
+  uc=-5.540982305e-11 luc=1.07711155026895e-16
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0225533225446134 lu0=6.10337219821866e-10 wu0=-9.32549089430616e-09 pu0=1.00637590260323e-14
+  a0=0.917652238179403 la0=-7.02134692747201e-08 wa0=-2.71452420997834e-07 pa0=9.65733956929998e-13
+  keta=-0.00498067579999999 lketa=-2.359763231238e-8
+  a1=0.0
+  a2=0.5
+  ags=0.104824129108753 lags=1.54030825611631e-07 wags=-1.38980175525042e-08 pags=1.19051416778944e-13
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.06358776784865+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=-1.10463035315009e-7
+  nfactor={1.95241773720061+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.35748002852696e-06 wnfactor=7.26039716739547e-07 pnfactor=-1.92772486519564e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.01798959 leta0=2.44562855999e-7
+  etab=-0.1233522794 letab=2.1041605472566e-7
+  dsub=0.8193648575 ldsub=-1.02290906149425e-6
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=1.0526917789172 lpclm=-8.68922843898544e-07 wpclm=5.69721661239028e-12 ppclm=-2.24692525980959e-17
+  pdiblc1=0.58503867943 lpdiblc1=-7.69213047803978e-7
+  pdiblc2=-0.0011773222896 lpdiblc2=9.73087237795344e-9
+  pdiblcb=0.16939 lpdiblcb=-7.66654721e-07 ppdiblcb=-2.01948391736579e-28
+  drout=0.132342 ldrout=1.6866403862e-6
+  pscbe1=-160819458.431 lpscbe1=1028.64586210602 ppscbe1=-4.33680868994202e-19
+  pscbe2=7.662008170125e-08 lpscbe2=-1.2067135725356e-13
+  pvag=0.0
+  delta=0.01
+  alpha0=4.445374715855e-05 lalpha0=-8.64134447115054e-11
+  alpha1=-9.7195e-11 lalpha1=3.833273605e-16
+  beta0=70.77889717255 lbeta0=-0.00013175539821372
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=1.27452823570094e-09 lagidl=1.74806567123903e-14 wagidl=2.38970772263074e-14 pagidl=-5.18464302914908e-20
+  bgidl=2485500315.0 lbgidl=-2459.8116723285
+  cgidl=846.079827500001 lcgidl=-0.00073388023167725
+  egidl=-1.617101386419 legidl=7.0312833850599e-06 wegidl=-4.2351647362715e-22 pegidl=2.42338070083895e-27
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.57697195 lkt1=3.83327360499981e-9
+  kt2=-0.019032
+  at=474951.874461442 lat=-0.908912631714993 wat=-0.55015874944261 pat=1.99948946586866e-6
+  ute=-1.659418285 lute=4.074769842115e-7
+  ua1=-4.933329728e-10 lua1=2.03280032582592e-15 wua1=9.86076131526265e-32 pua1=1.41059322098675e-36
+  ub1=-5.25840384761654e-18 lub1=4.74361029647927e-24 wub1=5.42242818018216e-24 pub1=-1.79178588698303e-29
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.44 pmos
* DC IV MOS Parameters
+  lmin=1e-06 lmax=2e-06 wmin=3.0e-06 wmax=5.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.06293228527081+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-4.88148223849926e-08 wvth0=-4.84612329469418e-08 pvth0=3.30971775741277e-13
+  k1=0.558687465 lk1=1.95411227865e-8
+  k2=0.0307358477030981 lk2=7.82286004334646e-09 wk2=-1.59638633043733e-08 pk2=3.87032628712393e-15
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=171842.794328 lvsat=-0.116999986466199 wvsat=0.138956502738259 pvsat=-1.31161042934643e-7
+  ua=3.36042486593186e-09 lua=-1.66689944841753e-15 wua=5.67204765303407e-16 pua=-2.26877125626624e-22
+  ub=6.41490862171316e-19 lub=8.8955520356231e-26 wub=-1.49118053166833e-24 pub=6.62756749948748e-31
+  uc=5.52615694e-13 luc=-1.0742296475666e-18
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0268154335725901 lu0=-7.67478040746212e-09 wu0=-4.52104797753868e-09 pu0=7.24402440128015e-16
+  a0=0.398878799642588 la0=9.38230217896995e-07 wa0=1.87245565097067e-06 pa0=-3.20180894416958e-12
+  keta=0.0466423328 lketa=-1.2394759872992e-07 pketa=-2.52435489670724e-29
+  a1=0.0
+  a2=0.5
+  ags=-0.152780981174146 lags=6.54789399490559e-07 wags=-3.21434220599336e-07 pags=7.16871041881681e-13
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.1606776136623+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=7.8269915962145e-8
+  nfactor={0.820500085300985+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=8.42854695000723e-07 wnfactor=-1.2388498622576e-07 pnfactor=-2.75556235101388e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.47195e-05 lcit=-9.17423605000001e-12
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.290368288598006 leta0=-2.84914096205664e-07 weta0=-5.56546148542895e-08 peta0=1.08187005815254e-13
+  etab=-0.0293684412 letab=2.772087164868e-8
+  dsub=0.287636937054122 ldsub=1.07168430604934e-08 wdsub=3.37365715638376e-12 pdsub=-6.55805214579416e-18
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.0417868163886008 lpclm=1.0961753127608e-06 wpclm=-1.13944332247806e-11 ppclm=1.07552055200395e-17
+  pdiblc1=-0.00906932782000014 lpdiblc1=3.85673507489298e-7
+  pdiblc2=0.00602058784087 lpdiblc2=-4.2611451246672e-9
+  pdiblcb=-0.41378 lpdiblcb=3.66969442e-7
+  drout=1.556250265901 ldrout=-1.08129489188495e-06 pdrout=-1.61558713389263e-27
+  pscbe1=433349461.692 lpscbe1=-126.359101721079
+  pscbe2=1.45323618864e-08 lpscbe2=2.0961294527044e-17
+  pvag=0.0
+  delta=0.01
+  alpha0=-6.40086482779e-05 lalpha0=1.2442660577741e-10 walpha0=-9.36496223633124e-27 palpha0=2.09860536254563e-32
+  alpha1=1.9439e-10 lalpha1=-1.83484721e-16
+  beta0=-41.5076459075 lbeta0=8.65184128795893e-05 pbeta0=-2.58493941422821e-26
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=6.72660953635165e-09 lagidl=6.88235587205537e-15 wagidl=1.65992944012306e-14 pagidl=-3.76602702578239e-20
+  bgidl=895681570.0 lbgidl=630.636986077001
+  cgidl=1321.8473949744 lcgidl=-0.00165872480609074 wcgidl=-0.00372451750089628 pcgidl=7.24008956999227e-9
+  egidl=3.152521570876 legidl=-2.24038668162586e-06 pegidl=-3.23117426778526e-27
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.5230855 lkt1=-1.0091659655e-7
+  kt2=-0.019032
+  at=-13970.6829493959 lat=0.0415039276359349 wat=0.930035872827167 pat=-8.77860860361563e-7
+  ute=-1.4394171 lute=-2.01833193100009e-8
+  ua1=5.524e-10
+  ub1=-2.08875043290252e-18 lub1=-1.41787897638331e-24 wub1=-7.37720073037417e-24 pub1=6.96333976940018e-30
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=2.81e-6
+  sbref=2.81e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.45 pmos
* DC IV MOS Parameters
+  lmin=8.0e-07 lmax=1e-06 wmin=3.0e-06 wmax=5.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.45967061626058+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=3.25666488236245e-07 wvth0=1.4261460898133e-06 pvth0=-1.06091007621211e-12
+  k1=0.59077167 lk1=-1.07431583129997e-8
+  k2=0.0404952874515038 lk2=-1.38907513517361e-09 wk2=-5.59898214293701e-08 pk2=4.16508281613085e-14
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=7438.69360000012 lvsat=0.03818104421096
+  ua=-1.41897961017227e-09 lua=2.84438043657716e-15 wua=1.54253726171631e-15 pua=-1.14749346899076e-21
+  ub=4.45372099579868e-18 lub=-3.50940850277464e-24 wub=-3.72384276946495e-24 pub=2.77016663620498e-30
+  uc=6.40846463e-12 luc=-6.601565458257e-18 wuc=-3.08148791101958e-33 puc=-2.93873587705572e-39
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0170081603085286 lu0=1.58230482648555e-09 wu0=-1.77150737293536e-08 pu0=1.31782433472661e-14
+  a0=3.43622413939817 la0=-1.9287200482983e-06 wa0=-7.17199027609182e-06 pa0=5.3352435663847e-12
+  keta=-0.157135299 lketa=6.83981079260999e-8
+  a1=0.0
+  a2=0.5
+  ags=-0.129308683198584 lags=6.32633897431426e-07 wags=2.06734640528983e-06 pags=-1.53789899089511e-12
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.0961094772139999+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=1.73240519685946e-8
+  nfactor={2.19564977158162+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-4.55149093879564e-07 wnfactor=-1.96245636799941e-06 pnfactor=1.45987129215477e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-1.35975e-05 lcit=1.755418025e-11
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=-0.0568240276050302 leta0=4.2800731058382e-08 weta0=2.78273074271448e-07 peta0=-2.0700733995053e-13
+  etab=0.00197847644 letab=-1.867483911716e-9
+  dsub=0.388880694284393 ldsub=-8.48471393891596e-08 wdsub=-1.68682857819188e-11 pdsub=1.25483177932974e-17
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=2.061963089575 lpclm=-8.10669071499841e-7
+  pdiblc1=0.185912130255 lpdiblc1=2.01630509212305e-7
+  pdiblc2=-0.03533450056535 lpdiblc2=3.47739228219639e-08 wpdiblc2=2.64697796016969e-23
+  pdiblcb=-0.025
+  drout=0.33218586617 ldrout=7.40994950211371e-8
+  pscbe1=-74402724.1499996 lpscbe1=352.908186495185
+  pscbe2=1.8463592403e-08 lpscbe2=-3.68972719009171e-15
+  pvag=0.0
+  delta=0.01
+  alpha0=0.000255919397305 lalpha0=-1.7755347644829e-10
+  alpha1=0.0
+  beta0=68.0295673025 lbeta0=-1.68737626693297e-5
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=4.02004606708838e-09 lagidl=9.43708113069296e-15 wagidl=-1.09960981362512e-13 pagidl=8.17999740355726e-20
+  bgidl=658101750.0 lbgidl=854.888578175
+  cgidl=-3989.305249872 lcgidl=0.00335447217537978 wcgidl=0.0186225875044814 pcgidl=-1.38533428445837e-8
+  egidl=1.887175135705 legidl=-1.04602618146795e-6
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.59094525 lkt1=-3.68637785249996e-8
+  kt2=-0.019032
+  at=48597.5 lat=-0.01755418025
+  ute=-1.3901295 lute=-6.67058849500003e-8
+  ua1=5.524e-10
+  ub1=-3.5909e-18
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=2.41e-6
+  sbref=2.41e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.46 pmos
* DC IV MOS Parameters
+  lmin=6e-07 lmax=8.0e-07 wmin=3.0e-06 wmax=5.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.794510848210322+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-1.69145863216341e-07 wvth0=-6.87511490840597e-07 pvth0=5.11439798036319e-13
+  k1=0.623676047152739 lk1=-3.52207244769235e-08 wk1=-1.37828888482153e-07 pk1=1.02530910141875e-13
+  k2=0.035106129386676 lk2=2.61991954925172e-09 wk2=2.604946552413e-09 pk2=-1.93781974034011e-15
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=134889.815414479 lvsat=-0.0566298453068312 wvsat=-0.357750529174642 pvsat=2.66130618653016e-7
+  ua=-8.98940456267072e-09 lua=8.47601955874075e-15 wua=3.31997949797888e-14 pua=-2.46973274854649e-20
+  ub=5.49088409895426e-18 lub=-4.28095413521208e-24 wub=-1.50809959229616e-23 pub=1.12187528670911e-29
+  uc=1.12986107745032e-11 luc=-1.02393451751529e-17 wuc=-4.00695211480132e-17 puc=2.9807716782007e-23
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=-0.0229725026656818 lu0=3.13239200130007e-08 wu0=1.30466998486639e-07 pu0=-9.70544001742109e-14
+  a0=1.09413019035858 la0=-1.86436359607747e-07 wa0=-7.295794336721e-07 pa0=5.42734140708675e-13
+  keta=0.23433552940968 lketa=-2.22817041327861e-07 wketa=-1.04742179286578e-06 pketa=7.79177071712855e-13
+  a1=0.0
+  a2=0.5
+  ags=-2.81066807025968 lags=2.62729714546618e-06 wags=1.02813741241807e-05 pags=-7.64831421097801e-12
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={0.147858053872035+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=-1.64163394406307e-07 wvoff=-6.42418874583443e-07 pvoff=4.77895400802623e-13
+  nfactor={3.11295353513887+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.13753136358981e-06 wnfactor=-4.06394990056009e-06 pnfactor=3.02317233102665e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=-0.154734473195029 leta0=1.15636311532782e-07 weta0=4.5623636555851e-07 peta0=-3.39394232338976e-13
+  etab=-0.00197847644 letab=1.076093335716e-9
+  dsub=0.050598035854696 ldsub=1.66801330216692e-07 wdsub=6.52769668589256e-07 pdsub=-4.85595356463547e-13
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-0.996088780204323 lpclm=1.46421571442899e-06 wpclm=5.72988126047699e-06 ppclm=-4.26245866966883e-12
+  pdiblc1=-0.278964204284975 lpdiblc1=5.47452014476593e-07 wpdiblc1=2.14233817654894e-06 ppdiblc1=-1.59368536953475e-12
+  pdiblc2=0.0515505201311965 lpdiblc2=-2.98598440741971e-08 wpdiblc2=-1.1685021191695e-07 ppdiblc2=8.69248726450188e-14
+  pdiblcb=-0.025
+  drout=-2.6369920523285 ldrout=2.28287094859217e-06 wdrout=8.93353473176889e-06 pdrout=-6.64565648696288e-12
+  pscbe1=484512627.389013 lpscbe1=-62.8689435146869 wpscbe1=-246.024371541647 ppscbe1=0.000183017529989831
+  pscbe2=5.74592176791542e-09 lpscbe2=5.77094799534771e-15 wpscbe2=2.25833897371485e-14 ppscbe2=-1.67997836254647e-20
+  pvag=0.0
+  delta=0.01
+  alpha0=-0.000346986191715301 lalpha0=2.70947991223912e-10 walpha0=1.06029790759506e-09 palpha0=-7.88755613459967e-16
+  alpha1=0.0
+  beta0=-4.17051739180334 lbeta0=3.68358803347625e-05 wbeta0=0.000144149460813289 pbeta0=-1.07232783899006e-10
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=6.48800504056994e-08 lagidl=-3.58366760967998e-14 wagidl=-1.00560656872966e-13 pagidl=7.48070726477994e-20
+  bgidl=2475754064.8786 lbgidl=-497.262978863189 wbgidl=-1945.93395445184 pbgidl=0.00144758026871672
+  cgidl=2456.58020794 lcgidl=-0.00144062201668657 wcgidl=-0.0056375708970133 pcgidl=4.1937889902882e-9
+  egidl=-1.42766449638101 legidl=1.41988302084083e-06 wegidl=5.55641320397588e-06 pegidl=-4.13341578243766e-12
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.807259185222 lkt1=1.24052157886645e-07 wkt1=5.24877290411585e-07 pkt1=-3.90456216337177e-13
+  kt2=-0.019032
+  at=44036.5 lat=-0.01416125235
+  ute=-1.74132463358 lute=1.94548174920162e-07 wute=5.83196989346206e-07 pute=-4.33840240374643e-13
+  ua1=5.534878e-10 lua1=-8.09214420000127e-19
+  ub1=-4.38417815e-18 lub1=5.90119615785001e-25
+  uc1=-2.93321028e-10 luc1=1.369676327292e-16
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=2.02e-6
+  sbref=2.01e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.47 pmos
* DC IV MOS Parameters
+  lmin=5e-07 lmax=6e-07 wmin=3.0e-06 wmax=5.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.1686037948853+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=3.43232904801773e-08 wvth0=1.02286720165441e-06 pvth0=-4.18835172811714e-13
+  k1=0.32315978510016 lk1=1.28230070453475e-07 wk1=8.35083475457027e-07 pk1=-4.26636124604646e-13
+  k2=0.0736703908582881 lk2=-1.83551822651581e-08 wk2=-9.6279192859455e-08 pk2=5.18452636857749e-14
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=366812.2049719 lvsat=-0.182772432987112 wvsat=-1.75640532016131 pvsat=1.02685895947066e-6
+  ua=2.23031054528687e-08 lua=-8.54397663871115e-15 wua=-6.14866074923271e-14 pua=2.6802606819119e-20
+  ub=-1.55265845692765e-17 lub=7.15044707343863e-24 wub=3.36416323831332e-23 pub=-1.52814846685939e-29
+  uc=-1.66201021665222e-10 luc=8.63027049088139e-17 wuc=9.09989790718668e-16 puc=-4.86929542942281e-22
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0766274493521475 lu0=-2.28484938894967e-08 wu0=-2.05540064124968e-07 pu0=8.5699841180242e-14
+  a0=1.3607214084968 la0=-3.31435323153127e-07 wa0=-2.56851577302341e-06 pa0=1.54293161568185e-12
+  keta=-0.134908216002467 lketa=-2.19853681981945e-08 wketa=-2.76859908619734e-07 pketa=3.6006846287143e-13
+  a1=0.0
+  a2=0.5
+  ags=-1.41185040580065 lags=1.86648021776691e-06 wags=1.30726028805259e-05 pags=-9.16646353155419e-12
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.166202722473177+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=6.6542618478538e-09 wvoff=8.86841745270929e-07 pvoff=-3.5386945033617e-13
+  nfactor={-2.00601446961707+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.64667533419695e-06 wnfactor=1.64196484836575e-05 pnfactor=-8.1178568301493e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=6.45008878600001e-05 lcit=-2.96430329070541e-11 wcit=-1.58657316645695e-10 pcit=8.62937145235935e-17
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.804308189527616 leta0=-4.05986992722065e-07 weta0=-4.19582243617302e-06 peta0=2.1908605499228e-12
+  etab=0.0138824456262119 letab=-7.55066217609668e-09 wetab=1.54817809582869e-07 petab=-8.42054066321225e-14
+  dsub=0.670927996690821 ldsub=-1.70596135482077e-07 wdsub=-1.38997517452419e-06 pdsub=6.25453563705853e-13
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.229997833001498 lpclm=7.97347205506351e-07 wpclm=6.89695247787957e-06 ppclm=-4.8972287048141e-12
+  pdiblc1=0.90013089329261 lpdiblc1=-9.3857809095856e-08 wpdiblc1=2.16822070230123e-06 ppdiblc1=-1.60776287529142e-12
+  pdiblc2=-0.0803444652744428 lpdiblc2=4.18778384879301e-08 wpdiblc2=3.65091192316621e-07 ppdiblc2=-1.7520305711762e-13
+  pdiblcb=-1.3172355144 lpdiblcb=7.02846896282162e-07 wpdiblcb=6.3462926658278e-06 ppdiblcb=-3.45174858094374e-12
+  drout=7.07010980622698 ldrout=-2.99682175227616e-06 wdrout=-2.66673129420368e-05 pdrout=1.271764456282e-11
+  pscbe1=924817293.808384 lpscbe1=-302.350651580183 wpscbe1=-1118.75678997422 ppscbe1=0.000657696692375307
+  pscbe2=2.53191834945908e-08 lpscbe2=-4.87494905779102e-15 wpscbe2=-4.78294300251717e-14 ppscbe2=2.14977490432612e-20
+  pvag=0.0
+  delta=0.01
+  alpha0=0.000341727301490559 lalpha0=-1.03643277730755e-10 walpha0=-7.2183086745277e-10 palpha0=1.80544227288549e-16
+  alpha1=6.46117757200002e-10 lalpha1=-3.51423448141081e-16 walpha1=-3.1731463329139e-15 palpha1=1.72587429047187e-21
+  beta0=-185.771106560767 lbeta0=0.000135608440783762 wbeta0=0.00122002569378778 pbeta0=-6.92401867013833e-10
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-2.69796382604468e-08 lagidl=1.41258085687171e-14 wagidl=5.30623058521697e-14 pagidl=-8.74845677840189e-21
+  bgidl=-1846637539.02961 lbgidl=1853.68581450248 wbgidl=18224.9698946758 pbgidl=-0.00952337433482378
+  cgidl=-440.053374803758 lcgidl=0.000134856988967765 wcgidl=-0.000415363925694757 pcgidl=1.35343061858804e-9
+  egidl=12.0058178737334 legidl=-5.8865880402644e-06 wegidl=-5.31783233140011e-05 pegidl=2.781240740969e-11
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.598860474987999 lkt1=1.07040993903732e-08 wkt1=-8.59365800848335e-07 pkt1=3.62433600999092e-13
+  kt2=-0.019032
+  at=18000.0
+  ute=-0.787381575639998 lute=-3.24301454293405e-07 wute=-4.33954031160632e-06 pute=2.24363657761343e-12
+  ua1=5.52e-10
+  ub1=-5.0978828e-18 lub1=9.78303574919999e-25
+  uc1=-4.1496e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=1.81e-6
+  sbref=1.81e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.48 pmos
* DC IV MOS Parameters
+  lmin=2.0e-05 lmax=1.0e-04 wmin=1.5e-06 wmax=3.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.05900507992+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} wvth0=6.88884083987926e-8
+  k1=0.608210897813333 wk1=-3.78468616208035e-8
+  k2=0.028732595933776 wk2=-1.59468655163159e-9
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=218485.3576 wvsat=-0.0538126505679296
+  ua=2.7537687604592e-09 wua=-5.72640543089371e-17
+  ub=-7.85358136906667e-19 wub=6.4742232675645e-25
+  uc=-5.53294281333333e-11 wuc=4.47069476092341e-17
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0195546283130667 wu0=2.46196299544888e-10
+  a0=0.851800775034667 wa0=1.72427782071682e-7
+  keta=-0.00633154966613333 wketa=-4.64130687951792e-9
+  a1=0.0
+  a2=0.5
+  ags=0.11055232889056 wags=6.91087527176064e-8
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.0877395348729174+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} wvoff=-1.59094951636619e-8
+  nfactor={1.8568872856+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} wnfactor=-4.35841391241019e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.47036533333333e-05 wcit=-1.36927864040533e-11
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-0.62969404356336 wpclm=2.07626729919112e-6
+  pdiblc1=0.39
+  pdiblc2=0.00449373431354613 wpdiblc2=-4.5207766749077e-9
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=442271342.730453 wpscbe1=-316.024252175572
+  pscbe2=1.501581684088e-08 wpscbe2=-4.32555122504007e-17
+  pvag=0.0
+  delta=0.01
+  alpha0=7.93748430502346e-05 walpha0=-8.35707368750219e-11
+  alpha1=0.0
+  beta0=39.0156126693547 wbeta0=-2.18206053289173e-6
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=1.94551350666667e-08 wagidl=-1.36243224720331e-14
+  bgidl=1759707578.66667 wbgidl=46.5554737737812
+  cgidl=1500.46871466667 wcgidl=-0.00145691247339127
+  egidl=0.50686839579552 wegidl=5.43326533015245e-7
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.557185386666667 wkt1=-5.47711456162136e-8
+  kt2=-0.019032
+  at=549674.549386667 wat=-0.293655497221328
+  ute=-1.51728538666667 wute=-5.47711456162136e-8
+  ua1=2.2096e-11
+  ub1=-3.5771875824e-18 wub1=-2.48934856825689e-25
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.49 pmos
* DC IV MOS Parameters
+  lmin=8e-06 lmax=2.0e-05 wmin=1.5e-06 wmax=3.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.05900507992+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} wvth0=6.8888408398793e-8
+  k1=0.608210897813334 wk1=-3.78468616208035e-8
+  k2=0.028732595933776 wk2=-1.59468655163156e-9
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=218485.3576 wvsat=-0.0538126505679296
+  ua=2.7537687604592e-09 wua=-5.72640543089355e-17
+  ub=-7.85358136906667e-19 wub=6.4742232675645e-25
+  uc=-5.53294281333333e-11 wuc=4.47069476092341e-17
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0195546283130667 wu0=2.46196299544888e-10
+  a0=0.851800775034667 wa0=1.72427782071682e-7
+  keta=-0.00633154966613333 wketa=-4.64130687951792e-9
+  a1=0.0
+  a2=0.5
+  ags=0.11055232889056 wags=6.91087527176063e-8
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.0877395348729174+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} wvoff=-1.59094951636618e-8
+  nfactor={1.8568872856+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} wnfactor=-4.35841391241019e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.47036533333333e-05 wcit=-1.36927864040533e-11
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-0.62969404356336 wpclm=2.07626729919112e-6
+  pdiblc1=0.39
+  pdiblc2=0.00449373431354613 wpdiblc2=-4.5207766749077e-9
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=442271342.730453 wpscbe1=-316.024252175572
+  pscbe2=1.501581684088e-08 wpscbe2=-4.3255512250407e-17
+  pvag=0.0
+  delta=0.01
+  alpha0=7.93748430502347e-05 walpha0=-8.35707368750219e-11
+  alpha1=0.0
+  beta0=39.0156126693547 wbeta0=-2.1820605328917e-6
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=1.94551350666667e-08 wagidl=-1.36243224720331e-14
+  bgidl=1759707578.66667 wbgidl=46.5554737737812
+  cgidl=1500.46871466667 wcgidl=-0.00145691247339127
+  egidl=0.50686839579552 wegidl=5.43326533015245e-7
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.557185386666667 wkt1=-5.47711456162132e-8
+  kt2=-0.019032
+  at=549674.549386667 wat=-0.293655497221328
+  ute=-1.51728538666667 wute=-5.47711456162136e-8
+  ua1=2.2096e-11
+  ub1=-3.5771875824e-18 wub1=-2.48934856825688e-25
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.50 pmos
* DC IV MOS Parameters
+  lmin=4e-06 lmax=8e-06 wmin=1.5e-06 wmax=3.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.06995036809706+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=8.69482747497584e-08 wvth0=8.43332607642915e-08 pvth0=-1.22692362706286e-13
+  k1=0.625719531872793 lk1=-1.39086838104944e-07 wk1=-6.25532251075712e-08 pk1=1.96264880902534e-13
+  k2=0.0266112766202987 lk2=1.68515484943324e-08 wk2=1.39869864633901e-09 pk2=-2.37791526741585e-14
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=362170.967602716 lvsat=-1.14142411730058 wvsat=-0.256566840100322 pvsat=1.61065900622637e-6
+  ua=2.29870481856325e-09 lua=3.61498244802724e-15 wua=5.84874853844675e-16 pua=-5.10108727248145e-21
+  ub=-2.45652100133914e-19 lub=-4.28737078551907e-24 wub=-1.14154702909435e-25 pub=6.04989176596282e-30
+  uc=-7.80485551484119e-11 luc=1.80478473095082e-16 wuc=7.67658168637034e-17 puc=-2.54672451470578e-22
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0181348024691192 lu0=1.12789545217343e-08 wu0=2.24970686863577e-09 pu0=-1.59156876098011e-14
+  a0=0.890673769670506 la0=-3.08803182087643e-07 wa0=1.17574254833028e-07 pa0=4.35750935031148e-13
+  keta=-0.000518109104816901 lketa=-4.61813904750416e-08 wketa=-1.28446296018293e-08 pketa=6.51663753737694e-14
+  a1=0.0
+  a2=0.5
+  ags=0.0815000514769466 lags=2.30788386546004e-07 wags=1.10104305166847e-07 pags=-3.2566456910152e-13
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.0908170552274715+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=2.44475139445423e-08 wvoff=-1.1566818501432e-08 pvoff=-3.4497789137088e-14
+  nfactor={1.89027806858771+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-2.65253040976097e-07 wnfactor=-4.82958991551849e-07 pnfactor=3.74297505109207e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.47036533333333e-05 wcit=-1.36927864040533e-11
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-2.0626079646051 lpclm=1.13829248973635e-05 wpclm=4.09824640151743e-06 ppclm=-1.606239979097e-11
+  pdiblc1=0.39
+  pdiblc2=0.00765253625334478 lpdiblc2=-2.50932067295665e-08 wpdiblc2=-8.97814945694981e-09 ppdiblc2=3.54089236432644e-14
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=889483628.574255 lpscbe1=-3552.60967751458 wpscbe1=-947.083719880616 ppscbe1=0.00501307330550211
+  pscbe2=-4.4345459901337e-08 lpscbe2=4.71560046312498e-13 wpscbe2=8.3721204653585e-14 ppscbe2=-6.6541649511138e-19
+  pvag=0.0
+  delta=0.01
+  alpha0=0.000133190643613257 lalpha0=-4.27507338092597e-10 walpha0=-1.59509997786301e-10 palpha0=6.03253894753111e-16
+  alpha1=0.0
+  beta0=40.7273198809008 lbeta0=-1.35976309178014e-05 wbeta0=-4.59744373227562e-06 pbeta0=1.91875625975859e-11
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=2.974026163165e-08 lagidl=-8.17040169195711e-14 wagidl=-2.81376234273748e-14 pagidl=1.15292211459139e-19
+  bgidl=1594954202.43503 lbgidl=1308.78434544653 wbgidl=279.038303960742 pbgidl=-0.00184682035472221
+  cgidl=2151.06276714933 lcgidl=-0.00516825409351705 wcgidl=-0.00237496313847336 pcgidl=7.29290267834554e-9
+  egidl=1.51679065254119 legidl=-8.02272141536191e-06 wegidl=-8.81770723789539e-07 pegidl=1.13208300983315e-11
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.557185386666667 wkt1=-5.47711456162136e-8
+  kt2=-0.019032
+  at=969001.551330936 lat=-3.33109177074508 wat=-0.885366152356878 pat=4.7004902733313e-6
+  ute=-1.47901514828533 lute=-3.04014946677474e-07 wute=-1.0877412591516e-07 pute=4.28994275196799e-13
+  ua1=2.2096e-11
+  ub1=-3.40324934895684e-18 lub1=-1.38174793264912e-24 wub1=-4.94378402284398e-25 pub1=1.94977898076945e-30
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.51 pmos
* DC IV MOS Parameters
+  lmin=2e-06 lmax=4e-06 wmin=1.5e-06 wmax=3.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.02164710222827+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-1.03554975510157e-07 wvth0=2.37078175859632e-08 pvth0=1.16408322644723e-13
+  k1=0.623123809943136 lk1=-1.28849570386569e-07 wk1=-5.88904122755194e-08 pk1=1.81819113374206e-13
+  k2=0.0276705238596586 lk2=1.26739833070207e-08 wk2=2.83739486656649e-09 pk2=-2.94532266971136e-14
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=51440.7790024267 lvsat=0.0840646735201055 wvsat=0.181903286112792 pvsat=-1.18623324545527e-7
+  ua=3.82520147749203e-09 lua=-2.40536772512197e-15 wua=-1.59487437728059e-15 pua=3.49562572015347e-21
+  ub=-3.40986723168707e-18 lub=8.1919772718134e-24 wub=4.24907650223288e-24 pub=-1.11582557839979e-29
+  uc=-9.71143706464489e-11 luc=2.5567214283779e-16 wuc=1.21405941689832e-16 puc=-4.30728639772346e-22
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0191467344513647 lu0=7.28799597695614e-09 wu0=5.91414077597709e-10 pu0=-9.37554667122616e-15
+  a0=0.598732626936566 la0=8.42583490740742e-07 wa0=6.56953183612743e-07 pa0=-1.69150562218317e-12
+  keta=-0.000615662740984527 lketa=-4.57966486893601e-08 wketa=-1.27069720560477e-08 pketa=6.46234677789613e-14
+  a1=0.0
+  a2=0.5
+  ags=0.0621270100284493 lags=3.07193724714732e-07 wags=1.10397395013693e-07 pags=-3.26820486148496e-13
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.0302611298456251+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=-2.14379000168922e-07 wvoff=-9.7017042584054e-08 pvoff=3.02509349622365e-13
+  nfactor={2.75211978453893+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-3.66427058451609e-06 wnfactor=-1.60196971445884e-06 pnfactor=4.78756389518208e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.47036533333333e-05 wcit=-1.36927864040533e-11
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=-0.0403455043395735 leta0=4.74630634564843e-07 weta0=1.69819059791555e-07 peta0=-6.69749389911913e-13
+  etab=-0.173542404768148 letab=4.083608901651e-07 wetab=1.46108273198715e-07 petab=-5.76236418668412e-13
+  dsub=1.06335733280588 ldsub=-1.98519098485311e-06 wdsub=-7.10285518893047e-07 pdsub=2.80129505796229e-12
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=1.25118931397354 lpclm=-1.68636018962285e-06 wpclm=-5.77839683095772e-07 ppclm=2.37961611813604e-12
+  pdiblc1=0.76851754635597 lpdiblc1=-1.49283535107331e-06 wpdiblc1=-5.34124595592725e-07 ppdiblc1=2.10653399255815e-12
+  pdiblc2=-0.00349840803197694 lpdiblc2=1.88850024373138e-08 wpdiblc2=6.75690342029053e-09 ppdiblc2=-2.66485513992838e-14
+  pdiblcb=0.352258634293334 lpdiblcb=-1.48787032778948e-06 wpdiblcb=-5.32348149816786e-07 ppdiblcb=2.09952786806242e-12
+  drout=-0.269968995445334 ldrout=3.27331472113685e-06 wdrout=1.17116592959693e-06 pdrout=-4.61896130973733e-12
+  pscbe1=-517482635.084434 lpscbe1=1996.32456972893 wpscbe1=1038.2807469031 ppscbe1=-0.00281700561504621
+  pscbe2=1.34601939861023e-07 lpscbe2=-2.34190603610273e-13 wpscbe2=-1.68790755361482e-13 ppscbe2=3.30465423992042e-19
+  pvag=0.0
+  delta=0.01
+  alpha0=6.73162259229829e-05 lalpha0=-1.67705222163923e-10 walpha0=-6.65548704812254e-11 palpha0=2.36648168174623e-16
+  alpha1=-1.88629317146667e-10 lalpha1=7.43935163894739e-16 walpha1=2.66174074908393e-16 palpha1=-1.04976393403121e-21
+  beta0=102.114300000692 lbeta0=-0.000255701741812245 wbeta0=-9.12203658313922e-05 pbeta0=3.60819705064292e-10
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=1.85120406657223e-08 lagidl=-3.74210362520489e-14 wagidl=-2.62829762586781e-14 pagidl=1.07977668490516e-19
+  bgidl=2961776362.59237 lbgidl=-4081.82557199804 wbgidl=-1386.48529704197 pbgidl=0.00472183817527238
+  cgidl=1871.05031719089 lcgidl=-0.00406391299212597 wcgidl=-0.0029837874926572 pcgidl=9.69404504881122e-9
+  egidl=-3.97740258429835 legidl=1.36458272914096e-05 wegidl=6.87106337594179e-06 pegidl=-1.92555723075989e-11
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.553585620809333 lkt1=-1.41971165647363e-08 wkt1=-6.80798493616326e-08 pkt1=5.24881967015608e-14
+  kt2=-0.019032
+  at=187874.631921061 lat=-0.250405313284477 wat=0.285550663007722 pat=8.25114452148533e-8
+  ute=-1.62284455814133 lute=2.63233862853605e-07 wute=-1.06469629963358e-07 pute=4.19905573612487e-13
+  ua1=-4.933329728e-10 lua1=2.03280032582592e-15 wua1=-4.93038065763132e-32 pua1=1.88079096131566e-37
+  ub1=-3.51559839977928e-18 lub1=-9.38654511110496e-25 wub1=3.48954212204904e-25 pub1=-1.37624051751492e-30
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.52 pmos
* DC IV MOS Parameters
+  lmin=1e-06 lmax=2e-06 wmin=1.5e-06 wmax=3.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.13464341970687+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=1.16098566036488e-07 wvth0=1.60296763665322e-07 pvth0=-1.49106929638943e-13
+  k1=0.537330494114427 lk1=3.79240562528594e-08 wk1=6.21721925171089e-08 pk1=-5.35144840821846e-14
+  k2=0.0266938129427 lk2=1.45726116584966e-08 wk2=-4.19711208151758e-09 pk2=-1.5778848640733e-14
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=229838.803268882 lvsat=-0.262723245851456 wvsat=-0.0298754469055057 pvsat=2.93053354568742e-7
+  ua=4.32711975260349e-09 lua=-3.38104666011113e-15 wua=-2.24693685250683e-15 pua=4.76316996574575e-21
+  ub=5.53382798107872e-19 lub=4.8781553889502e-25 wub=-1.2346894988055e-24 pub=-4.98363054579445e-31
+  uc=6.66647392168721e-11 luc=-6.26980688255193e-17 wuc=-1.92458738338939e-16 puc=1.79392911735581e-22
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0301286736083654 lu0=-1.40597955503375e-08 wu0=-1.41662077927238e-08 pu0=1.93117944824919e-14
+  a0=1.17972406597633 la0=-2.86805767608665e-07 wa0=-4.00659880472434e-07 pa0=3.64388413092003e-13
+  keta=0.0995706931546326 lketa=-2.4054890591485e-07 wketa=-1.54079538114929e-07 pketa=3.39437598940821e-13
+  a1=0.0
+  a2=0.5
+  ags=-0.657189342525319 lags=1.705472782444e-06 wags=1.14694694249662e-06 pags=-2.34176915150055e-12
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.218686371038114+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=1.51900826185158e-07 wvoff=1.68869061561702e-07 pvoff=-2.14346648226571e-13
+  nfactor={0.00767275952989177+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.67065998739898e-06 wnfactor=2.24233339051717e-06 pnfactor=-2.68537691058078e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=2.38629317146667e-05 lcit=-1.78047212454739e-11 wcit=-2.66174074908393e-11 pcit=2.51241709306032e-17
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.451165112406808 leta0=-4.80816853328447e-07 weta0=-5.23749605456797e-07 peta0=6.78478738464358e-13
+  etab=0.00885491219762986 letab=5.37987457153239e-08 wetab=-1.11271851182427e-07 petab=-7.59151948839106e-14
+  dsub=0.0314189003784409 ldsub=2.07941339425889e-08 wdsub=7.45878675351584e-07 pdsub=-2.93425192298516e-14
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-0.710718331345165 lpclm=2.12739208211219e-06 wpclm=2.19060333111395e-06 ppclm=-3.00196025718623e-12
+  pdiblc1=-0.384486082626327 lpdiblc1=7.48488403305377e-07 wpdiblc1=1.09287421324968e-06 ppdiblc1=-1.0561889919506e-12
+  pdiblc2=0.0104707968941369 lpdiblc2=-8.26973501855878e-09 wpdiblc2=-1.2954985774129e-08 ppdiblc2=1.16693900057482e-14
+  pdiblcb=-0.779517268586667 lpdiblcb=7.12188849818955e-07 wpdiblcb=1.06469629963357e-06 ppdiblcb=-1.00496683722413e-12
+  drout=2.49345344270889 ldrout=-2.09850215639115e-06 wdrout=-2.72828841919275e-06 pdrout=2.96118799887492e-12
+  pscbe1=635639209.37849 lpscbe1=-245.228983722551 wpscbe1=-588.884875331149 ppscbe1=0.000346041638014956
+  pscbe2=1.41063979929357e-08 lpscbe2=4.068022710166e-17 wpscbe2=1.24002178640846e-15 ppscbe2=-5.74037057422394e-23
+  pvag=0.0
+  delta=0.01
+  alpha0=-0.000143180071080662 lalpha0=2.41478529581463e-10 walpha0=2.3047561223543e-10 palpha0=-3.40749387178284e-16
+  alpha1=3.77258634293333e-10 lalpha1=-3.56094424909477e-16 walpha1=-5.32348149816786e-16 palpha1=5.02483418612064e-22
+  beta0=-115.803637608749 lbeta0=0.000167908937106747 wbeta0=0.000216282764257539 pbeta0=-2.36935629515583e-10
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-1.61993393083622e-09 lagidl=1.71350916620121e-15 wagidl=4.08968837023873e-14 pagidl=-2.26132612877987e-20
+  bgidl=216638223.797227 lbgidl=1254.44845600585 wbgidl=1976.76036895751 pbgidl=-0.001815975074864
+  cgidl=-1600.62303317432 lcgidl=0.00268467283364897 wcgidl=0.00478307447260575 pcgidl=-5.40395792546344e-9
+  egidl=5.27915095736141 legidl=-4.34798713822287e-06 wegidl=-6.19082230048014e-06 pegidl=6.13542725879774e-12
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.469016534568 lkt1=-1.78590963309265e-07 wkt1=-1.57399948993234e-07 pkt1=2.26117538375429e-13
+  kt2=-0.019032
+  at=68728.0701815413 lat=-0.0187963119190234 wat=0.689291863382708 pat=-7.02321074194082e-7
+  ute=-1.45040765637867 lute=-7.19662304828435e-08 wute=3.19945647117119e-08 pute=1.50745025583618e-13
+  ua1=5.524e-10
+  ub1=-4.38317573044144e-18 lub1=7.47829061963677e-25 wub1=-6.97908424409807e-25 pub1=6.58755761800416e-31
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=2.81e-6
+  sbref=2.81e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.53 pmos
* DC IV MOS Parameters
+  lmin=8.0e-07 lmax=1e-06 wmin=1.5e-06 wmax=3.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.895522607182498+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-1.09607568905269e-07 wvth0=-2.16142922821868e-07 pvth0=2.06214490436316e-13
+  k1=0.584096513297573 lk1=-6.218389254113e-09 wk1=1.94320219758067e-08 pk1=-1.31720371082504e-14
+  k2=0.0294022146857447 lk2=1.20161512532367e-08 wk2=-2.36968216732599e-08 pk2=2.6269272429126e-15
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=-443869.467793432 lvsat=0.373189991204261 wvsat=1.31380138339977 pvsat=-9.75243205556412e-7
+  ua=-8.76687454415665e-09 lua=8.97837455660077e-15 wua=2.29329648124585e-14 pua=-1.9004139215815e-20
+  ub=1.02639083957859e-17 lub=-8.6779495727533e-24 wub=-2.06378560688182e-23 pub=1.78162858708556e-29
+  uc=1.23205222394029e-11 luc=-1.14025624204861e-17 wuc=-1.72105672585023e-17 puc=1.39761630527572e-23
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=-0.00820370044372129 lu0=2.21221323174272e-08 wu0=5.56790732590781e-08 pu0=-4.6615166302304e-14
+  a0=0.83003867988532 la0=4.32622683226459e-08 wa0=4.14865790354194e-07 pa0=-4.05386267601247e-13
+  keta=-0.488341483890459 lketa=3.14381397998011e-07 wketa=9.64173000009874e-07 pketa=-7.16080971795181e-13
+  a1=0.0
+  a2=0.5
+  ags=2.79469540147411 lags=-1.55276122741706e-06 wags=-6.4447101895845e-06 pags=4.82399601547081e-12
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.0394951063033218+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=-1.72378085980128e-08 wvoff=-1.64809868700592e-07 pvoff=1.00612894048008e-13
+  nfactor={1.68848013126916+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=8.41459092142792e-08 wnfactor=-4.8603685676439e-07 pnfactor=-1.10068234171711e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-1.35975e-05 lcit=1.755418025e-11
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=-0.256068819221202 leta0=1.86741254735232e-07 weta0=8.58293790166119e-07 peta0=-6.26032022664112e-13
+  etab=0.300297325726016 letab=-2.2129374841412e-07 wetab=-8.68434808881125e-07 petab=6.38770920887891e-13
+  dsub=-0.803606631610877 ldsub=8.08974733587306e-07 wdsub=3.47142821617863e-06 pdsub=-2.6019887308165e-12
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=4.29808375447819 lpclm=-2.60041620669647e-06 wpclm=-6.50956192311701e-06 ppclm=5.21012572628236e-12
+  pdiblc1=0.21832819866173 lpdiblc1=1.7949200319758e-07 wpdiblc1=-9.43662870745572e-08 ppdiblc1=6.44473163054426e-14
+  pdiblc2=-0.0511958210929221 lpdiblc2=4.99373856994262e-08 wpdiblc2=4.61738267425332e-08 ppdiblc2=-4.41422961287291e-14
+  pdiblcb=-0.025
+  drout=0.0692316924848506 ldrout=1.89720753645325e-07 wdrout=7.65484843198145e-07 pdrout=-3.3658458349584e-13
+  pscbe1=177203717.134327 lpscbe1=187.488277406715 wpscbe1=-732.450504797039 ppscbe1=0.000481553235667809
+  pscbe2=1.64844728078746e-08 lpscbe2=-2.20398459071914e-15 wpscbe2=5.76140713689137e-15 ppscbe2=-4.32513933806306e-21
+  pvag=0.0
+  delta=0.01
+  alpha0=0.000520769267904426 lalpha0=-3.85223251486562e-10 walpha0=-7.71003398902507e-10 palpha0=6.04546651434815e-16
+  alpha1=0.0
+  beta0=131.693313972747 lbeta0=-6.57034354910272e-05 wbeta0=-0.00018533127827677 pbeta0=1.42147865232552e-10
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-9.25349756400139e-08 lagidl=8.7528217035494e-14 wagidl=1.71119956108947e-13 pagidl=-1.4553081933235e-19
+  bgidl=506981834.976002 lbgidl=980.393121414207 wbgidl=439.924580146711 pbgidl=-0.000365355773805481
+  cgidl=3900.093286032 lcgidl=-0.00250745330004987 wcgidl=-0.00434420901579461 pcgidl=3.21128495923766e-9
+  egidl=0.269883035323943 legidl=3.80260853388298e-07 wegidl=4.70809256425089e-06 pegidl=-4.15205848202188e-12
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.724138601440001 lkt1=6.22187556112168e-08 wkt1=3.87738632603579e-07 pkt1=-2.88438768793802e-13
+  kt2=-0.019032
+  at=119897.829053333 lat=-0.067095447318108 wat=-0.207562102705843 pat=1.44219384396901e-7
+  ute=-1.70091398669333 lute=1.64486694701171e-07 wute=9.04723476075018e-07 pute=-6.73023793852205e-13
+  ua1=5.524e-10
+  ub1=-3.5909e-18
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=2.41e-6
+  sbref=2.41e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.54 pmos
* DC IV MOS Parameters
+  lmin=6e-07 lmax=8.0e-07 wmin=1.5e-06 wmax=3.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.02862658583924+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-1.05915191825193e-08 wvth0=-5.97810349201635e-09 pvth0=4.98728813368385e-14
+  k1=0.70465093572872 lk1=-9.58988241006425e-08 wk1=-3.73554562716134e-07 pk1=2.79170683244085e-13
+  k2=0.0110325251852878 lk2=2.56813632726266e-08 wk2=7.26855194486576e-08 pk2=-6.90718963176819e-14
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=16975.2351048947 lvsat=0.0303676167181963 wvsat=-0.0144898660937309 pvsat=1.28726549418066e-8
+  ua=3.96786712628672e-09 lua=-4.94999772042065e-16 wua=-4.52006680484848e-15 pua=1.41817100429965e-21
+  ub=-1.4504259530004e-18 lub=3.63437493088538e-26 wub=5.12582400404346e-24 pub=-1.34931573534624e-30
+  uc=-5.21806584618427e-12 luc=1.6443932563822e-18 wuc=8.01211009576364e-18 puc=-4.78698663108121e-24
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0265851294483591 lu0=-3.75727823929148e-09 wu0=-1.38000261300169e-08 pu0=5.07033573324381e-15
+  a0=1.00587729087467 la0=-8.75440743923313e-08 wa0=-4.72666770996079e-07 pa0=2.54849204787218e-13
+  keta=-0.149113475749536 lketa=6.20296827419791e-08 wketa=6.88350722571913e-08 pketa=-5.00390873399598e-14
+  a1=0.0
+  a2=0.5
+  ags=0.672743314091913 lags=2.57589303865584e-08 wags=1.4082917684029e-07 pags=-7.4986719212588e-14
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.0533360795669392+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=-6.94150858720771e-09 wvoff=-5.67234375057776e-08 pvoff=2.0207397882186e-14
+  nfactor={2.47485455920586+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-5.00838027727829e-07 wnfactor=-2.2063825241174e-06 pnfactor=1.16969690777219e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.0257190304886185 leta0=-2.28807266639039e-08 weta0=-6.90811072009412e-08 peta0=6.38421634872439e-14
+  etab=0.0104871609673172 letab=-5.70396685012381e-09 wetab=-3.62886671938914e-08 petab=1.97374060867575e-14
+  dsub=0.300809479024667 ldsub=-1.2600411114475e-08 wdsub=-7.56198627770735e-08 pdsub=3.66603351186467e-14
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.667317290607857 lpclm=1.00510965776667e-07 wpclm=8.87546501359935e-07 ppclm=-2.92583230686034e-13
+  pdiblc1=0.317425897875466 lpdiblc1=1.05773224752482e-07 wpdiblc1=4.06189335710084e-07 ppdiblc1=-3.07916011484052e-13
+  pdiblc2=0.0191169730567227 lpdiblc2=-2.36830186849457e-09 wpdiblc2=-2.24330427626372e-08 ppdiblc2=6.89435409616708e-15
+  pdiblcb=-0.025
+  drout=0.570347228843731 ldrout=-1.83059093852046e-07 wdrout=-4.03337820294467e-07 pdrout=5.32902595876315e-13
+  pscbe1=351466585.545357 lpscbe1=57.8541295957491 wpscbe1=141.285428685253 ppscbe1=-0.000168418925249667
+  pscbe2=1.64149662757392e-08 lpscbe2=-2.15227868146367e-15 wpscbe2=-8.47522305339931e-15 ppscbe2=6.26548986049417e-21
+  pvag=0.0
+  delta=0.01
+  alpha0=-4.23801992141437e-06 lalpha0=5.32966992708075e-12 walpha0=6.25250756785657e-11 palpha0=-1.55151808060451e-17
+  alpha1=0.0
+  beta0=45.23147742094 lbeta0=-1.38447528013778e-06 wbeta0=3.35511321891257e-07 pbeta0=4.03034045010795e-12
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=1.51979351981126e-07 lagidl=-9.43659912818723e-14 wagidl=-3.54115085291985e-13 pagidl=2.45191527965803e-19
+  bgidl=1211407235.35627 lbgidl=456.371066071327 wbgidl=1734.70104358331 pbgidl=-0.00132853998495598
+  cgidl=1695.99988055467 lcgidl=-0.000867828215715283 wcgidl=-0.00342344854828317 pcgidl=2.5263312474559e-9
+  egidl=3.47005626849778 legidl=-2.00034801476972e-06 wegidl=-8.70132212377969e-06 pegidl=5.82320510440407e-12
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.647423426384 lkt1=5.15033688705675e-09 wkt1=5.95800522013155e-08 pkt1=-4.4321600832559e-14
+  kt2=-0.019032
+  at=41065.2021893333 lat=-0.00845185619397841 wat=0.00864973317144052 pat=-1.66206003122099e-8
+  ute=-1.2439681407272 lute=-1.75435320113037e-07 wute=-8.64655507571611e-07 pute=6.43217232082523e-13
+  ua1=5.534878e-10 lua1=-8.09214420000522e-19
+  ub1=-7.26808098179201e-19 lub1=-2.1305979657645e-24 wub1=-1.06469553283753e-23 pub1=7.92027006877841e-30
+  uc1=-4.66529325417792e-10 luc1=2.65817285178296e-16 wuc1=5.04225981779745e-16 puc1=-3.75093707845952e-22
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=2.02e-6
+  sbref=2.01e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.55 pmos
* DC IV MOS Parameters
+  lmin=5e-07 lmax=6e-07 wmin=1.5e-06 wmax=3.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.778216308142747+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-1.4678966922164e-07 wvth0=-1.13588249451883e-07 pvth0=1.08402039724409e-13
+  k1=0.440256587387308 lk1=4.79052619622514e-08 wk1=4.9420344270612e-07 pk1=-1.92802895905079e-13
+  k2=0.128555937615153 lk2=-3.8239620747977e-08 wk2=-2.56056288481177e-07 pk2=1.09730773015355e-13
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=-510216.811962977 lvsat=0.317107371118412 wvsat=0.796710342921749 pvsat=-4.28339138741713e-7
+  ua=1.25191715270904e-09 lua=9.82205418586836e-16 wua=-2.04577436485465e-16 pua=-9.29023663152995e-22
+  ub=-8.34325113504028e-18 lub=3.78535136582034e-24 wub=1.27302591560619e-23 pub=-5.48536801452908e-30
+  uc=2.82874665477458e-10 luc=-1.55049243310547e-16 wuc=-3.97312645819642e-16 puc=2.15669148111308e-22
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=-0.000736936539163291 lu0=1.1103193451322e-08 wu0=1.96750901856838e-08 pu0=-1.31367800308658e-14
+  a0=0.0254332938542401 la0=4.45719415587079e-07 wa0=1.3186361163601e-06 pa0=-7.19440435645807e-13
+  keta=-0.383888412194913 lketa=1.8972377067462e-07 wketa=4.47945344595313e-07 pketa=-2.56237164464664e-13
+  a1=0.0
+  a2=0.5
+  ags=5.81395912795155 lags=-2.7705483507717e-06 wags=-7.96242234994195e-06 pags=4.33237178620427e-12
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={0.295043641987348+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=-1.96425239140585e-07 wvoff=-4.55890701324647e-07 pvoff=2.37314472673269e-13
+  nfactor={5.47478504231172+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-2.13250021748911e-06 wnfactor=-5.35767705232038e-06 pnfactor=2.88368600166179e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=-1.08015108272097 leta0=5.78602027910793e-07 weta0=1.29001941343276e-06 peta0=-6.75372609685427e-13
+  etab=0.071837469619728 letab=-3.90723997261701e-08 wetab=-1.38948289445597e-08 petab=7.55739746294602e-15
+  dsub=0.127292160329826 ldsub=8.17756585236495e-08 wdsub=1.92600934162968e-07 pdsub=-1.09224956337041e-13
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=3.7387475926299 lpclm=-1.57003997549312e-06 wpclm=-3.31735491237565e-06 ppclm=1.99446264824475e-12
+  pdiblc1=1.93398804539203 lpdiblc1=-7.73474927281778e-07 wpdiblc1=-8.41436717746791e-07 ppdiblc1=3.70667798991143e-13
+  pdiblc2=0.0635275279132733 lpdiblc2=-2.65232026549724e-08 wpdiblc2=-5.37339915641669e-08 ppdiblc2=2.39189401493191e-14
+  pdiblcb=1.69798068586667 lpdiblcb=-9.37129195042879e-07 wpdiblcb=-2.43129115390371e-06 ppdiblcb=1.32237925860823e-12
+  drout=-3.16747236083941 ldrout=1.84994098097661e-06 wdrout=3.13527155418154e-06 pdrout=-1.39174704290119e-12
+  pscbe1=741229513.334433 lpscbe1=-154.137926828729 wpscbe1=-584.315136587622 ppscbe1=0.00022623522220225
+  pscbe2=4.06725141993201e-09 lpscbe2=4.56364342860987e-15 wpscbe2=1.40369844296393e-14 ppscbe2=-5.97889978953056e-21
+  pvag=0.0
+  delta=0.01
+  alpha0=0.000106203181103928 lalpha0=-5.47392993106031e-11 walpha0=-3.61975426917301e-11 palpha0=3.81800513255588e-17
+  alpha1=-8.61490342933333e-10 lalpha1=4.6856459752144e-16 walpha1=1.21564557695185e-15 palpha1=-6.61189629304113e-22
+  beta0=398.26396383871 lbeta0=-0.000193398844642763 wbeta0=-0.000480156463511855 pbeta0=2.65369925562183e-10
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-2.22087636667168e-07 lagidl=1.09089043843935e-13 wagidl=6.21040419581983e-13 pagidl=-2.85195551135148e-19
+  bgidl=7686677615.31466 lbgidl=-3065.52849358805 wbgidl=-9527.42571787525 pbgidl=0.00479693076060134
+  cgidl=-3985.65118531765 lcgidl=0.00222242179901267 wcgidl=0.00990621167810099 pcgidl=-4.72367094967445e-9
+  egidl=-15.6780969133639 legidl=8.41433250084487e-06 wegidl=2.74122102870589e-05 pegidl=-1.3818945173851e-11
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-1.03687067812267 lkt1=2.16970697107719e-07 wkt1=4.15723949456183e-07 pkt1=-2.38028266549482e-13
+  kt2=-0.019032
+  at=4646.32818666671 lat=0.011356369376072 wat=0.0388738206011073 pat=-3.30594814652057e-8
+  ute=-2.98569689182347 lute=7.71890947608224e-07 wute=2.05996661207413e-06 pute=-9.47484738792796e-13
+  ua1=5.52e-10
+  ub1=-9.34750978651093e-18 lub1=2.55820168251914e-24 wub1=1.2371072121924e-23 pub1=-4.59923506143941e-30
+  uc1=2.21952290559999e-11 wuc1=-1.85411282140005e-16
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=1.81e-6
+  sbref=1.81e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.56 pmos
* DC IV MOS Parameters
+  lmin=2.0e-05 lmax=1.0e-04 wmin=1e-06 wmax=1.5e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.012257832304+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} wvth0=2.92355427684563e-9
+  k1=0.57508521568 wk1=8.89665593481486e-9
+  k2=0.02920354177888 wk2=-2.25923634987447e-9
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=362922.705248 wvsat=-0.257627614084632
+  ua=3.5189278207248e-09 wua=-1.13697694361348e-15
+  ub=-1.43755868432e-18 wub=1.56773991040922e-24
+  uc=1.5460123027744e-11 wuc=-5.51839048759574e-17
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0213840147744 wu0=-2.33524361849673e-9
+  a0=1.075963042128 wa0=-1.43886696374653e-7
+  keta=-0.0122424698496 wketa=3.69956894769116e-9
+  a1=0.0
+  a2=0.5
+  ags=0.16570511887456 wags=-8.71712861765621e-9
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.083222932284432+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} wvoff=-2.22828550098632e-8
+  nfactor={1.60190221744+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} wnfactor=-7.60329815007141e-8
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=5.0e-6
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=2.22320713069008 wpclm=-1.94945013619321e-6
+  pdiblc1=0.39
+  pdiblc2=-0.0026241897739872 wpdiblc2=5.52329753331424e-9
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=206647509.73088 wpscbe1=16.4635960747942
+  pscbe2=1.496045407648e-08 wpscbe2=3.48666631433759e-17
+  pvag=0.0
+  delta=0.01
+  alpha0=-6.0192853181488e-05 walpha0=1.13372681006777e-10
+  alpha1=0.0
+  beta0=34.608004388992 wbeta0=4.03749788109497e-6
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-8.7863584e-09 wagidl=2.62271359928064e-14
+  bgidl=2288882881.6 wbgidl=-700.161679494234
+  cgidl=-1230.282944 wcgidl=0.00239644026914662
+  egidl=-0.25248076426096 wegidl=1.6148410953743e-6
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.66888768 wkt1=1.0285151369728e-7
+  kt2=-0.019032
+  at=688661.13216 wat=-0.489778908226447
+  ute=-1.5561
+  ua1=2.2096e-11
+  ub1=-4.9870417648e-18 wub1=1.74050474054222e-24
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.57 pmos
* DC IV MOS Parameters
+  lmin=8e-06 lmax=2.0e-05 wmin=1e-06 wmax=1.5e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.012257832304+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} wvth0=2.92355427684521e-9
+  k1=0.57508521568 wk1=8.89665593481465e-9
+  k2=0.02920354177888 wk2=-2.25923634987447e-9
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=362922.705248 wvsat=-0.257627614084632
+  ua=3.5189278207248e-09 wua=-1.13697694361348e-15
+  ub=-1.43755868432e-18 wub=1.56773991040921e-24
+  uc=1.5460123027744e-11 wuc=-5.51839048759575e-17
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0213840147744 wu0=-2.33524361849674e-9
+  a0=1.075963042128 wa0=-1.43886696374652e-7
+  keta=-0.0122424698496 wketa=3.69956894769115e-9
+  a1=0.0
+  a2=0.5
+  ags=0.16570511887456 wags=-8.71712861765621e-9
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.0832229322844319+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} wvoff=-2.22828550098631e-8
+  nfactor={1.60190221744+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} wnfactor=-7.60329815007132e-8
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=5.0e-6
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=2.22320713069008 wpclm=-1.94945013619321e-6
+  pdiblc1=0.39
+  pdiblc2=-0.0026241897739872 wpdiblc2=5.52329753331424e-9
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=206647509.73088 wpscbe1=16.4635960747943
+  pscbe2=1.496045407648e-08 wpscbe2=3.48666631433823e-17
+  pvag=0.0
+  delta=0.01
+  alpha0=-6.0192853181488e-05 walpha0=1.13372681006777e-10
+  alpha1=0.0
+  beta0=34.608004388992 wbeta0=4.03749788109497e-6
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-8.78635840000001e-09 wagidl=2.62271359928064e-14
+  bgidl=2288882881.6 wbgidl=-700.161679494234
+  cgidl=-1230.282944 wcgidl=0.00239644026914662
+  egidl=-0.25248076426096 wegidl=1.6148410953743e-6
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.66888768 wkt1=1.0285151369728e-7
+  kt2=-0.019032
+  at=688661.13216 wat=-0.489778908226448
+  ute=-1.5561
+  ua1=2.2096e-11
+  ub1=-4.9870417648e-18 wub1=1.74050474054222e-24
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.58 pmos
* DC IV MOS Parameters
+  lmin=4e-06 lmax=8e-06 wmin=1e-06 wmax=1.5e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.991957644883398+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-1.61262658850528e-07 wvth0=-2.57219589916179e-08 pvth0=2.27557092853341e-13
+  k1=0.6114670897633 lk1=-2.89013969530326e-07 wk1=-4.24416610566331e-08 pk1=4.07826456348366e-13
+  k2=0.0168597845552095 lk2=9.8057573009116e-08 wk2=1.51589900934181e-08 pk2=-1.38368649042872e-13
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=434921.086582033 lvsat=-0.571947941479424 wvsat=-0.35922424199156 pvsat=8.07073452429849e-7
+  ua=3.07621790547527e-09 lua=3.51684329575074e-15 wua=-5.12270753044532e-16 pua=-4.9626035072607e-21
+  ub=-1.3146148994548e-18 lub=-9.76653132590631e-25 wub=1.39425442736108e-24 pub=1.37815132878611e-30
+  uc=4.27807006023209e-11 luc=-2.17031936194682e-16 wuc=-9.37358626091327e-17 puc=3.06252897036571e-22
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0199701881979866 lu0=1.12312969403704e-08 wu0=-3.40198591826108e-10 pu0=-1.58484381873689e-14
+  a0=1.03010391442547 la0=3.64300324556126e-07 wa0=-7.9175064710123e-08 pa0=-5.14062730779852e-13
+  keta=-0.0151984746609212 lketa=2.34822066206542e-08 wketa=7.8707755129272e-09 pketa=-3.31356478335786e-14
+  a1=0.0
+  a2=0.5
+  ags=0.180147034048018 lags=-1.14725129946436e-07 wags=-2.90960573512626e-08 pags=1.61888171966896e-13
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.0641612575196907+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=-1.51424038163628e-07 wvoff=-4.91807080236904e-08 pvoff=2.13673854556543e-13
+  nfactor={1.72299546747528+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-9.61952668955258e-07 wnfactor=-2.46907182252498e-07 pnfactor=1.35740756335209e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.3983178786e-05 lcit=-7.13614739581054e-11 wcit=-1.26761276522095e-11 pcit=1.00697890456387e-16
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=3.71457851861628 lpclm=-1.18473051685469e-05 wpclm=-4.05391833621031e-06 ppclm=1.67176849341159e-11
+  pdiblc1=0.39
+  pdiblc2=-0.00648348303639423 lpdiblc2=3.06578397472352e-08 wpdiblc2=1.09691308187238e-08 ppdiblc2=-4.32611550359646e-14
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=207260270.322231 lpscbe1=-4.86770886163049 wpscbe1=15.5989320553817 ppscbe1=6.86880450381094e-6
+  pscbe2=1.49760237219519e-08 lpscbe2=-1.23683706664227e-16 wpscbe2=1.28963986965499e-17 ppscbe2=1.74529583739067e-22
+  pvag=0.0
+  delta=0.01
+  alpha0=-0.000175613299475475 lalpha0=9.16888483314804e-10 walpha0=2.76242011090437e-10 palpha0=-1.29381767125159e-15
+  alpha1=1.7966357572e-10 lalpha1=-1.42722947916211e-15 walpha1=-2.53522553044189e-16 palpha1=2.01395780912773e-21
+  beta0=-30.1418104566307 lbeta0=0.000514366054152143 wbeta0=9.54057026104938e-05 pbeta0=-7.25819881549872e-10
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=1.564788789792e-08 lagidl=-1.94103209166047e-13 wagidl=-8.25193122120332e-15 pagidl=2.73898262041372e-19
+  bgidl=2202464701.67868 lbgidl=686.497379476976 wbgidl=-578.217331479978 pbgidl=-0.000968713706190442
+  cgidl=-2861.6282115376 lcgidl=0.0129592436707919 wcgidl=0.00469842505078786 pcgidl=-1.82867369068798e-8
+  egidl=0.610020821192107 legidl=-6.85162634468062e-06 wegidl=3.97768558147824e-07 pegidl=9.66830252847344e-12
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.704820395144 lkt1=2.85445895832422e-07 wkt1=1.53556024306118e-07 pkt1=-4.02791561825544e-13
+  kt2=-0.019032
+  at=811838.479673632 lat=-0.978508530913542 wat=-0.663593970593544 pat=1.38076947393797e-6
+  ute=-1.29433017017596 lute=-2.07947335113919e-06 wute=-3.69382359785384e-07 pute=2.9343365278991e-12
+  ua1=2.2096e-11
+  ub1=-3.77089902075132e-18 lub1=-9.66091634444831e-24 wub1=2.4410578986104e-26 pub1=1.36324804099856e-29
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.59 pmos
* DC IV MOS Parameters
+  lmin=2e-06 lmax=4e-06 wmin=1e-06 wmax=1.5e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.00778414493964+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-9.88445252787055e-08 wvth0=4.14585400780561e-09 pvth0=1.09761425164918e-13
+  k1=0.517605883722672 lk1=8.11652409733055e-08 wk1=9.00055113424721e-08 pk1=-1.14531946876467e-13
+  k2=0.0571286306222665 lk2=-6.075872899475e-08 wk2=-3.87308217537224e-08 pk2=7.41673799010658e-14
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=114272.854074038 lvsat=0.692656622708856 wvsat=0.0932411963075406 pvsat=-9.77404989677976e-7
+  ua=3.34839408331171e-09 lua=2.4434076679816e-15 wua=-9.22053370582323e-16 pua=-3.3464618419534e-21
+  ub=-1.39039577847626e-18 lub=-6.77780923817926e-25 wub=1.39940841249292e-24 pub=1.35782452682463e-30
+  uc=5.43673736140794e-11 luc=-2.62728615885756e-16 wuc=-9.23493417092227e-17 puc=3.00784597259416e-22
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0205017262128699 lu0=9.13496416347205e-09 wu0=-1.32060937709519e-09 pu0=-1.19817960913461e-14
+  a0=1.51708171600811 la0=-1.55629142710565e-06 wa0=-6.38925542579758e-07 pa0=1.6935371788902e-12
+  keta=-0.19530127936236 lketa=7.33789658082659e-07 wketa=2.62013122815909e-07 pketa=-1.03544765136181e-12
+  a1=0.0
+  a2=0.5
+  ags=1.02840962834401 lags=-3.46018797559041e-06 wags=-1.25312014256093e-06 pags=4.98931676162529e-12
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.0832282087966044+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=-7.62258890226084e-08 wvoff=-2.22754093446428e-08 pvoff=1.07562047096246e-13
+  nfactor={1.65645172828243+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-6.99510815952587e-07 wnfactor=-5.58769029475216e-08 pnfactor=6.04003244801201e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-9.5198729669997e-06 lcit=2.13322118505501e-11 wcit=2.04889346642414e-11 pcit=-3.01017988134638e-17
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0={-0.0616863611519999+5e-17} leta0=5.58796839747372e-07 weta0=1.99933057476143e-07 peta0=-7.88515985380159e-13
+  etab=0.0528279064826688 letab=-4.84420980376997e-07 wetab=-1.73321967526068e-07 petab=6.8356450772606e-13
+  dsub=0.0286761456800004 ldsub=2.09548814905265e-06 wdsub=7.49748965535534e-07 pdsub=-2.9569349451756e-12
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=2.46383535837796 lpclm=-6.91449921888303e-06 wpclm=-2.28899966577067e-06 ppclm=9.75702218976897e-12
+  pdiblc1=0.391608671522929 lpdiblc1=-6.34443961928124e-09 wpdiblc1=-2.26998995131948e-09 ppdiblc1=8.95261336900995e-15
+  pdiblc2=0.00129
+  pdiblcb=-0.025
+  drout=0.698144503206717 ldrout=-5.44828106196973e-07 wdrout=-1.94935155896986e-07 pdrout=7.68804761342123e-13
+  pscbe1=356291166.742006 lpscbe1=-592.630661251581 wpscbe1=-194.697969758977 ppscbe1=0.000836258755569462
+  pscbe2=1.45205283806585e-08 lpscbe2=1.67274436986279e-15 wpscbe2=6.55644052814284e-16 ppscbe2=-2.36040288933589e-21
+  pvag=0.0
+  delta=0.01
+  alpha0=0.000623202687782588 lalpha0=-2.23356188883227e-09 walpha0=-8.50964033265466e-10 palpha0=3.15177024708366e-15
+  alpha1=-3.5932715144e-10 lalpha1=6.98496049684216e-16 walpha1=5.07045106088378e-16 palpha1=-9.85644981725198e-22
+  beta0=192.983424289945 lbeta0=-0.000365617559164877 wbeta0=-0.00021944542363946 pbeta0=5.15921475267322e-10
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-5.021216175472e-08 lagidl=6.56422406590002e-14 wagidl=7.06934708799984e-14 pagidl=-3.74545093055576e-20
+  bgidl=3139002579.88288 lbgidl=-3007.11435837257 wbgidl=-1636.56850335573 pbgidl=0.00320531748057034
+  cgidl=-967.294541529599 lcgidl=0.00548818110964739 wcgidl=0.00102138958410385 pcgidl=-3.78487672982476e-9
+  egidl=-2.08882249462395 legidl=3.79234180856631e-06 wegidl=4.20609556572259e-06 pegidl=-5.35135835670069e-12
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.717974118148 lkt1=3.37322863987898e-07 wkt1=1.6388810167897e-07 pkt1=-4.43540241776339e-13
+  kt2=-0.019032
+  at=341875.415792487 lat=0.874978796727309 wat=0.0682407728898893 pat=-1.50551357088634e-6
+  ute=-2.21120946756168 lute=1.53660690982035e-06 wute=7.23769740260057e-07 pute=-1.3769460394701e-12
+  ua1=-1.01995243298176e-10 lua1=4.89403454443677e-16 wua1=-5.52215104749105e-16 pua1=2.17788115162e-21
+  ub1=-5.56126888628592e-18 lub1=-2.59987663176641e-24 wub1=3.23559165303247e-24 pub1=9.67903372054147e-31
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.60 pmos
* DC IV MOS Parameters
+  lmin=1e-06 lmax=2e-06 wmin=1e-06 wmax=1.5e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.049606097227+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-1.75468322273063e-08 wvth0=4.03009380632684e-08 pvth0=3.94795572695022e-14
+  k1=0.564158406730352 lk1=-9.32820850132312e-09 wk1=2.43154323364275e-08 pk1=1.31629977033827e-14
+  k2=0.02157975420417 lk2=8.34473187438773e-09 wk2=3.01931574818715e-09 pk2=-6.99071238889613e-15
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=593232.582453334 lvsat=-0.238393193287658 wvsat=-0.54265895513757 pvsat=2.58721314716176e-7
+  ua=3.42728534049076e-09 lua=2.29005095315125e-15 wua=-9.77184112912203e-16 pua=-3.23929319193834e-21
+  ub=-7.64189450626385e-19 lub=-1.89506340452529e-24 wub=6.24531431094415e-25 pub=2.86410789096519e-30
+  uc=-1.56967729137593e-10 luc=1.4808569035322e-16 wuc=1.23108143226174e-16 puc=-1.18043207706502e-22
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.022831869101247 lu0=4.60539940275584e-09 wu0=-3.86971613994708e-09 pu0=-7.02658745503828e-15
+  a0=0.676045898581525 la0=7.85980983898919e-08 wa0=3.10078366825713e-07 pa0=-1.51231520603096e-13
+  keta=0.229388169458045 lketa=-9.17641614793255e-08 wketa=-3.37264459656769e-07 pketa=1.2948804120683e-13
+  a1=0.0
+  a2=0.5
+  ags=-0.777757072085547 lags=5.08194733746114e-08 wags=1.31707958340814e-06 pags=-6.89448568597277e-15
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.111238985682306+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=-2.17757398344939e-08 wvoff=1.72504858756625e-08 pvoff=3.07276593774949e-14
+  nfactor={1.4395046381311+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-2.77787367407421e-07 wnfactor=2.21881153950511e-07 pnfactor=6.40693579971145e-14
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-1.89296921000061e-06 lcit=6.50627363731958e-12 wcit=9.72664128035502e-12 pcit=-9.18097670452711e-18
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.29378629625281 leta0=-1.32206458981837e-07 weta0=-3.01672987497155e-07 peta0=1.86556005443434e-13
+  etab=-0.196610290228699 letab=4.61930210230406e-10 wetab=1.78659274100556e-07 petab=-6.51827871935287e-16
+  dsub=1.18906739503144 ldsub=-1.60196400561619e-07 wdsub=-8.87674484859288e-07 pdsub=2.26052500046898e-13
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-2.18637803083799 lpclm=2.12505058841387e-06 wpclm=4.27290083042948e-06 ppclm=-2.9986561847945e-12
+  pdiblc1=0.275412985873961 lpdiblc1=2.19528353713749e-07 wpdiblc1=1.61693277285197e-07 ppdiblc1=-3.09775581812056e-13
+  pdiblc2=0.0025330225796676 lpdiblc2=-2.41631159261585e-09 wpdiblc2=-1.75402419007863e-09 ppdiblc2=3.40964762309386e-15
+  pdiblcb=-0.025
+  drout=1.04049591866945 ldrout=-1.21032502271497e-06 wdrout=-6.78025868850781e-07 pdrout=1.70788479825301e-12
+  pscbe1=53375503.2923212 lpscbe1=-3.79290307174051 wpscbe1=232.745111272218 ppscbe1=5.35215035292079e-6
+  pscbe2=1.477988530028e-08 lpscbe2=1.16858045381057e-15 wpscbe2=2.89666540964093e-16 ppscbe2=-1.64897920405029e-21
+  pvag=0.0
+  delta=0.01
+  alpha0=-0.00094811931468297 lalpha0=8.20930951760527e-10 walpha0=1.36632215912567e-09 palpha0=-1.15841238230547e-15
+  alpha1=0.0
+  beta0=-4.37485550059802 lbeta0=1.8027200919959e-05 wbeta0=5.90460555398559e-05 pbeta0=-2.54381111093506e-11
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-6.12280683659699e-08 lagidl=8.7056061520609e-14 wagidl=1.25009683771267e-13 pagidl=-1.43039795544894e-19
+  bgidl=1531533988.80688 lbgidl=117.643835820067 wbgidl=121.316214535446 pbgidl=-0.000211834622538318
+  cgidl=2692.96756621238 lcgidl=-0.00162700240159225 wcgidl=-0.00127559404782643 pcgidl=6.80229752284515e-10
+  egidl=-2.47204537237979 legidl=4.5372887606359e-06 wegidl=4.74685983563235e-06 pegidl=-6.40255002097827e-12
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.5573657713744 lkt1=2.51162986946962e-08 wkt1=-3.27306943326695e-08 pkt1=-6.13329642093128e-14
+  kt2=-0.019032
+  at=1564510.75806232 lat=-1.50170204511103 wat=-1.42140110435511 pat=1.39020127429022e-6
+  ute=-1.550465108872 lute=2.5218595096348e-07 wute=1.73185235695244e-07 pute=-3.06664821046564e-13
+  ua1=-2.30275459003648e-10 lua1=7.38767365753544e-16 wua1=1.10443020949821e-15 pua1=-1.04247167474536e-21
+  ub1=-1.00209767098176e-17 lub1=6.06934940639684e-24 wub1=7.25756998638398e-24 pub1=-6.85042031014784e-30
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=2.81e-6
+  sbref=2.81e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.61 pmos
* DC IV MOS Parameters
+  lmin=8.0e-07 lmax=1e-06 wmin=1e-06 wmax=1.5e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.32337513199936+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=2.40863759694323e-07 wvth0=3.87598063537109e-07 pvth0=-2.88334199465255e-13
+  k1=0.469901838057278 lk1=7.96405666691899e-08 wk1=1.80571671428684e-07 pk1=-1.34327266375798e-13
+  k2=0.0272812247585189 lk2=2.96311381813778e-09 wk2=-2.07039012709116e-08 pk2=1.54016321554311e-14
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=1385399.23440022 lvsat=-0.986119296060325 wvsat=-1.26747236519088 pvsat=9.42872692465498e-7
+  ua=2.22311944696024e-08 lua=-1.54589588738172e-14 wua=-2.08082863805808e-14 pua=1.54792842385141e-20
+  ub=-1.65988079698577e-17 lub=1.30512330157771e-23 wub=1.7268015543876e-23 pub=-1.28456767630893e-29
+  uc=6.64875314508049e-12 luc=-6.35190727339537e-18 wuc=-9.20715657658034e-18 puc=6.84920377731812e-24
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0690944676871143 lu0=-3.90618674024444e-08 wu0=-5.33960625976716e-08 pu0=3.97213309664079e-14
+  a0=0.622829915304962 la0=1.28828665004636e-07 wa0=7.07257249218472e-07 pa0=-5.26128667693621e-13
+  keta=0.864119589860614 lketa=-6.90887149197311e-07 wketa=-9.4427941131597e-07 pketa=7.0244945407795e-13
+  a1=0.0
+  a2=0.5
+  ags=-6.15309755878468 lags=5.12460335876992e-06 wags=6.18148466546483e-06 pags=-4.59840644263929e-12
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.32286479460111+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=1.77977861203966e-07 wvoff=2.35051964977664e-07 pvoff=-1.74855156746884e-13
+  nfactor={0.374925452622637+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=7.27068925794019e-07 wnfactor=1.367514896055e-06 pnfactor=-1.01729433117532e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-1.35975e-05 lcit=1.755418025e-11
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.700109518355951 leta0=-5.15734948324992e-07 weta0=-4.90965637275652e-07 peta0=3.65229337569358e-13
+  etab=-0.910363120933192 letab=6.74173227112201e-07 wetab=8.39923304757898e-07 petab=-6.248189464094e-13
+  dsub=3.82438852055279 ldsub=-2.64767601094122e-06 wdsub=-3.05911723105891e-06 pdsub=2.27567730818472e-12
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-3.98075515397057 lpclm=3.8187631549387e-06 wpclm=5.1726745452394e-06 ppclm=-3.84795259420359e-12
+  pdiblc1=0.708302091180901 lpdiblc1=-1.89075672785472e-07 wpdiblc1=-7.85766486912789e-07 ppdiblc1=5.84531689614424e-13
+  pdiblc2=-0.024688974080288 lpdiblc2=2.32785310547162e-08 wpdiblc2=8.77012095039316e-09 ppdiblc2=-6.52409297499747e-15
+  pdiblcb=-0.025
+  drout=-3.1722175498244 ldrout=2.76605522019637e-06 wdrout=5.33948090322375e-06 pdrout=-3.97203984390815e-12
+  pscbe1=-1139256544.40059 lpscbe1=1121.9324867456 wpscbe1=1125.20130441384 ppscbe1=-0.000837037250353453
+  pscbe2=2.54414976432243e-08 lpscbe2=-8.89491543669457e-15 wpscbe2=-6.87781478017134e-15 ppscbe2=5.11640641496949e-21
+  pvag=0.0
+  delta=0.01
+  alpha0=-0.000490713237445142 lalpha0=3.89185355455741e-10 walpha0=6.56295518466248e-10 palpha0=-4.88218236187042e-16
+  alpha1=0.0
+  beta0=-106.992489013277 lbeta0=0.000114887985192577 wbeta0=0.000151477303573597 pbeta0=-1.12683966128399e-10
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=1.17468972549849e-07 lagidl=-8.1616075399833e-14 wagidl=-1.25215775165977e-13 pagidl=9.31480151459701e-20
+  bgidl=1163596139.27439 lbgidl=464.940371993773 wbgidl=-486.62123819155 pbgidl=0.000361997539090692
+  cgidl=2677.50342077808 lcgidl=-0.00161240579471681 wcgidl=-0.00261901734729426 pcgidl=1.9482870046522e-9
+  egidl=10.4166325653881 legidl=-7.62833434482317e-06 wegidl=-9.60994511062446e-06 pegidl=7.14883816779354e-12
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.122566514528 lkt1=-3.8529071984262e-07 wkt1=-4.61137332949598e-07 pkt1=3.43040061981205e-13
+  kt2=-0.019032
+  at=-199191.70288 lat=0.163056707772432 wat=0.242703859447156 pat=-1.80547401042739e-7
+  ute=-0.552374226504 lute=-6.89912032903675e-07 wute=-7.1597638536911e-07 pute=5.32614833076081e-13
+  ua1=5.524e-10
+  ub1=-3.5909e-18
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=2.41e-6
+  sbref=2.41e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.62 pmos
* DC IV MOS Parameters
+  lmin=6e-07 lmax=8.0e-07 wmin=1e-06 wmax=1.5e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.0328630825+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=2.47518460717498e-8
+  k1=0.439924394999999 lk1=1.019407865595e-7
+  k2=0.0625425000195 lk2=-2.3267748848506e-8
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=6706.71609999996 lvsat=0.0394900683032101
+  ua=7.64635875649998e-10 lua=5.10014064223967e-16
+  ub=2.18208665e-18 lub=-9.19874491935e-25
+  uc=4.59868253100002e-13 luc=-1.74799580225109e-18
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.016805478645 lu0=-1.64088454015499e-10
+  a0=0.670912999999999 la0=9.30596583000004e-8
+  keta=-0.1003321935 lketa=2.656853244465e-8
+  a1=0.0
+  a2=0.5
+  ags=0.772544586889999 lags=-2.73818333974715e-8
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.0935342216534999+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=7.37884798823869e-9
+  nfactor={0.9112596485+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=3.2808991748085e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=-0.0232366091 leta0=2.236223588949e-08 peta0=6.31088724176809e-30
+  etab=-0.01522949275 letab=8.283321106725e-9
+  dsub=0.247220026019999 ldsub=1.33796321417223e-8
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=1.2962939877 lpclm=-1.06833701550031e-7
+  pdiblc1=0.60527969075 lpdiblc1=-1.12437309104925e-7
+  pdiblc2=0.00321937093564999 lpdiblc2=2.51751319735996e-9
+  pdiblcb=-0.025
+  drout=0.284514216564999 ldrout=1.94592459179297e-7
+  pscbe1=451591189.885 lpscbe1=-61.4991427894518
+  pscbe2=1.0408838377e-08 lpscbe2=2.28787979144971e-15
+  pvag=0.0
+  delta=0.01
+  alpha0=4.00715633235e-05 lalpha0=-5.66545783605163e-12
+  alpha1=0.0
+  beta0=45.4692438959999 lbeta0=1.47170208136561e-6
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-9.89710336e-08 lagidl=7.939364517504e-14 wagidl=1.26217744835362e-29 pagidl=1.20370621524202e-35
+  bgidl=2440736100.0 lbgidl=-485.12404479
+  cgidl=-730.092000000001 lcgidl=0.0009225044388
+  egidl=-2.696301033755 legidl=2.12637695957935e-06 pegidl=-3.02922587604869e-28
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.60520089 lkt1=-2.6259007929e-8
+  kt2=-0.019032
+  at=47195.0 lat=-0.0202303605
+  ute=-1.8567227 lute=2.8039279653e-7
+  ua1=5.534878e-10 lua1=-8.09214420000127e-19
+  ub1=-8.27197535e-18 lub1=3.482251952865e-24
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=2.02e-6
+  sbref=2.01e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.63 pmos
* DC IV MOS Parameters
+  lmin=5e-07 lmax=6e-07 wmin=1e-06 wmax=1.5e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.990437427040082+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=1.6765320670989e-09 wvth0=1.85876122539671e-07 pvth0=-1.01098023049327e-13
+  k1=0.538681698734559 lk1=4.82266890582729e-08 wk1=3.55316161784459e-07 pk1=-1.93256460394566e-13
+  k2=-0.0197473355697587 lk2=2.14896927284918e-08 wk2=-4.67861329030411e-08 pk2=2.5446977685964e-14
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=521840.96238278 lvsat=-0.240691448249994 wvsat=-0.659622254226451 pvsat=3.58768544073767e-7
+  ua=-2.64636689744616e-09 lua=2.36525847251097e-15 wua=5.29627559355234e-15 pua=-2.88064429533312e-21
+  ub=7.80258233036177e-18 lub=-3.97686209248377e-24 wub=-1.0053061863633e-23 pub=5.46786034763002e-30
+  uc=-1.71278180753186e-11 luc=7.81794679177577e-18 wuc=2.6019658711747e-17 puc=-1.41520923733192e-23
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0094808536597587 lu0=3.81977507545722e-09 wu0=5.25680730714581e-09 pu0=-2.85917749435662e-15
+  a0=0.193828088623521 la0=3.52546141597667e-07 wa0=1.08101489504035e-06 pa0=-5.87964001412444e-13
+  keta=0.254075759517144 lketa=-1.66193953201375e-07 wketa=-4.52283346250884e-07 pketa=2.45996912025856e-13
+  a1=0.0
+  a2=0.5
+  ags=-5.73785969588298 lags=3.51362705600275e-06 wags=8.33830298509563e-06 pags=-4.53520299359352e-12
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.202059890659656+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=6.64059593606869e-08 wvoff=2.4557010517941e-07 pvoff=-1.33565580207081e-13
+  nfactor={-0.848494756195077+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.2852203381945e-06 wnfactor=3.56507777823336e-06 pnfactor=-1.93904580358113e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-3.04435514400001e-05 lcit=2.1997247628216e-11 wcit=5.70697336627783e-11 pcit=-3.10402281391851e-17
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.619774921666033 leta0=-3.27371735694155e-07 weta0=-1.10873937165372e-06 peta0=6.03043344242461e-13
+  etab=0.0864104513594721 letab=-4.69986444944169e-08 wetab=-3.44587051855855e-08 petab=1.874208975044e-14
+  dsub=0.300745533230177 ldsub=-1.57328912298931e-08 wdsub=-5.21584265232269e-08 pdsub=2.83689681859832e-14
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-1.8009477350913 lpclm=1.57775607147616e-06 wpclm=4.49968700579042e-06 ppclm=-2.44737976244941e-12
+  pdiblc1=0.899469101041139 lpdiblc1=-2.72446929362276e-07 wpdiblc1=6.18368826550975e-07 ppdiblc1=-3.36330804761075e-13
+  pdiblc2=0.0108465546776569 lpdiblc2=-1.63091203991761e-09 wpdiblc2=2.06039190447184e-08 ppdiblc2=-1.12064715684223e-14
+  pdiblcb=-1.6427420576 lpdiblcb=8.79889905128641e-07 wpdiblcb=2.28278934651113e-06 ppdiblcb=-1.2416091255674e-12
+  drout=-0.94560258431 ldrout=8.63652987175208e-7
+  pscbe1=4039186262.82716 lpscbe1=-2012.79210296269 wpscbe1=-5238.04871396981 ppscbe1=0.00284897469552818
+  pscbe2=-5.93000950364422e-08 lpscbe2=4.02025686750209e-14 wpscbe2=1.03454393544843e-13 ppscbe2=-5.62688446490402e-20
+  pvag=0.0
+  delta=0.01
+  alpha0=-3.42222855691506e-05 lalpha0=3.4742966576661e-11 walpha0=1.61956271628785e-10 palpha0=-8.8088016138896e-17
+  alpha1=0.0
+  beta0=-5.70284798958539 lbeta0=2.93042028579355e-05 wbeta0=8.98794887918049e-05 pbeta0=-4.88854539538627e-11
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=2.49794487698178e-07 lagidl=-1.10299921859039e-13 wagidl=-4.48305585814589e-14 pagidl=2.43833408124555e-20
+  bgidl=3840351035.44961 lbgidl=-1246.37460818104 wbgidl=-4099.88966633399 pbgidl=0.00222992998951906
+  cgidl=1416.8319424 lcgidl=-0.000245207493471359 wcgidl=0.00228278934651113 pcgidl=-1.2416091255674e-9
+  egidl=-0.352356484516434 legidl=8.51505519248489e-07 wegidl=5.78611927087391e-06 pegidl=-3.14707027142832e-12
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.499598691359999 lkt1=-8.36960437692964e-08 wkt1=-3.42418401976669e-07 pkt1=1.86241368835111e-13
+  kt2=-0.019032
+  at=-159.841152000008 lat=0.00552593760257282 wat=0.0456557869302226 pat=-2.48321825113481e-8
+  ute=-0.8884720293056 lute=-2.46238743260684e-07 wute=-8.99419002525384e-07 pute=4.89193995473556e-13
+  ua1=5.52e-10
+  ub1=-5.80514400000002e-19 lub1=-7.01133657839997e-25
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=1.81e-6
+  sbref=1.81e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.64 pmos
* DC IV MOS Parameters
+  lmin=2.0e-05 lmax=1.0e-04 wmin=7.5e-07 wmax=1.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.019777265888+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} wvth0=9.77448013749257e-9
+  k1=0.62142183072 wk1=-3.33204486816693e-8
+  k2=0.022422366410784 wk2=3.91906540329634e-9
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=-184795.410496 wvsat=0.241396170297264
+  ua=1.6719378577344e-09 wua=5.4580822370722e-16
+  ub=1.25092521248e-18 wub=-8.81727014029678e-25
+  uc=-7.8082945127488e-11 wuc=3.00428103480018e-17
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.01756796441696 wu0=1.14154459796541e-9
+  a0=1.027397144704 wa0=-9.96385014952353e-8
+  keta=-0.0094623107328 wketa=1.16657709701115e-9
+  a1=0.0
+  a2=0.5
+  ags=0.24006319987392 wags=-7.6464478783849e-8
+  b0=2.508198224e-07 wb0=-2.2852093690935e-13
+  b1=-8.7777682496e-07 wb1=7.99738954113756e-13
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.10410066537376+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} wvoff=-3.26123590310883e-9
+  nfactor={1.54470873312+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} wnfactor=-2.39242267106999e-8
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.22192e-06 wcit=1.204643842432e-11
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-2.3266099098 wpclm=2.19586997012914e-6
+  pdiblc1=0.39
+  pdiblc2=0.0091183795479744 wpdiblc2=-5.17531040564768e-9
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=222383306.46784 wpscbe1=2.12677461093688
+  pscbe2=1.5010196982176e-08 wpscbe2=-1.04538992646255e-17
+  pvag=0.0
+  delta=0.01
+  alpha0=0.000183938006643392 walpha0=-1.09053968856232e-10
+  alpha1=0.0
+  beta0=42.617242287328 wbeta0=-3.2596867311274e-6
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-8.5593472e-09 wagidl=2.60203069965312e-14
+  bgidl=1040444304.0 wbgidl=437.285714802816
+  cgidl=1928.8768 wcgidl=-0.0004818575369728
+  egidl=2.6592854993344 wegidl=-1.03805750032237e-6
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.52955616 wkt1=-2.40928768486399e-8
+  kt2=-0.019032
+  at=-378712.3344 wat=0.482700787662502
+  ute=-1.9413867488 wute=3.51033215684685e-7
+  ua1=2.2096e-11
+  ub1=-4.8666835296e-18 wub1=1.63084683388444e-24
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.65 pmos
* DC IV MOS Parameters
+  lmin=8e-06 lmax=2.0e-05 wmin=7.5e-07 wmax=1.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.02687928850364+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=1.41642028844068e-07 wvth0=1.62451045345126e-08 pvth0=-1.29049485911713e-13
+  k1=0.645632077891384 lk1=-4.82846748561366e-07 wk1=-5.53783080385286e-08 pk1=4.39919741227266e-13
+  k2=0.0195748194584279 lk2=5.67911916630944e-08 wk2=6.51345404140014e-09 pk2=-5.17422275594788e-14
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=-360191.036315931 lvsat=3.49807282179012 wvsat=0.4011984233993 pvsat=-3.1870801556417e-6
+  ua=1.27536000458576e-09 lua=7.90930904541121e-15 wua=9.07128719399534e-16 pua=-7.20613983403796e-21
+  ub=1.89157771843166e-18 lub=-1.27771095134492e-23 wub=-1.46542294959221e-24 pub=1.16411733692655e-29
+  uc=-9.99116987315257e-11 luc=4.35350479003567e-16 wuc=4.99309004416261e-17 puc=-3.96646080018233e-22
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0167385315021174 lu0=1.65421271103297e-08 wu0=1.89723760894686e-09 pu0=-1.50714658417129e-14
+  a0=1.09979331115518 la0=-1.4438619040856e-06 wa0=-1.65598359164236e-07 pa0=1.31549680536477e-12
+  keta=-0.0103099319678242 lketa=1.69048731491984e-08 wketa=1.93884141375672e-09 pketa=-1.5401962306742e-14
+  a1=0.0
+  a2=0.5
+  ags=0.295621393248623 lags=-1.10804705284573e-06 wags=-1.27083326534767e-07 pags=1.00953723765954e-12
+  b0=4.16860454663613e-07 lb0=-3.31149776580228e-12 wb0=-3.79799892802199e-13 pb0=3.01709236843139e-18
+  b1=-1.45885776827665e-06 lb1=1.15890202254128e-11 wb1=1.32915947724578e-12 pb1=-1.05587099712927e-17
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.101731089620061+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=-4.72585818741972e-08 wvoff=-5.42014689400093e-09 pvoff=4.3057104911254e-14
+  nfactor={1.56209179562267+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-3.46686060246875e-07 wnfactor=-3.9761865424627e-08 pnfactor=3.15864282746692e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-1.69747208573333e-05 lcit=1.7456498501857e-10 wcit=2.0021080274233e-11 pcit=-1.59045459590479e-16
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-3.92210327307793 lpclm=3.18203600878788e-05 wpclm=3.64951759143821e-06 ppclm=-2.8991402794626e-11
+  pdiblc1=0.39
+  pdiblc2=0.0128786993835922 lpdiblc2=-7.49954427695782e-08 wpdiblc2=-8.60132276659974e-09 ppdiblc2=6.83280479255916e-14
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=220838016.98208 lpscbe1=30.8190989750583 wpscbe1=3.5346816802554 ppscbe1=-2.80791577997805e-5
+  pscbe2=1.501779266276e-08 lpscbe2=-1.51487493999108e-16 wpscbe2=-1.73742934619766e-17 ppscbe2=1.38019649832622e-22
+  pvag=0.0
+  delta=0.01
+  alpha0=0.000263175341237937 lalpha0=-1.58030147742015e-09 walpha0=-1.81246787455984e-10 palpha0=1.43980635487159e-15
+  alpha1=0.0
+  beta0=44.9856924308367 lbeta0=-4.7236132817124e-05 wbeta0=-5.41757218307763e-06 pbeta0=4.30366516651504e-11
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-2.746539705184e-08 lagidl=3.77060367640112e-13 wagidl=4.32455333923432e-14 pagidl=-3.43538192715435e-19
+  bgidl=722717632.878801 lbgidl=6336.7089561741 wbgidl=726.765213954657 pbgidl=-0.0057733501831344
+  cgidl=2278.98883429333 lcgidl=-0.00698259940074281 wcgidl=-0.000800843210969318 pcgidl=6.36181838361917e-9
+  egidl=3.41352590290795 legidl=-1.50424951848304e-05 wegidl=-1.72524291505662e-06 pegidl=1.37051571929183e-11
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.512050558285334 lkt1=-3.49129970037136e-07 wkt1=-4.00421605484654e-08 pkt1=3.18090919180956e-13
+  kt2=-0.019032
+  at=-729437.064753346 lat=6.99481894969411 wat=0.802244686588515 pat=-6.3729515657905e-6
+  ute=-2.19644336578269 lute=5.08682366344113e-06 wute=5.83414279191148e-07 pute=-4.63458469246656e-12
+  ua1=2.2096e-11
+  ub1=-6.05163770966579e-18 lub1=2.3632607671814e-23 wub1=2.71045384752566e-24 pub1=-2.15315743193591e-29
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.66 pmos
* DC IV MOS Parameters
+  lmin=4e-06 lmax=8e-06 wmin=7.5e-07 wmax=1.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.03907157288229+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=2.38496316719585e-07 wvth0=1.72033523524571e-08 pvth0=-1.36661710752683e-13
+  k1=0.476027341039248 lk1=8.64476320518317e-07 wk1=8.09569522468553e-08 pk1=-6.43113932953795e-13
+  k2=0.0556525217151932 lk2=-2.29806467294423e-07 wk2=-2.01849175620944e-08 pk2=1.60346966621522e-13
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=197394.704295728 lvsat=-0.931332543054834 wvsat=-0.142814905196037 pvsat=1.1345073253868e-6
+  ua=3.74709124767939e-09 lua=-1.17258767766003e-14 wua=-1.12350077163333e-15 pua=8.92497777977804e-21
+  ub=-9.16919875105361e-19 lub=9.53331451984947e-24 wub=1.0319160814564e-24 pub=-8.19743815948146e-30
+  uc=-6.72378394645289e-11 luc=1.75792608372471e-16 wuc=6.50158917161398e-18 puc=-5.16479742203841e-23
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0228839163143147 lu0=-3.22761952992841e-08 wu0=-2.99488462370012e-09 pu0=2.37910639622114e-14
+  a0=0.901926900755534 la0=1.27969073488119e-07 wa0=3.76064997365022e-08 pa0=-2.98742273256795e-13
+  keta=-0.00100743740508521 lketa=-5.69932134077437e-08 wketa=-5.05862176671591e-09 pketa=4.01851854526146e-14
+  a1=0.0
+  a2=0.5
+  ags=0.0445047894028949 lags=8.86798136444342e-07 wags=9.44870491759308e-08 pags=-7.50595669948677e-13
+  b0=-2.4730207439084e-07 lb0=1.96454294875339e-12 wb0=2.25315930769197e-13 pb0=-1.78988722243742e-18
+  b1=8.65466004989936e-07 lb1=-6.87517539703955e-12 wb1=-7.88522615282311e-13 pb1=6.26394480354115e-18
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.149332742164339+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=3.30884185772296e-07 wvoff=2.84186909501103e-08 pvoff=-2.25755239038582e-13
+  nfactor={1.25037304554145+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=2.12957651852328e-06 wnfactor=1.83697215881728e-07 pnfactor=-1.45927231324286e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=7.01250000000132e-08 lcit=3.91624340125e-11
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-0.522872595818586 lpclm=4.81721151079827e-06 wpclm=-1.93193575653167e-07 ppclm=1.53471044563119e-12
+  pdiblc1=0.39
+  pdiblc2=0.005556006565935 lpdiblc2=-1.6824703295391e-8
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=225793653.74242 lpscbe1=-8.54798388541258 wpscbe1=-1.28675944521933 ppscbe1=1.0221888356878e-5
+  pscbe2=1.49562706494802e-08 lpscbe2=3.37237227294089e-16 wpscbe2=3.08933440132141e-17 ppscbe2=-2.45413635506642e-22
+  pvag=0.0
+  delta=0.01
+  alpha0=0.000177066895447731 lalpha0=-8.96264594907328e-10 walpha0=-4.50835037833161e-11 palpha0=3.58138845704285e-16
+  alpha1=-3.5932715144e-10 lalpha1=2.85445895832422e-15 walpha1=2.37549742508378e-16 palpha1=-1.88707139951231e-21
+  beta0=165.011521548047 lbeta0=-0.00100070931674133 wbeta0=-8.23977175656403e-05 pbeta0=6.5455922856969e-10
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-7.09690240319974e-10 lagidl=1.64515708300078e-13 wagidl=6.6513927902346e-15 pagidl=-5.28379991863447e-20
+  bgidl=2166460677.20624 lbgidl=-5132.24141365865 wbgidl=-545.414208799236 pbgidl=0.00433271593328025
+  cgidl=4141.2312321952 lcgidl=-0.0217760667854354 wcgidl=-0.00168185217695932 pcgidl=1.33604655085471e-8
+  egidl=-1.32843888229237 legidl=2.26271988723224e-05 wegidl=2.16389144015372e-06 pegidl=-1.71897372114371e-11
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.510207534856 lkt1=-3.63770763857422e-07 wkt1=-2.37549742508382e-08 pkt1=1.88707139951232e-13
+  kt2=-0.019032
+  at=427107.161632776 lat=-2.19265273029461 wat=-0.313066805651792 pat=2.48697139741727e-6
+  ute=-1.6997565575 lute=1.14119332712424e-06 wute=8.470329472543e-22
+  ua1=2.2096e-11
+  ub1=-3.7441064775e-18 lub1=5.30181031661224e-24
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.67 pmos
* DC IV MOS Parameters
+  lmin=2e-06 lmax=4e-06 wmin=7.5e-07 wmax=1.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.925980967666947+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-2.07521721189188e-07 wvth0=-7.03846935926389e-08 pvth0=2.08776783650177e-13
+  k1=0.707645557692672 lk1=-4.90027641411201e-08 wk1=-8.3138875452899e-08 pk1=4.06360191126618e-15
+  k2=-0.00652088613447346 lk2=1.53992359238771e-08 wk2=1.92599983652764e-08 pk2=4.78016269556425e-15
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=-52850.9215919964 lvsat=0.0556111808837638 wvsat=0.245506999821763 pvsat=-3.96995435812902e-7
+  ua=8.70283729668738e-10 lua=-3.80035606318085e-16 wua=1.33574306018037e-15 pua=-7.74033968512046e-22
+  ub=-1.80111578247041e-20 lub=5.98810842976629e-24 wub=1.49034274155773e-25 pub=-4.71544059966853e-30
+  uc=-8.25156209799935e-12 luc=-5.68433709333848e-17 wuc=-3.52974798576905e-17 puc=1.1320337412429e-22
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0119089625623944 lu0=1.10079248029142e-08 wu0=6.50822321379846e-09 pu0=-1.36882430380992e-14
+  a0=0.30185508905808 la0=2.49459229164171e-06 wa0=4.68262576327908e-07 pa0=-1.99720677372564e-12
+  keta=0.280856502761671 lketa=-1.16863640703141e-06 wketa=-1.71812327846167e-07 pketa=6.97845126859363e-13
+  a1=0.0
+  a2=0.5
+  ags=-0.801841753518978 lags=4.22470426707392e-06 wags=4.14414570448918e-07 pags=-2.01235782109721e-12
+  b0=5.49118282282528e-07 lb0=-1.1764592959307e-12 wb0=-5.00299470514482e-13 pb0=1.07186735868528e-18
+  b1=-1.08611796883453e-06 lb1=8.21676637326751e-13 wb1=9.89557736933263e-13 pb1=-7.48626297561853e-19
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.0185031232293883+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=-1.85094748345258e-07 wvoff=-8.12461759045913e-08 pvoff=2.06752029349675e-13
+  nfactor={2.43699875477211+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-2.55035661611152e-06 wnfactor=-7.67030176594163e-07 pnfactor=2.2903014499428e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=2.08178259339994e-05 lcit=-4.26644237011002e-11 wcit=-7.15162145366326e-12 pcit=2.82052798511025e-17
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.311968541728 leta0=-9.14860731721059e-07 weta0=-1.40502429918214e-07 peta0=5.54127533354444e-13
+  etab=-0.135741180949338 letab=2.59276643546093e-07 wetab=-1.51742624311673e-09 petab=5.98457736022796e-15
+  dsub=0.995402871054915 ldsub=-1.71718538315348e-06 wdsub=-1.31031887046648e-07 pdsub=5.16776659323276e-13
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-2.35599842986424 lpclm=1.20468764876909e-05 wpclm=2.10233161936165e-06 ppclm=-7.51861137098776e-12
+  pdiblc1=0.789328332407172 lpdiblc1=-1.57491101018064e-06 wpdiblc1=-3.64630782104309e-07 ppdiblc1=1.43806734154119e-12
+  pdiblc2=0.00319363714014225 lpdiblc2=-7.50775451700703e-09 wpdiblc2=-1.73439618383505e-09 ppdiblc2=6.84028510942704e-15
+  pdiblcb=-0.025
+  drout=-0.0611043172974277 ldrout=2.44957331698933e-06 wdrout=4.96813407469059e-07 pdrout=-1.95938239771722e-12
+  pscbe1=58125008.024431 lpscbe1=652.720387961767 wpscbe1=76.9600247839703 ppscbe1=-0.000298375603964623
+  pscbe2=1.465527626283e-08 lpscbe2=1.52432898880398e-15 wpscbe2=5.32875796359405e-16 ppscbe2=-2.22518222931475e-21
+  pvag=0.0
+  delta=0.01
+  alpha0=-0.00123163192355892 lalpha0=4.659502677373e-09 walpha0=8.38968361789335e-10 palpha0=-3.12847330692769e-15
+  alpha1=9.7567520576e-10 lalpha1=-2.41065683823686e-15 walpha1=-7.09270201547113e-16 palpha1=1.84709177784815e-21
+  beta0=-363.285181264348 lbeta0=0.00108284004948047 wbeta0=0.000287368677806634 pbeta0=-8.03762458139024e-10
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-6.05565665979186e-08 lagidl=4.00545803966812e-13 wagidl=8.01182167550174e-14 pagidl=-3.42583806221051e-19
+  bgidl=-1337799124.93296 lbgidl=8688.20881999814 wbgidl=2442.22762269516 pbgidl=-0.0074502446859505
+  cgidl=-1404.8969704864 lcgidl=9.73082331205124e-05 wcgidl=0.00142008740671668 pcgidl=1.12672598448737e-9
+  egidl=5.87086179154466 legidl=-5.76612305522352e-06 wegidl=-3.04594094866848e-06 pegidl=3.35732074683877e-12
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.675056778238401 lkt1=2.86378167118426e-07 wkt1=1.24786284956693e-07 pkt1=-3.97124732237351e-13
+  kt2=-0.019032
+  at=-224284.912972188 lat=0.37637247273991 wat=0.58406718378607 pat=-1.05123534352672e-6
+  ute=-1.5350444853248 lute=4.91585385672478e-07 wute=1.07718529603964e-07 pute=-4.24831108905073e-13
+  ua1=-1.27600843180365e-09 lua1=5.11959406859041e-15 wua1=5.17423615245476e-16 pua1=-2.04066699616663e-21
+  ub1=-4.040415987752e-18 lub1=6.4704253940951e-24 wub1=1.84994866058982e-24 pub1=-7.29601252250018e-30
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.68 pmos
* DC IV MOS Parameters
+  lmin=1e-06 lmax=2e-06 wmin=7.5e-07 wmax=1.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.09131144872361+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=1.13864200936864e-07 wvth0=7.8298516990427e-08 pvth0=-8.02485094022407e-14
+  k1=0.672839661739296 lk1=1.86564170026462e-08 wk1=-7.47036243772023e-08 pk1=-1.23336826547814e-14
+  k2=0.00468361082748295 lk2=-6.38118572046996e-09 wk2=1.84133243941132e-08 pk2=6.42601222810835e-15
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=-31488.202622176 lvsat=0.0140841914783296 wvsat=0.0265216532615869 pvsat=2.86901793654239e-8
+  ua=3.04871135479424e-09 lua=-4.61468106679953e-15 wua=-6.32266868840042e-16 pua=3.05158053251074e-21
+  ub=6.79663728614944e-19 lub=4.63189821801626e-24 wub=-6.90957425099641e-25 pub=-3.08258073548593e-30
+  uc=-7.22217563773396e-11 luc=6.75082897262247e-17 wuc=4.58964264281977e-17 puc=-4.46294603048483e-23
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0229296421925194 lu0=-1.04151743300859e-08 wu0=-3.95879681231302e-09 pu0=6.65859719065886e-15
+  a0=1.74898545679898 la0=-3.18484430209837e-07 wa0=-6.67472572907981e-07 pa0=2.10548782874003e-13
+  keta=-0.40333787994783 lketa=1.61369053517586e-07 wketa=2.39209713052726e-07 pketa=-1.01140618443996e-13
+  a1=0.0
+  a2=0.5
+  ags=1.29038342995906 lags=1.57627732910969e-07 wags=-5.67194955442691e-07 pags=-1.0420706371651e-13
+  b0=-1.1676572297685e-07 lb0=1.17952621893003e-13 wb0=1.06384783141316e-13 pb0=-1.07466161996228e-19
+  b1=-2.52898387291081e-06 lb1=3.62646366826064e-12 wb1=2.30414709067355e-12 pb1=-3.3040565422976e-18
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.136125546200861+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=4.35514796689877e-08 wvoff=3.99245316178764e-08 pvoff=-2.87917090032491e-14
+  nfactor={1.01418613022125+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=2.15448844752891e-07 wnfactor=6.09387145233145e-07 pnfactor=-3.853161819573e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=5.56401842000122e-06 lcit=-1.30125472746391e-11 wcit=2.93260967861087e-12 pcit=8.60254295307484e-18
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=-0.354312670107625 leta0=3.80323315966213e-07 weta0=2.88807388357972e-07 peta0=-2.80407822392635e-13
+  etab=-0.0127208345764263 letab=2.01373922317903e-08 wetab=1.11183266135932e-08 petab=-1.85780626179304e-14
+  dsub=-0.0527879742955222 ldsub=3.20392801123238e-07 wdsub=2.43774974713033e-07 pdsub=-2.11810399251368e-13
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=6.02766372521723 lpclm=-4.25012437557193e-06 wpclm=-3.21087975734541e-06 ppclm=2.8097402241931e-12
+  pdiblc1=0.205011082161199 lpdiblc1=-4.39056707427497e-07 wpdiblc1=2.2583617015028e-07 ppdiblc1=2.90258633053489e-13
+  pdiblc2=-0.0031546203331016 lpdiblc2=4.83262318523169e-09 wpdiblc2=3.42796451717373e-09 ppdiblc2=-3.19482785726393e-15
+  pdiblcb=-0.025
+  drout=-0.0462253258064109 ldrout=2.42065004542994e-06 wdrout=3.12081510106195e-07 pdrout=-1.60028206243355e-12
+  pscbe1=390001432.644157 lpscbe1=7.58580614348102 wpscbe1=-73.9534264565218 ppscbe1=-5.01494609823081e-6
+  pscbe2=1.6641741562704e-08 lpscbe2=-2.33716090762115e-15 wpscbe2=-1.40666325230536e-15 ppscbe2=1.54508772738472e-21
+  pvag=0.0
+  delta=0.01
+  alpha0=0.00200997751154271 lalpha0=-1.64186190352105e-09 walpha0=-1.32878802686124e-09 palpha0=1.08542833697015e-15
+  alpha1=-2.644384e-10 walpha1=2.409287684864e-16
+  beta0=212.307416770732 lbeta0=-3.6054401839918e-05 wbeta0=-0.000138372295997464 pbeta0=2.38354208387625e-11
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=2.7662089543082e-07 lagidl=-2.54893464470853e-13 wagidl=-1.82803155748133e-13 pagidl=1.68509049787823e-19
+  bgidl=3347013878.40576 lbgidl=-418.599177191996 wbgidl=-1532.76025095853 pbgidl=0.00027673424164492
+  cgidl=-1391.45882137651 lcgidl=7.11858150658001e-05 wcgidl=0.00244571049620026 pcgidl=-8.66982739159773e-10
+  egidl=7.57282921067541 legidl=-9.07457752127178e-06 wegidl=-4.40498521749091e-06 pegidl=5.99916690100269e-12
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.4486168446752 lkt1=-1.53798419735078e-07 wkt1=-1.31811406452604e-07 pkt1=1.01675520093182e-13
+  kt2=-0.019032
+  at=-87931.9695867263 lat=0.111315986092911 wat=0.0841328550350264 pat=-7.94130018675615e-8
+  ute=-1.1239213693504 lute=-3.07596839470157e-07 wute=-2.15437059207927e-07 pute=2.03351040186364e-13
+  ua1=2.1177509180073e-09 lua1=-1.47753473150709e-15 wua1=-1.03484723049095e-15 pua1=9.76792300860409e-22
+  ub1=2.00571126550399e-18 lub1=-5.28264137350922e-24 wub1=-3.69989732117963e-24 pub1=3.49233308146145e-30
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=2.81e-6
+  sbref=2.81e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.69 pmos
* DC IV MOS Parameters
+  lmin=8.0e-07 lmax=1e-06 wmin=7.5e-07 wmax=1.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.642138254675405+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-3.10110376925236e-07 wvth0=-2.33074130445234e-07 pvth0=2.1365613251228e-13
+  k1=0.954357487341278 lk1=-2.47068258583066e-07 wk1=-2.6081393281137e-07 pk1=1.6333583747623e-13
+  k2=-0.0576453864965935 lk2=5.24511548537258e-08 wk2=5.66723945371764e-08 pk2=-2.9686724079929e-14
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=-64616.1888341903 lvsat=0.0453536976638498 wvsat=0.0536308868562966 pvsat=3.10177377537734e-9
+  ua=-7.68226391551368e-09 lua=5.51428649084411e-15 wua=6.44574590026487e-15 pua=-3.62935572024738e-21
+  ub=1.12908557451704e-17 lub=-5.38400592641044e-24 wub=-8.14214550823122e-24 pub=3.95059569618196e-30
+  uc=-5.20166542109638e-12 luc=4.24802587262675e-18 wuc=1.58971237738913e-18 puc=-2.80835291229005e-24
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=-0.00491747055040193 lu0=1.58697153879576e-08 wu0=1.40359182827765e-08 pu0=-1.03266143875961e-14
+  a0=3.14376150837266 la0=-1.63501354529023e-06 wa0=-1.58955344149913e-06 pa0=1.08090091473719e-12
+  keta=-0.541668943041296 lketa=2.91939743971508e-07 wketa=3.36528897856829e-07 pketa=-1.93000196980588e-13
+  a1=0.0
+  a2=0.5
+  ags=1.15819889390733 lags=2.82396716490194e-07 wags=-4.79808287397039e-07 pags=-1.86691339684802e-13
+  b0=3.86872798757712e-08 lb0=-2.87794674995862e-14 wb0=-3.52478259456957e-14 pb0=2.6220857721003e-20
+  b1=6.19677895310065e-06 lb1=-4.60978386321157e-12 wb1=-5.64586051705419e-12 pb1=4.19995563863661e-18
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.036165341803603+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=-5.08009572615841e-08 wvoff=-2.61587596683333e-08 pvoff=3.35843096418042e-14
+  nfactor={2.51063049750819+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.19704499352925e-06 wnfactor=-5.78317427520043e-07 pnfactor=7.35758164264435e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-7.59983514400001e-05 lcit=6.39741736362161e-11 wcit=5.68531661435783e-11 pcit=-4.22930702942079e-17
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.492114027217527 leta0=-4.18618843638998e-07 weta0=-3.01461777281398e-07 peta0=2.76747243054367e-13
+  etab=0.053458904541402 letab=-4.23296635215278e-08 wetab=-3.82110873639027e-08 petab=2.79839712354279e-14
+  dsub=0.86556318561798 ldsub=-5.46438858719117e-07 wdsub=-3.63343303701143e-07 pdsub=3.61248543743773e-13
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=3.08735930694654 lpclm=-1.47477103516623e-06 wpclm=-1.26705626764433e-06 ppclm=9.74965232264255e-13
+  pdiblc1=-2.00721384547582 lpdiblc1=1.64906240176909e-06 wpdiblc1=1.68832922091141e-06 ppdiblc1=-1.09018855755994e-12
+  pdiblc2=-0.0602654488468101 lpdiblc2=5.87395342193212e-08 wpdiblc2=4.11837048042724e-08 ppdiblc2=-3.88324711142564e-14
+  pdiblcb=-0.025
+  drout=8.67105620132828 ldrout=-5.80759198803249e-06 wdrout=-5.45087843835644e-06 pdrout=3.83937583292033e-12
+  pscbe1=-386582947.288653 lpscbe1=740.60380236206 wpscbe1=439.44340077954 ppscbe1=-0.000489610211326349
+  pscbe2=2.6826825714991e-08 lpscbe2=-1.19508618389648e-14 wpscbe2=-8.13998164504566e-15 ppscbe2=7.90066695829225e-21
+  pvag=0.0
+  delta=0.01
+  alpha0=0.000836834338293315 lalpha0=-5.34532062290952e-10 walpha0=-5.53227767598758e-10 palpha0=3.53377008252299e-16
+  alpha1=-2.644384e-10 walpha1=2.409287684864e-16
+  beta0=208.054347214226 lbeta0=-3.20399294855316e-05 wbeta0=-0.000135560608725936 pbeta0=2.1181469223167e-11
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-7.17183738800897e-08 lagidl=7.39039718317142e-14 wagidl=4.7152059416955e-14 pagidl=-4.85456778065036e-20
+  bgidl=-425642744.332806 lbgidl=3142.41140901093 wbgidl=961.327951707441 pbgidl=-0.00207743561285149
+  cgidl=-3346.89512158816 lcgidl=0.00191692213883558 wcgidl=0.00286978806706145 pcgidl=-1.26726955829565e-9
+  egidl=-2.88309891679771 legidl=7.94773038250096e-07 wegidl=2.50738704386906e-06 pegidl=-5.25421276494985e-13
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.572750051136001 lkt1=-3.66290861567287e-08 wkt1=-5.09769134801944e-08 pkt1=2.5375842176525e-14
+  kt2=-0.019032
+  at=-31162.8628800001 lat=0.0577316262724321 wat=0.0896134554385166 pat=-8.45861405884158e-8
+  ute=-1.338215 lute=-1.05325081500001e-7
+  ua1=5.524e-10
+  ub1=-3.5909e-18
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=2.41e-6
+  sbref=2.41e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.70 pmos
* DC IV MOS Parameters
+  lmin=6e-07 lmax=8.0e-07 wmin=7.5e-07 wmax=1.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.57816948656872+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=3.86203256480201e-07 wvth0=4.96826483521397e-07 pvth0=-3.29316934217497e-13
+  k1=0.200848202612479 lk1=3.13467298326687e-07 wk1=2.178213625795e-07 pk1=-1.92720958765038e-13
+  k2=0.101842014621781 lk2=-6.61915228382334e-08 wk2=-3.58056305560802e-08 pk2=3.91076787869446e-14
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=-293249.779558146 lvsat=0.2154342258034 wvsat=0.273289163368154 pvsat=-1.60302018121793e-7
+  ua=-1.10122784352354e-08 lua=7.99148429206512e-15 wua=1.07298995209905e-14 pua=-6.81633759870516e-21
+  ub=2.10580288149203e-17 lub=-1.26498059729974e-23 wub=-1.71977954026903e-23 pub=1.068709365267e-29
+  uc=8.72638351441749e-12 luc=-6.11304973050201e-18 wuc=-7.53158898852531e-18 puc=3.97698317381371e-24
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0114503740510774 lu0=3.69367578891711e-09 wu0=4.87901437510449e-09 pu0=-3.51479357067893e-15
+  a0=1.00033955641136 la0=-4.05219552262188e-08 wa0=-3.00139217840164e-07 pa0=1.21705673757283e-13
+  keta=-0.570923394583824 lketa=3.13702130473995e-07 wketa=4.28753760942668e-07 pketa=-2.61606272630144e-13
+  a1=0.0
+  a2=0.5
+  ags=5.4215167543229 lags=-2.88908543987295e-06 wags=-4.23565994585945e-06 pags=2.60728670904539e-12
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.367589868055089+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=1.95745747816897e-07 wvoff=2.49691003213903e-07 pvoff=-1.71620328966291e-13
+  nfactor={-2.67902178024871+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=2.66353733589411e-06 wnfactor=3.27109104860723e-06 pnfactor=-2.12781680112664e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-2.595701144e-05 lcit=2.6748420810216e-11 wcit=3.27602892949383e-11 pcit=-2.43703792065046e-17
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=-0.289685151083959 leta0=1.62961565099477e-07 weta0=2.42760200807417e-07 peta0=-1.28099486445902e-13
+  etab=-0.0128079221658944 letab=6.96622886602996e-09 wetab=-2.20628327289628e-09 petab=1.19999747212829e-15
+  dsub=-0.117527741347609 ldsub=1.84882481850585e-07 wdsub=3.32320231857559e-07 pdsub=-1.56255560358346e-13
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=1.97761146997746 lpclm=-6.49229619244932e-07 wpclm=-6.20745632833067e-07 ppclm=4.94174751028155e-13
+  pdiblc1=1.14089119122192 lpdiblc1=-6.92812935030361e-07 wpdiblc1=-4.8799349563396e-07 ppdiblc1=5.28777911278161e-13
+  pdiblc2=0.0244476836856485 lpdiblc2=-4.27856507157486e-09 wpdiblc2=-1.93410308332727e-08 ppdiblc2=6.19187972651345e-15
+  pdiblcb=-0.025
+  drout=4.03351920012437 ldrout=-2.3577282128369e-06 wdrout=-3.41570344450101e-06 pdrout=2.32540915499127e-12
+  pscbe1=1786640957.47623 lpscbe1=-876.057460392536 wpscbe1=-1216.3585030533 ppscbe1=0.000742140824934901
+  pscbe2=-6.92068717669786e-10 lpscbe2=8.52044372949154e-15 wpscbe2=1.01139920503253e-14 ppscbe2=-5.67846407369416e-21
+  pvag=0.0
+  delta=0.01
+  alpha0=0.000392466817447044 lalpha0=-2.0396706353341e-10 walpha0=-3.21065906450944e-10 palpha0=1.80671799744441e-16
+  alpha1=-9.83578628800001e-10 lalpha1=5.3496841620432e-16 walpha1=8.96134554385165e-16 palpha1=-4.87407584130092e-22
+  beta0=492.171800094041 lbeta0=-0.000243394902682826 wbeta0=-0.00040698891214181 pbeta0=2.23096984134236e-10
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-1.53779233443623e-07 lagidl=1.34949045261026e-13 wagidl=4.99355316447251e-14 pagidl=-5.06163027967418e-20
+  bgidl=11296947356.576 lbgidl=-5578.02336705513 wbgidl=-8068.85865102137 pbgidl=0.00464012020091847
+  cgidl=-6684.97549037729 lcgidl=0.00440012012517781 wcgidl=0.00542547052854878 pcgidl=-3.16844174139607e-9
+  egidl=-11.9184028836308 legidl=7.51613565917726e-06 wegidl=8.40222010701447e-06 pegidl=-4.91058759216886e-12
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.176780271584001 lkt1=-3.31191005165462e-07 wkt1=-3.90332311756344e-07 pkt1=2.77822322954152e-13
+  kt2=-0.019032
+  at=145552.86288 lat=-0.073727202120432 wat=-0.0896134554385165 pat=4.87407584130092e-8
+  ute=-1.8567227 lute=2.80392796530002e-7
+  ua1=5.53487800000001e-10 lua1=-8.09214420000522e-19
+  ub1=-8.27197535e-18 lub1=3.482251952865e-24
+  uc1=4.09098745700737e-10 luc1=-3.85562436926778e-16 wuc1=-4.72219914012958e-16 puc1=3.5128439403424e-22
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=2.02e-6
+  sbref=2.01e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.71 pmos
* DC IV MOS Parameters
+  lmin=5e-07 lmax=6e-07 wmin=7.5e-07 wmax=1.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.0961596996004701+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-4.19861866651829e-07 wvth0=-6.28896737819645e-07 pvth0=2.82963925869896e-13
+  k1=1.42396183499168 lk1=-3.51784206324359e-07 wk1=-4.5125902923886e-07 pk1=1.71191866344967e-13
+  k2=-0.192691250344499 lk2=9.40051199769265e-08 wk2=1.10782376072566e-07 pk2=-4.06215380183758e-14
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=-753433.33077003 lvsat=0.465728059307544 wvsat=0.502275053167901 pvsat=-2.84847443583876e-7
+  ua=2.06206028587491e-08 lua=-9.21363984373306e-15 wua=-1.59021674834381e-14 pua=7.66884364500355e-21
+  ub=-2.92004245700714e-17 lub=1.46857668230996e-23 wub=2.3660229711324e-23 pub=-1.15355862068423e-29
+  uc=2.28443773953897e-11 luc=-1.37918266023628e-17 wuc=-1.03988486928334e-17 puc=5.53648572698687e-24
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0294959328004253 lu0=-6.12130361485319e-09 wu0=-1.29788512375989e-08 pu0=6.19809953607045e-15
+  a0=1.38644615858688 la0=-2.50525336149485e-07 wa0=-5.57465803099354e-09 pa0=-3.85079903229251e-14
+  keta=-0.392122891580656 lketa=2.16452536890572e-07 wketa=1.36465659969717e-07 pketa=-1.02630774510956e-13
+  a1=0.0
+  a2=0.5
+  ags=10.331231612736 lags=-5.55947935136383e-06 wags=-6.30218182982186e-06 pags=3.73126796173254e-12
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={0.623869398165448+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=-3.43508947080454e-07 wvoff=-5.06930766151987e-07 pvoff=2.39906251391817e-13
+  nfactor={8.04289772241223+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-3.16811468160318e-06 wnfactor=-4.53583434345584e-06 pnfactor=2.11836991961646e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=0.00016280112576 lcit=-7.59171300128641e-11 wcit=-1.18994718755433e-10 pcit=5.81691696720924e-17
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=-1.67609071843309 leta0=9.1702755318067e-07 weta0=9.83014629578026e-07 peta0=-5.30723870254237e-13
+  etab=0.125754149340451 letab=-6.83976818262715e-08 wetab=-7.03045910412638e-08 petab=3.82386670673434e-14
+  dsub=-0.125462402745114 ldsub=1.89198144184687e-07 wdsub=3.36157919112116e-07 pdsub=-1.58342878456099e-13
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=6.09644639655989 lpclm=-2.88946393581312e-06 wpclm=-2.69559719798046e-06 ppclm=1.62268651731182e-12
+  pdiblc1=-0.75328143840188 lpdiblc1=3.37427558222022e-07 wpdiblc1=2.12418323203535e-06 ppdiblc1=-8.91985010901178e-13
+  pdiblc2=0.100061509046729 lpdiblc2=-4.54049246854666e-08 wpdiblc2=-6.06794690211258e-08 ppdiblc2=2.86758562568868e-14
+  pdiblcb=3.2104841152 lpdiblcb=-1.75977981025728e-06 wpdiblcb=-2.13896560662226e-06 ppdiblcb=1.16338339344185e-12
+  drout=-6.07797119889259 ldrout=3.14191141518842e-06 wdrout=4.67608051527174e-06 pdrout=-2.07571214072913e-12
+  pscbe1=-7289602666.61215 lpscbe1=4060.51144674914 wpscbe1=5083.56556448663 ppscbe1=-0.00268438787540007
+  pscbe2=1.62485305663535e-07 lpscbe2=-8.02317301964457e-14 wpscbe2=-9.86133978913032e-14 ppscbe2=5.34583633155576e-20
+  pvag=0.0
+  delta=0.01
+  alpha0=0.000258395852343585 lalpha0=-1.31045865613639e-10 walpha0=-1.04646943350957e-10 palpha0=6.29615257143573e-17
+  alpha1=0.0
+  beta0=174.052992371366 lbeta0=-7.03700831624633e-05 wbeta0=-7.38953383376964e-05 pbeta0=4.19273893421784e-11
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=7.022007498912e-07 lagidl=-3.30618467674784e-13 wagidl=-4.57016094440473e-13 pagidl=2.25114686630998e-19
+  bgidl=-6496302731.10401 lbgidl=4099.72535563403 wbgidl=5317.79423375793 pbgidl=-0.00264088030311299
+  cgidl=12648.666670656 lcgidl=-0.00611544784620821 wcgidl=-0.00795049034706401 pcgidl=4.10674337884972e-9
+  egidl=19.0579251309104 legidl=-9.33188914793175e-06 wegidl=-1.18985106678151e-05 pegidl=6.13097987626093e-12
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-2.12279915472 lkt1=7.27248665372208e-07 wkt1=1.13647304738877e-06 pkt1=-5.52607111884878e-13
+  kt2=-0.019032
+  at=96904.682304 lat=-0.0472674567051456 wat=-0.0427793121324452 pat=2.3267667868837e-8
+  ute=-3.6223325817088 lute=1.24070801119142e-06 wute=1.59139041132696e-06 pute=-8.65557244720734e-13
+  ua1=5.52e-10
+  ub1=-6.6657116265984e-18 lub1=2.60860511370687e-24 wub1=5.5441988523649e-24 pub1=-3.01548975580127e-30
+  uc1=-1.14579749140147e-09 luc1=4.60145626433114e-16 wuc1=9.44439828025916e-16 puc1=-4.19236839660704e-22
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=1.81e-6
+  sbref=1.81e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.72 pmos
* DC IV MOS Parameters
+  lmin=2.0e-05 lmax=1.0e-04 wmin=7e-07 wmax=7.5e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.004992+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+  k1=0.57102
+  k2=0.0283505
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=180350.0
+  ua=2.497549e-9
+  ub=-8.281e-20
+  uc=-3.2639e-11
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.01929471
+  a0=0.87668
+  keta=-0.0076977
+  a1=0.0
+  a2=0.5
+  ags=0.1244
+  b0=-9.485e-8
+  b1=3.3194e-7
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.10903374+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.50852+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.99495
+  pdiblc1=0.39
+  pdiblc2=0.00129
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=225600350.0
+  pscbe2=1.4994384e-8
+  pvag=0.0
+  delta=0.01
+  alpha0=1.8978653e-5
+  alpha1=0.0
+  beta0=37.686511
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=3.08e-8
+  bgidl=1701900000.0
+  cgidl=1200.0
+  egidl=1.0890786
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.566
+  kt2=-0.019032
+  at=351440.0
+  ute=-1.4104
+  ua1=2.2096e-11
+  ub1=-2.3998e-18
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.73 pmos
* DC IV MOS Parameters
+  lmin=8e-06 lmax=2.0e-05 wmin=7e-07 wmax=7.5e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.00230629980834+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-5.35633360526048e-8
+  k1=0.56186465525 lk1=1.8259328015953e-7
+  k2=0.0294273280825916 lk2=-2.14761515964003e-8
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=246677.59305 lvsat=-1.32283088302989
+  ua=2.64751884293833e-09 lua=-2.99098355057783e-15
+  ub=-3.2507909025e-19 lub=4.83179050903698e-24 wub=-1.83670992315982e-40
+  uc=-2.43842406291833e-11 luc=-1.64632095415631e-16
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0196083682715832 lu0=-6.25556920263095e-9
+  a0=0.849302672633335 la0=5.46010679268076e-7
+  keta=-0.00737716363499999 lketa=-6.39274520992324e-9
+  a1=0.0
+  a2=0.5
+  ags=0.103390118918166 lags=4.19018967307977e-7
+  b0=-1.57639909583334e-07 lb0=1.25227567773904e-12
+  b1=5.51681513833333e-07 lb1=-4.38250277774061e-12
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.109929818539917+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=1.78713007922409e-8
+  nfactor={1.50194642275+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.31102767316307e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.33099583333333e-05 lcit=-6.60134780041667e-11
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=1.59830161734375 lpclm=-1.2033184321142e-5
+  pdiblc1=0.39
+  pdiblc2=-0.000132002188645002 lpdiblc2=2.8360269450117e-8
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=226184716.523832 lpscbe1=-11.6545475146777
+  pscbe2=1.49915116181583e-08 lpscbe2=5.72864962118343e-17 wpscbe2=-2.52435489670724e-29
+  pvag=0.0
+  delta=0.01
+  alpha0=-1.09857298561001e-05 lalpha0=5.97606655243774e-10
+  alpha1=0.0
+  beta0=36.7908581207249 lbeta0=1.78628114589734e-5
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=3.794951e-08 lagidl=-1.42589112489e-13 wagidl=5.04870979341448e-29
+  bgidl=1822051487.5 lbgidl=-2396.28925155132
+  cgidl=1067.60166666667 lcgidl=0.00264053912016668
+  egidl=0.803855121271667 legidl=5.68846853741002e-6
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.572619916666666 lkt1=1.32026956008326e-07 wkt1=8.470329472543e-22
+  kt2=-0.019032
+  at=484070.030416666 lat=-2.64516006362696
+  ute=-1.31394781416666 lute=-1.9236327490414e-6
+  ua1=2.2096e-11
+  ub1=-1.95169784083332e-18 lub1=-8.93690465220408e-24
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.74 pmos
* DC IV MOS Parameters
+  lmin=4e-06 lmax=8e-06 wmin=7e-07 wmax=7.5e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.013049100575+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=3.17763989577253e-8
+  k1=0.598486034250001 lk1=-1.08323292478583e-7
+  k2=0.025120015752225 lk2=1.27407068248004e-8
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=-18632.7791499998 lvsat=0.784768182689687
+  ua=2.04763947118501e-09 lua=1.77439819069343e-15
+  ub=6.43997270749998e-19 lub=-2.86645519511093e-24
+  uc=-5.74032781124501e-11 luc=9.76678364476925e-17
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.01835373518525 lu0=3.71111057189243e-9
+  a0=0.958811982099999 la0=-3.23920324204192e-7
+  keta=-0.00865930909499998 lketa=3.79249010977054e-9
+  a1=0.0
+  a2=0.5
+  ags=0.1874296432455 lags=-2.48582609995927e-7
+  b0=9.35197287499998e-08 lb0=-7.42911373217127e-13
+  b1=-3.272845415e-07 lb1=2.59991566922185e-12
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.10634550438025+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=-1.06021324607301e-8
+  nfactor={1.52824073175+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-7.77765939488086e-8
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=7.01249999999793e-08 lcit=3.91624340125001e-11
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-0.81510485203125 lpclm=7.13867533092605e-06 wpclm=2.11758236813575e-22 ppclm=-1.61558713389263e-27
+  pdiblc1=0.39
+  pdiblc2=0.005556006565935 lpdiblc2=-1.68247032953911e-8
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=223847250.428501 lpscbe1=6.91404940003849
+  pscbe2=1.5003001145525e-08 lpscbe2=-3.39851602360616e-17
+  pvag=0.0
+  delta=0.01
+  alpha0=0.0001088718015683 lalpha0=-3.54529588638518e-10
+  alpha1=0.0
+  beta0=40.3734696378249 lbeta0=-1.05970961717175e-5
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=9.35147e-09 lagidl=8.4590857467e-14
+  bgidl=1341445537.5 lbgidl=1421.59635465374
+  cgidl=1597.195 lcgidl=-0.00156649736049999
+  egidl=1.944749036185 legidl=-3.37467863327002e-6
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.546140250000001 lkt1=-7.83248680249999e-8
+  kt2=-0.019032
+  at=-46450.0912499996 lat=1.56923873088087
+  ute=-1.6997565575 lute=1.14119332712427e-6
+  ua1=2.2096e-11
+  ub1=-3.7441064775e-18 lub1=5.30181031661227e-24
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.75 pmos
* DC IV MOS Parameters
+  lmin=2e-06 lmax=4e-06 wmin=7e-07 wmax=7.5e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.0324476436+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=1.08282312794046e-7
+  k1=0.581886401 lk1=-4.28559989039009e-8
+  k2=0.0226125504092 lk2=2.26298993911562e-8
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=318512.6925 lvsat=-0.54489984295075
+  ua=2.89078160014499e-09 lua=-1.55087005171188e-15
+  ub=2.074239895e-19 lub=-1.14465383118905e-24 wub=-1.83670992315982e-40
+  uc=-6.1643928498175e-11 luc=1.14392537503952e-16
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0217535588295 lu0=-9.69745389866518e-9
+  a0=1.010167613 la0=-5.26461796910697e-7
+  keta=0.020966369035 lketa=-1.13048221867136e-07 pketa=1.0097419586829e-28
+  a1=0.0
+  a2=0.5
+  ags=-0.1749818565465 lags=1.18073210403374e-06 pags=8.07793566946316e-28
+  b0=-2.07654517e-07 lb0=4.448897345963e-13 pb0=-3.85185988877447e-34
+  b1=4.10726267e-07 lb1=-3.107251584213e-13
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.1413993076029+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=1.27646562069078e-07 wvoff=2.11758236813575e-22
+  nfactor={1.2767585225+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=9.14044091112243e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.0994389999999998 leta0=-7.66654720999996e-8
+  etab=-0.1380365 letab=2.6832915235e-7
+  dsub=0.797198847665502 ldsub=-9.35488535307965e-7
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.824071664889999 lpclm=6.73927065840326e-7
+  pdiblc1=0.237773365950998 lpdiblc1=6.0036662202585e-7
+  pdiblc2=0.000570120761530006 lpdiblc2=2.83913172860183e-9
+  pdiblcb=-0.025
+  drout=0.690395324916501 ldrout=-5.14266121938182e-7
+  pscbe1=174537790.41 lpscbe1=201.385628767002
+  pscbe2=1.546132530315e-08 lpscbe2=-1.84156980549338e-15
+  pvag=0.0
+  delta=0.01
+  alpha0=3.742485758835e-05 lalpha0=-7.27499862759935e-11
+  alpha1=-9.71949999999999e-11 lalpha1=3.833273605e-16
+  beta0=71.40006536645 lbeta0=-0.000132962887065842
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=6.063342208e-08 lagidl=-1.17660033341312e-13
+  bgidl=2356411130.00001 lbgidl=-2581.32644560702
+  cgidl=743.183500000003 lcgidl=0.00180163859435001
+  egidl=1.263450842653 legidl=-6.87706687799169e-7
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.486300099999999 lkt1=-3.14328435609998e-7
+  kt2=-0.019032
+  at=659198.248 lat=-1.2137677542872
+  ute=-1.37210517 lute=-1.51030980036996e-7
+  ua1=-4.933329728e-10 lua1=2.03280032582592e-15 wua1=3.45126646034193e-31 pua1=1.50463276905253e-36
+  ub1=-1.242110355e-18 lub1=-4.56581219091547e-24
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.76 pmos
* DC IV MOS Parameters
+  lmin=1e-06 lmax=2e-06 wmin=7e-07 wmax=7.5e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.972874010000002+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-7.52287356099563e-9
+  k1=0.55984
+  k2=0.03253633478 lk2=3.33905495275805e-9
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=8629.50079999992 lvsat=0.05748209339488
+  ua=2.0923194407e-09 lua=1.26054003326808e-18
+  ub=-3.65505846000001e-19 lub=-3.09355239605989e-26
+  uc=-2.7970035e-12
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0169414093 lu0=-3.43116428270012e-10
+  a0=0.73934
+  keta=-0.0414997913 lketa=8.37974720806995e-9
+  a1=0.0
+  a2=0.5
+  ags=0.43242187
+  b0=4.415611461e-08 lb0=-4.4604952190379e-14
+  b1=9.56360298999998e-07 lb1=-1.3713831532261e-12 wb1=-8.07793566946316e-28
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.075734118+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.93596926797001+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-3.67395677006884e-07 wnfactor=3.3881317890172e-21
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.0825488271000001 leta0=-4.38326649996901e-8
+  etab=0.00409718673 letab=-7.96452128444701e-9
+  dsub=0.31595571
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=1.1707598
+  pdiblc1=0.54661982
+  pdiblc2=0.0020306546
+  pdiblcb=-0.025
+  drout=0.42584153
+  pscbe1=278136550.0
+  pscbe2=1.4513967e-8
+  pvag=0.0
+  delta=0.01
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=3.0
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=1.056e-10
+  bgidl=1028500000.0
+  cgidl=2308.019766 lcgidl=-0.0012402466231274
+  egidl=0.90967406
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.648
+  kt2=-0.019032
+  at=39330.72 lat=-0.00880726660799991
+  ute=-1.4498
+  ua1=5.524e-10
+  ub1=-3.5909e-18
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=2.81e-6
+  sbref=2.81e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.77 pmos
* DC IV MOS Parameters
+  lmin=8.0e-07 lmax=1e-06 wmin=7e-07 wmax=7.5e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.994695417999992+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=1.30743534501967e-8
+  k1=0.55984
+  k2=0.0280795226499997 lk2=7.5458399222648e-9
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=16508.0152999992 lvsat=0.0500455635583297
+  ua=2.067826692e-09 lua=2.43792455311992e-17
+  ub=-1.025276115e-18 lub=5.91821632948499e-25
+  uc=-2.7970035e-12
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0163138155 lu0=2.49269359549936e-10
+  a0=0.73934
+  keta=-0.032622
+  a1=0.0
+  a2=0.5
+  ags=0.43242187
+  b0=-1.462997805e-08 lb0=1.0883240671395e-14
+  b1=-2.343373335e-06 lb1=1.7432354239065e-12
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.075734118+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.63584464564998+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-8.41080459990356e-8
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.036111
+  etab=-0.0043407
+  dsub=0.31595571
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=1.1707598
+  pdiblc1=0.54661982
+  pdiblc2=0.0020306546
+  pdiblcb=-0.025
+  drout=0.42584153
+  pscbe1=278136550.0
+  pscbe2=1.4513967e-8
+  pvag=0.0
+  delta=0.01
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=3.0
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-3.94300800000001e-10 lagidl=4.7185636512e-16
+  bgidl=1028500000.0
+  cgidl=994.06
+  egidl=0.90967406
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.649859749999997 lkt1=1.75541802500059e-9
+  kt2=-0.019032
+  at=104390 lat=-0.070216721
+  ute=-1.33821499999999 lute=-1.05325081499995e-7
+  ua1=5.524e-10
+  ub1=-3.5909e-18
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=2.41e-6
+  sbref=2.41e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.78 pmos
* DC IV MOS Parameters
+  lmin=6e-07 lmax=8.0e-07 wmin=7e-07 wmax=7.5e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.826650064999988+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-1.11934584646502e-7
+  k1=0.530333425000002 lk1=2.19499411425018e-8
+  k2=0.0476809993440004 lk2=-7.03569859040166e-9
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=120138.23575 lvsat=-0.0270449574344251
+  ua=5.218192662745e-09 lua=-2.31917800010601e-15
+  ub=-4.95603783000001e-18 lub=3.515915272737e-24 wub=2.93873587705572e-39 pub=2.80259692864963e-45
+  uc=-2.66619636585002e-12 luc=-9.73074270941982e-20
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0188305644850001 lu0=-1.6229402103915e-9
+  a0=0.546337084999998 la0=1.43574868468504e-7
+  keta=0.0776265300000001 lketa=-8.20138814670004e-8
+  a1=0.0
+  a2=0.5
+  ags=-0.985510282385004 lags=1.0547997281592e-6
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={0.0101026353239995+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=-6.38539607977236e-8
+  nfactor={2.26896012949999+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-5.55082654435051e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=2.35975e-05 lcit=-1.011518025e-11
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.0775235459999999 leta0=-3.08067929693999e-8
+  etab=-0.01614523365 letab=8.78139258223501e-9
+  dsub=0.38515300677 ldsub=-5.14758690672026e-8
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=1.0386470339 lpclm=9.82786867017858e-8
+  pdiblc1=0.402732897065 lpdiblc1=1.07037481971348e-7
+  pdiblc2=-0.00480832577935002 lpdiblc2=5.08751750419848e-9
+  pdiblcb=-0.025
+  drout=-1.13320914871 ldrout=1.15977779989237e-06 pdrout=8.07793566946316e-28
+  pscbe1=-53271102.2749996 lpscbe1=246.534152527372
+  pscbe2=1.46067563400001e-08 lpscbe2=-6.9025990026001e-17
+  pvag=0.0
+  delta=0.01
+  alpha0=-9.31901922020003e-05 lalpha0=6.93242583690678e-11 walpha0=-7.57503684238477e-27 palpha0=2.73502740803562e-32
+  alpha1=3.71950000000001e-10 lalpha1=-2.02303605e-16
+  beta0=-123.4557519435 lbeta0=9.40704338707698e-05 wbeta0=9.48676900924816e-20
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-7.82447700000002e-08 lagidl=5.83848204030001e-14 wagidl=3.62876016401665e-29 pagidl=2.40741243048404e-35
+  bgidl=-908327900.0 lbgidl=1440.80627481
+  cgidl=1521.80617 lcgidl=-0.000392590375862999
+  egidl=0.791128117940005 legidl=8.81863262984351e-8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.767212390000001 lkt1=8.90540469210002e-8
+  kt2=-0.019032
+  at=10000.0
+  ute=-1.85672269999999 lute=2.80392796529993e-7
+  ua1=5.53487799999998e-10 lua1=-8.09214419998155e-19
+  ub1=-8.27197534999998e-18 lub1=3.482251952865e-24
+  uc1=-3.05199803999999e-10 luc1=1.458042541956e-16
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=2.02e-6
+  sbref=2.01e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.79 pmos
* DC IV MOS Parameters
+  lmin=5e-07 lmax=6e-07 wmin=7e-07 wmax=7.5e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.04745382+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=8.16057769799985e-9
+  k1=0.741369550000009 lk1=-9.28326072449988e-8
+  k2=-0.0251174394720004 lk2=3.25593722816208e-8
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=6327.81309999991 lvsat=0.0348565314449099
+  ua=-3.43364566709001e-09 lua=2.38655686749125e-15
+  ub=6.58897623000002e-18 lub=-2.763417874497e-24
+  uc=7.11466689520002e-12 luc=-5.41711895477929e-18
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.00986360823999988 lu0=3.25418729126401e-9
+  a0=1.37801371 la0=-3.08774047868998e-7
+  keta=-0.185699528000001 lketa=6.12091614792e-8
+  a1=0.0
+  a2=0.5
+  ags=0.798301705699998 lags=8.45843878397766e-8
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.142934161608+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=1.93827530535911e-8
+  nfactor={1.181815+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=3.6215581500003e-8
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-1.7195e-05 lcit=1.20718605e-11
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=-0.189143846 leta0=1.142336015394e-07 weta0=1.05879118406788e-22 peta0=-1.0097419586829e-28
+  etab=0.0194086397 letab=-1.055635913283e-8
+  dsub=0.38302338315 ldsub=-5.03175667802839e-8
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=2.01897928439999 lpclm=-4.34924024345167e-7
+  pdiblc1=2.45984227137001 lpdiblc1=-1.01182430671314e-6
+  pdiblc2=0.00827534028889998 lpdiblc2=-2.0286884703227e-9
+  pdiblcb=-0.025
+  drout=0.995253439089993 ldrout=2.10699838794419e-9
+  pscbe1=400000000.0
+  pscbe2=1.33187732819999e-08 lpscbe2=6.3150799522026e-16
+  pvag=0.0
+  delta=0.01
+  alpha0=0.000100102740071 lalpha0=-3.58077674942169e-11
+  alpha1=0.0
+  beta0=62.275976117 lbeta0=-6.94905302133625e-6
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=1.09001000000001e-08 lagidl=9.89892561000003e-15
+  bgidl=1547603499.99998 lbgidl=105.025186350002
+  cgidl=622.440000000002 lcgidl=9.65748840000002e-5
+  egidl=1.05976651579999 legidl=-5.79260982976206e-8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.403725000000001 lkt1=-1.08646744499999e-7
+  kt2=-0.019032
+  at=32195.0000000001 lat=-0.0120718605
+  ute=-1.21513240000002 lute=-6.85681676400044e-8
+  ua1=5.52e-10
+  ub1=1.7206632e-18 lub1=-1.95274415448001e-24
+  uc1=2.82799608000001e-10 luc1=-1.740086259912e-16
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=1.81e-6
+  sbref=1.81e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.80 pmos
* DC IV MOS Parameters
+  lmin=2.0e-05 lmax=1.0e-04 wmin=4.2e-07 wmax=7.0e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.9842405582+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} wvth0=-1.26811230782126e-8
+  k1=0.533428779142857 wk1=2.29718447009167e-8
+  k2=0.0330459994132571 wk2=-2.86940090944379e-9
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=362016.462771429 wvsat=-0.111015648733769
+  ua=3.57327410982e-09 wua=-6.57371311710562e-16
+  ub=-9.91202620628571e-19 wub=5.55115096895637e-25
+  uc=-2.19106346628286e-11 wuc=-6.5560611440841e-18
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0215120007877143 wu0=-1.35497753120905e-9
+  a0=0.843960620285714 wa0=1.99946820658811e-8
+  keta=-0.0118293050857143 wketa=2.52480734145966e-9
+  a1=0.0
+  a2=0.5
+  ags=0.144013050978 wags=-1.19854570004519e-8
+  b0=-8.98078809142857e-08 wb0=-3.08121880480365e-15
+  b1=1.33211450857143e-07 wb1=1.21442221467003e-13
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.0934891375457143+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} wvoff=-9.49924438140418e-9
+  nfactor={1.05990856971429+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} wnfactor=2.74144650601879e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=2.17162144007122e-05 wcit=-7.15973175541762e-12
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=2.07268965160714 wpclm=-6.58602390138518e-7
+  pdiblc1=0.39
+  pdiblc2=0.00129
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=226310255.298571 wpscbe1=-0.433820288335795
+  pscbe2=1.49877431602286e-08 wpscbe2=4.05819062096117e-18
+  pvag=0.0
+  delta=0.01
+  alpha0=4.14205208003143e-05 walpha0=-1.37141356453009e-11
+  alpha1=-1.18248571428571e-10 walpha1=7.22612290057143e-17
+  beta0=78.7028147359143 wbeta0=-2.50648991478023e-5
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.53957028571428e-08 wagidl=-1.50303356331886e-14
+  bgidl=2240640491.42857 wbgidl=-329.222159350034
+  cgidl=963.502857142857 wcgidl=0.000144522458011428
+  egidl=0.0119270576628572 wegidl=6.58242998916059e-7
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.578144128285714 wkt1=7.42122821888682e-9
+  kt2=-0.019032
+  at=711672.448 wat=-0.220136608043008
+  ute=-1.36972249142857 wute=-2.48578627779657e-8
+  ua1=-7.87272901942857e-10 wua1=4.94602098501672e-16
+  ub1=-1.51861164571429e-18 wub1=-5.38490678550583e-25
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.81 pmos
* DC IV MOS Parameters
+  lmin=8e-06 lmax=2.0e-05 wmin=4.2e-07 wmax=7.0e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.984107554749542+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-2.65260751560221e-09 wvth0=-1.11211803104473e-08 pvth0=-3.11113425660315e-14
+  k1=0.476280230711945 lk1=1.13976493505127e-06 wk1=5.23002994975072e-08 pk1=-5.84923769617722e-13
+  k2=0.0444539465967597 lk2=-2.27518957833057e-07 wk2=-9.18270646753405e-09 pk2=1.25911934719996e-13
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=548605.740288925 lvsat=-3.72131789188119 wvsat=-0.184507083065118 pvsat=1.46570581716099e-6
+  ua=4.39426557591542e-09 lua=-1.63737717006604e-14 wua=-1.06742994153536e-15 pua=8.17816830736285e-21
+  ub=-1.8694799005096e-18 lub=1.75162742422192e-23 wub=9.43777157546401e-25 pub=-7.75143727141275e-30
+  uc=4.06294387687678e-12 luc=-5.18014453038029e-16 wuc=-1.73839606629153e-17 puc=2.15950545213617e-22
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0239813531389688 lu0=-4.92485163581857e-08 wu0=-2.67231356051981e-09 pu0=2.62728180349709e-14
+  a0=0.765148919390129 la0=1.57181268149146e-06 wa0=5.14260219919094e-08 pa0=-6.26863500350709e-13
+  keta=-0.0118726904364418 lketa=8.65273096375103e-10 wketa=2.7471984462539e-09 pketa=-4.43534595490588e-15
+  a1=0.0
+  a2=0.5
+  ags=0.107001972769599 lags=7.38145242680524e-07 wags=-2.20718944119502e-09 pags=-1.95016790375063e-13
+  b0=-1.83110383651726e-07 lb0=1.86081578434523e-12 wb0=1.55649048212982e-14 pb0=-3.71876424986612e-19
+  b1=4.55272189174769e-07 lb1=-6.42314715893291e-12 wb1=5.89153526615499e-14 pb1=1.24702961876908e-18
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.0993412521506218+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=1.16713988468816e-07 wvoff=-6.47063056623251e-09 pvoff=-6.0402371068402e-14
+  nfactor={0.913198908253605+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=2.92596281720567e-06 wnfactor=3.59781251118689e-07 pnfactor=-1.70792779704721e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=3.08252198101732e-05 lcit=-1.81669092985749e-10 wcit=-1.07035062274509e-11 pcit=7.06766836927852e-17
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=3.38949574145214 lpclm=-2.62622489752596e-05 wpclm=-1.09459156446614e-06 ppclm=8.69532449387262e-12
+  pdiblc1=0.39
+  pdiblc2=0.00159345102002661 lpdiblc2=-6.05199679830869e-09 wpdiblc2=-1.05441755400639e-09 ppdiblc2=2.1029198255348e-14
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=227585626.888744 lpscbe1=-25.4358834572522 wpscbe1=-0.856090720355724 ppscbe1=8.42171926916224e-6
+  pscbe2=1.49814742278932e-08 lpscbe2=1.25026959604226e-16 wpscbe2=6.13380904148516e-18 ppscbe2=-4.1395926217136e-23
+  pvag=0.0
+  delta=0.01
+  alpha0=-2.39763167205118e-05 lalpha0=1.3042679878316e-09 walpha0=7.93849567049458e-12 palpha0=-4.31837913699092e-16
+  alpha1=-1.18248571428571e-10 walpha1=7.22612290057143e-17
+  beta0=76.7480651219377 lbeta0=3.8985330826187e-05 wbeta0=-2.44176893696131e-05 pbeta0=-1.29078870952272e-11
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=1.17967147624857e-07 lagidl=-1.24791863730282e-12 wagidl=-4.88984582819997e-14 pagidl=6.75462451295625e-19
+  bgidl=2544905524.93657 lbgidl=-6068.2314017802 wbgidl=-441.733210861339 pbgidl=0.00224390916023631
+  cgidl=741.083019596429 lcgidl=0.00443591899804222 wcgidl=0.000199534239150034 pcgidl=-1.09714946185024e-9
+  egidl=-0.610569110040606 legidl=1.24150013190611e-05 wegidl=8.64348990058005e-07 pegidl=-4.11055727673585e-12
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.584975399788359 lkt1=1.36242195721608e-07 wkt1=7.55038631373397e-09 pkt1=-2.57591612782215e-15
+  kt2=-0.019032
+  at=1082773.3570556 lat=-7.40119942011399 wat=-0.365865208095746 pat=2.90639662659179e-6
+  ute=-1.24634213390019 lute=-2.46068551251027e-06 wute=-4.13135607881226e-08 pute=3.28190795544766e-13
+  ua1=-1.32306837028818e-09 lua1=1.06858512411323e-14 wua1=8.22024566025625e-16 pua1=-6.53008095005097e-21
+  ub1=-4.87170139246762e-19 lub1=-2.05709662608377e-23 wub1=-8.94967020328747e-25 pub1=7.10952851278954e-30
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.82 pmos
* DC IV MOS Parameters
+  lmin=4e-06 lmax=8e-06 wmin=4.2e-07 wmax=7.0e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.997304754939704+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=1.02184631075026e-07 wvth0=-9.62130664034661e-09 pvth0=-4.30261890139464e-14
+  k1=0.69048720175015 lk1=-5.61873822179132e-07 wk1=-5.62215454546716e-08 pk1=2.77162914497891e-13
+  k2=-0.00305980628874036 lk2=1.49925543714067e-07 wk2=1.72205765299458e-08 pk2=-8.38331050836837e-14
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=-88726.7684408283 lvsat=1.3415878242171 wvsat=0.0428341564796681 pvsat=-3.40270255658836e-7
+  ua=1.729178104132e-09 lua=4.79741666643989e-15 wua=1.94610467560618e-16 pua=-1.84735449845473e-21
+  ub=1.39035178232345e-18 lub=-8.37950266303819e-24 wub=-4.56094256604487e-25 pub=3.36900125546048e-30
+  uc=-8.32112319812993e-11 luc=1.75282872561736e-16 wuc=1.57711373774383e-17 puc=-4.7430238109148e-23
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0170630596607568 lu0=5.70971520338282e-09 wu0=7.88726650315686e-10 pu0=-1.22133929588523e-15
+  a0=0.970392930397791 la0=-5.86252175523062e-08 wa0=-7.07707118098685e-09 pa0=-1.62120778494539e-13
+  keta=-0.0126972771811011 lketa=7.41570773727422e-09 wketa=2.46758614554406e-09 pketa=-2.21413379929702e-15
+  a1=0.0
+  a2=0.5
+  ags=0.263236975782276 lags=-5.02969997751882e-07 wags=-4.63255576838939e-08 pags=1.55455115108112e-13
+  b0=2.47361706307178e-07 lb0=-1.55881145107931e-12 wb0=-9.4012217117281e-14 pb0=4.98593273981268e-19
+  b1=-7.39430498613314e-07 lb1=3.06745152258685e-12 wb1=2.51860745808118e-13 pb1=-2.85709289847938e-19
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.0942818424831241+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=7.65225440111805e-08 wvoff=-7.37205553068603e-09 pvoff=-5.32415412932798e-14
+  nfactor={0.982552238947723+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=2.37502689350468e-06 wnfactor=3.33468055197501e-07 pnfactor=-1.49889839996889e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.11585905357149e-07 lcit=6.23169433907191e-11 wcit=-2.53365934201313e-14 pcit=-1.41496280629922e-17
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-0.463968355627997 lpclm=4.34928446553531e-06 wpclm=-2.14578108406042e-07 ppclm=1.70458560027682e-12
+  pdiblc1=0.39
+  pdiblc2=0.000379646939920181 lpdiblc2=3.59034143364881e-09 wpdiblc2=3.16325266201915e-09 ppdiblc2=-1.24755521737373e-14
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=222485819.425999 lpscbe1=15.0764770460487 wpscbe1=0.831965039904105 ppscbe1=-4.98802688476594e-6
+  pscbe2=1.50065627821497e-08 lpscbe2=-7.42740065541786e-17 wpscbe2=-2.17650189479598e-18 ppscbe2=2.4620352829619e-23
+  pvag=0.0
+  delta=0.01
+  alpha0=0.000263331131984429 lalpha0=-9.78073653935575e-10 walpha0=-9.43894789799746e-11 palpha0=3.8104528412677e-16
+  alpha1=-2.34838706642857e-10 lalpha1=9.26180375128763e-16 walpha1=1.43508994274623e-16 palpha1=-5.65985122519687e-22
+  beta0=124.165287064102 lbeta0=-0.000337692338560171 wbeta0=-5.12048444619281e-05 pbeta0=1.99886594242614e-10
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-6.97097288359285e-08 lagidl=2.42967701614019e-13 wagidl=4.83139823638406e-14 pagidl=-9.67834559508665e-20
+  bgidl=1723947084.01969 lbgidl=453.380357019396 wbgidl=-233.745165071998 pbgidl=0.000591672923290364
+  cgidl=1397.58209935357 lcgidl=-0.00077924404164055 wcgidl=0.00012198264513343 pcgidl=-4.81087354141735e-10
+  egidl=1.09728801061836 legidl=-1.15204486174164e-06 wegidl=5.17880042879673e-07 pegidl=-1.35824260724591e-12
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.569624120664286 lkt1=1.42931694878775e-08 wkt1=1.43508994274624e-08 pkt1=-5.65985122519689e-14
+  kt2=-0.019032
+  at=-200104.230448907 lat=2.78985184726307 wat=0.0938974298478952 pat=-7.45911792968695e-7
+  ute=-1.73706540076857 lute=1.43757104716545e-06 wute=2.27992848860506e-08 pute=-1.81115239206298e-13
+  ua1=2.2096e-11
+  ub1=-3.7441064775e-18 lub1=5.30181031661225e-24
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.83 pmos
* DC IV MOS Parameters
+  lmin=2e-06 lmax=4e-06 wmin=4.2e-07 wmax=7.0e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.03958725087928+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=2.68942566811102e-07 wvth0=4.36298544993564e-09 pvth0=-9.81788385888104e-14
+  k1=0.572793789436142 lk1=-9.77027733539172e-08 wk1=5.55645855622697e-09 pk1=3.35166444793081e-14
+  k2=0.0182154642762419 lk2=6.60180041328334e-08 wk2=2.68704174750615e-09 pk2=-2.651429725522e-14
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=565184.890205157 lvsat=-1.2373743663168 wvsat=-0.150740393328831 pvsat=4.23168411330903e-7
+  ua=3.61850171779593e-09 lua=-2.65388673348927e-15 wua=-4.44706853016011e-16 pua=6.74049082167442e-22
+  ub=-1.6440041341739e-19 lub=-2.24771547825592e-24 wub=2.27220405325205e-25 pub=6.74076560275973e-31
+  uc=-8.37276186182824e-11 luc=1.77319449819333e-16 wuc=1.34952546976371e-17 puc=-3.84543844082801e-23
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0229122862855888 lu0=-1.73590496822921e-08 wu0=-7.08093713506057e-10 pu0=4.68197053699136e-15
+  a0=1.32731514513517 la0=-1.46629074025506e-06 wa0=-1.93807588297675e-07 pa0=5.74325707961965e-13
+  keta=0.0472134033124747 lketa=-2.2886602506134e-07 wketa=-1.60394576588277e-08 pketa=7.07757962607647e-14
+  a1=0.0
+  a2=0.5
+  ags=-0.534745384067152 lags=2.64419263125828e-06 wags=2.1985005261376e-07 pags=-8.94314874344806e-13
+  b0=-4.23478259749314e-07 lb0=1.08691429105089e-12 wb0=1.31889025899135e-13 pb0=-3.92338638351175e-19
+  b1=-4.11894526961079e-07 lb1=1.7756824039876e-12 wb1=5.0270027670644e-13 pb1=-1.27499531575783e-18
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.153027683480443+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=3.08210266320505e-07 wvoff=7.10605398526281e-09 pvoff=-1.1034175741323e-13
+  nfactor={0.859430688314401+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=2.86060597704744e-06 wnfactor=2.55027370159483e-07 pnfactor=-1.18953618224745e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.59124285714286e-05 wcit=-3.61306145028571e-12
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.593645305699999 leta0=-2.02576572115023e-06 weta0=-3.02007496588047e-07 peta0=1.1910873657936e-12
+  etab=-1.352289899935 letab=5.05722313635364e-06 wetab=7.42025395686679e-07 petab=-2.92647395804869e-12
+  dsub=0.732887999474988 ldsub=-6.81852981129402e-07 wdsub=3.93001020858297e-08 pdsub=-1.54995672616304e-13
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.928664736892841 lpclm=-1.14312118805762e-06 wpclm=-6.39164079286478e-08 ppclm=1.11039091976402e-12
+  pdiblc1=0.280052772869484 lpdiblc1=4.33620869080041e-07 wpdiblc1=-2.58367764502582e-08 ppdiblc1=1.01897662642173e-13
+  pdiblc2=-0.000281126153971653 lpdiblc2=6.19636443864881e-09 wpdiblc2=5.20193585075399e-10 ppdiblc2=-2.05159148017887e-15
+  pdiblcb=-0.025
+  drout=0.557580954635464 ldrout=9.54047301319364e-09 wdrout=8.116233042126e-08 pdrout=-3.20096114948408e-13
+  pscbe1=192833565.579826 lpscbe1=132.022000989969 wpscbe1=-11.1804750231803 ppscbe1=4.23878354800329e-5
+  pscbe2=1.57099244156618e-08 lpscbe2=-2.84826195296262e-15 wpscbe2=-1.51917923259513e-16 ppscbe2=6.15185544549921e-22
+  pvag=0.0
+  delta=0.01
+  alpha0=3.68696372155151e-05 lalpha0=-8.49321647164565e-11 walpha0=3.39292948957914e-13 palpha0=7.44448051625315e-18
+  alpha1=-2.12126699e-10 lalpha1=8.366064881861e-16 walpha1=7.0234301532104e-17 palpha1=-2.76997061812465e-22
+  beta0=110.174986932431 lbeta0=-0.000282515993870875 wbeta0=-2.36951994692847e-05 pbeta0=9.13913053561281e-11
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=6.2638890748856e-08 lagidl=-2.79002019166413e-13 wagidl=-1.22553388166323e-15 pagidl=9.8595442169776e-20
+  bgidl=3247727147.06331 lbgidl=-5556.25583361834 wbgidl=-544.679652763323 pbgidl=0.00181796744929618
+  cgidl=147.837299180001 lcgidl=0.004149624475764 wcgidl=0.000363813681936298 pcgidl=-1.43484478018857e-9
+  egidl=1.35461152545574 legidl=-2.1669030719088e-06 wegidl=-5.57079286180244e-08 pegidl=9.03930993543863e-13
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.4173410806 lkt1=-5.86295912221661e-07 wkt1=-4.21405809192624e-08 pkt1=1.66198237087479e-13
+  kt2=-0.019032
+  at=1137984.62130581 lat=-2.48743677517237 wat=-0.29258443758169 pat=7.78334043986845e-7
+  ute=-1.18278564786086 lute=-7.48452870327278e-07 wute=-1.15692402701141e-07 pute=3.65082127468828e-13
+  ua1=-4.933329728e-10 lua1=2.03280032582592e-15 wua1=-6.16297582203915e-33 pua1=7.05296610493373e-38
+  ub1=-7.96979884773e-19 lub1=-6.32136225244376e-24 wub1=-2.72017449833839e-25 pub1=1.07280962039968e-30
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.84 pmos
* DC IV MOS Parameters
+  lmin=1e-06 lmax=2e-06 wmin=4.2e-07 wmax=7.0e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.795555927916648+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-2.05429921895948e-07 wvth0=-1.08358370688808e-07 pvth0=1.20940205609293e-13
+  k1=0.512470086124013 lk1=1.95604735145309e-08 wk1=2.89475648899601e-08 pk1=-1.19533271228358e-14
+  k2=0.0596916178446797 lk2=-1.46074907888527e-08 wk2=-1.65944848596935e-08 pk2=1.09670623165153e-14
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=-181973.558498617 lvsat=0.215026942118462 wvsat=0.116476767125148 pvsat=-9.6275026875586e-8
+  ua=2.14112513944004e-09 lua=2.17985597176734e-16 wua=-2.98249672772466e-17 pua=-1.32439815520142e-22
+  ub=-2.65901606382116e-18 lub=2.60156788456397e-24 wub=1.40155492006964e-24 pub=-1.60871230293573e-30
+  uc=1.55283901134655e-11 luc=-1.56243055543113e-17 wuc=-1.11985747356143e-17 puc=9.54795062701741e-24
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.00987557499279867 lu0=7.98301339976266e-09 wu0=4.3179030817935e-09 pu0=-5.08806463339144e-15
+  a0=0.297744294928933 la0=5.35092035460848e-07 wa0=2.69857368986109e-07 pa0=-3.26992602501982e-13
+  keta=-0.0839431700948643 lketa=2.60892379851867e-08 wketa=2.59369790080264e-08 pketa=-1.08221989759329e-14
+  a1=0.0
+  a2=0.5
+  ags=0.856897652364357 lags=-6.10222672609312e-08 wags=-2.59395452699729e-07 pags=3.7290463434086e-14
+  b0=-2.87939802866084e-07 lb0=8.2344108471558e-13 wb0=2.02942486785965e-13 pb0=-5.30459460969084e-19
+  b1=5.7425538298745e-06 lb1=-1.01879497568651e-11 wb1=-2.92482372194329e-12 pb1=5.38776858521737e-18
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={0.132897168013787+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=-2.47599052499129e-07 wvoff=-1.27493744357881e-07 pvoff=1.51306790586008e-13
+  nfactor={3.4027750176073+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-2.08340106466502e-06 wnfactor=-8.96359126380354e-07 pnfactor=1.04864402837634e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.59124285714286e-05 wcit=-3.61306145028571e-12
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=-0.625343356826294 leta0=3.43826339934633e-07 weta0=4.32590082028623e-07 peta0=-2.36896867279345e-13
+  etab=2.43658660451876 letab=-2.30797390065401e-06 wetab=-1.48648455325304e-06 petab=1.40552653169522e-12
+  dsub=0.391402908723753 ldsub=-1.80401132180775e-08 wdsub=-4.61054813512905e-08 pdsub=1.10242410271142e-14
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-0.663901306511656 lpclm=1.95266794371638e-06 wpclm=1.12115406354485e-06 ppclm=-1.19326756973331e-12
+  pdiblc1=0.321386109861017 lpdiblc1=3.53272995302199e-07 wpdiblc1=1.37639419331092e-07 ppdiblc1=-2.15883714337193e-13
+  pdiblc2=0.00277541341441945 lpdiblc2=2.54757171653334e-10 wpdiblc2=-4.5511913245647e-10 ppdiblc2=-1.55681088568666e-16
+  pdiblcb=-0.025
+  drout=1.19382536675318 ldrout=-1.22725503970243e-06 wdrout=-4.69311850704522e-07 pdrout=7.49970645741999e-13
+  pscbe1=278763719.572086 lpscbe1=-35.0176253555846 wpscbe1=-0.383260816823736 ppscbe1=2.13991307842963e-5
+  pscbe2=1.44032515084451e-08 lpscbe2=-3.08220488624123e-16 wpscbe2=6.76577940272174e-17 ppscbe2=1.88352307716245e-22
+  pvag=0.0
+  delta=0.01
+  alpha0=-1.50395478404369e-06 lalpha0=-1.03377392285142e-11 walpha0=9.19121862309966e-13 palpha0=6.3173510915881e-18
+  alpha1=2.18248571428571e-10 walpha1=-7.22612290057143e-17
+  beta0=-29.6460280657749 lbeta0=-1.0717922815862e-05 wbeta0=1.99498571668828e-05 pbeta0=6.54967976108199e-12
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-1.01648407250857e-07 lagidl=4.03560594152292e-14 wagidl=6.21814668149698e-14 pagidl=-2.46614264844089e-20
+  bgidl=630425122.659754 lbgidl=-468.482428380266 wbgidl=243.261965243115 pbgidl=0.000286287738053467
+  cgidl=3505.34208833834 lcgidl=-0.0023770290838809 wcgidl=-0.000731678881891672 pcgidl=6.94683214636624e-10
+  egidl=-0.555217860916413 legidl=1.54561427226003e-06 wegidl=8.95189593304336e-07 pegidl=-9.44518699321014e-13
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.776988852674286 lkt1=1.12823391913544e-07 wkt1=7.88245719138454e-08 pkt1=-6.89459235047991e-14
+  kt2=-0.019032
+  at=-325948.435130286 lat=0.358302693233762 wat=0.223220630583497 pat=-2.24339428019462e-7
+  ute=-1.679203671204 lute=2.16534125249455e-07 wute=1.40187665858079e-07 pute=-1.32323137803441e-13
+  ua1=5.524e-10
+  ub1=-3.70543789578257e-18 lub1=-6.67610724842258e-25 wub1=6.99936499611455e-26 pub1=4.07974243508206e-31
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=2.81e-6
+  sbref=2.81e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.85 pmos
* DC IV MOS Parameters
+  lmin=8.0e-07 lmax=1e-06 wmin=4.2e-07 wmax=7.0e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.46431627084779+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=4.25812965796756e-07 wvth0=2.86983424691873e-07 pvth0=-2.52222915050531e-13
+  k1=0.283761272748497 lk1=2.35438722459681e-07 wk1=1.68710605908484e-07 pk1=-1.43875661540221e-13
+  k2=0.0681020858048794 lk2=-2.25461314964853e-08 wk2=-2.44576282536942e-08 pk2=1.83890833661126e-14
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=-84957.9086913415 lvsat=0.123453870265374 wvsat=0.0620054202874128 pvsat=-4.48595225954479e-8
+  ua=1.52232983088148e-09 lua=8.02066488925167e-16 wua=3.33350949842084e-16 pua=-4.7524156368908e-22
+  ub=2.72327613478046e-18 lub=-2.4787777216961e-24 wub=-2.29072528563184e-24 pub=1.87643098322589e-30
+  uc=-1.28600421124015e-12 luc=2.46801248778366e-19 wuc=-9.2336562136399e-19 puc=-1.50819255923465e-25
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0276685615227823 lu0=-8.81178658588894e-09 wu0=-6.93883987553819e-09 pu0=5.53717504403394e-15
+  a0=1.44479090552983 la0=-5.47605260285341e-07 wa0=-4.31098226565658e-07 pa0=3.34639384139331e-13
+  keta=-0.131209373527985 lketa=7.07038074057092e-08 wketa=6.02463496134575e-08 pketa=-4.32068138903993e-14
+  a1=0.0
+  a2=0.5
+  ags=2.01421311411026 lags=-1.15341233160289e-06 wags=-9.66626302110806e-07 pags=7.04845662193201e-13
+  b0=2.75827352395142e-06 lb0=-2.05187967446746e-12 wb0=-1.69451023845906e-12 pb0=1.26054616638969e-18
+  b1=-2.38377659842327e-05 lb1=1.77329141156707e-11 wb1=1.31351373703755e-11 pb1=-9.77122868982235e-18
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.480134223122378+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=3.31041277594298e-07 wvoff=2.47127286639865e-07 pvoff=-2.02298000572765e-13
+  nfactor={-1.54133853300296+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=2.583347715756e-06 wnfactor=1.94156393174211e-06 pnfactor=-1.63007154618545e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.59124285714286e-05 wcit=-3.61306145028572e-12
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.629828705144 leta0=-8.40930569359127e-07 weta0=-3.62818514742678e-07 peta0=5.13889307213085e-13
+  etab=-0.00518977054644128 letab=-3.18118022997047e-09 wetab=5.18863614648084e-10 petab=1.94400651381403e-15
+  dsub=1.25582656478186 ldsub=-8.33969602171324e-07 wdsub=-5.74351319873775e-07 pdsub=5.09635488008487e-13
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=1.50138756485271 lpclm=-9.11482219644497e-08 wpclm=-2.02045304590434e-07 ppclm=5.57003138495864e-14
+  pdiblc1=0.612442519987914 lpdiblc1=7.85448497834213e-08 wpdiblc1=-4.02239886718145e-08 ppdiblc1=-4.79984435232498e-14
+  pdiblc2=0.0264402026372479 lpdiblc2=-2.20824373757745e-08 wpdiblc2=-1.49165771673701e-08 ppdiblc2=1.34944891505863e-14
+  pdiblcb=-0.025
+  drout=-1.71215985295285 ldrout=1.51570440917808e-06 wdrout=1.30652409311695e-06 pdrout=-9.2624090163109e-13
+  pscbe1=241367569.395887 lpscbe1=0.280600795729697 wpscbe1=22.4693769712505 ppscbe1=-1.71474023867124e-7
+  pscbe2=1.21282629341076e-08 lpscbe2=1.83914122669303e-15 wpscbe2=1.45789421185056e-15 ppscbe2=-1.12389184706721e-21
+  pvag=0.0
+  delta=0.01
+  alpha0=-5.87869826958651e-05 lalpha0=4.37317108174541e-11 walpha0=3.59245510871124e-11 palpha0=-2.67242735537029e-17
+  alpha1=6.58074132857143e-10 lalpha1=-4.15151347432429e-16 walpha1=-3.41036870292469e-16 palpha1=2.53697327810567e-22
+  beta0=-204.662543535735 lbeta0=0.000154480166136233 wbeta0=0.000126901749704513 pbeta0=-9.44022116051875e-11
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=2.72147200889687e-06 lagidl=-2.62438730138661e-12 wagidl=-1.66332161439052e-12 pagidl=1.60404093186545e-18
+  bgidl=-702319682.45652 lbgidl=789.495393168986 wbgidl=1057.69698467045 pbgidl=-0.000482457476783995
+  cgidl=21870.8333426086 lcgidl=-0.0197122162787866 wcgidl=-0.0127577126825747 pcgidl=1.20460565191014e-8
+  egidl=6.51972018754148 legidl=-5.13241975167938e-06 wegidl=-3.42827674835609e-06 pegidl=3.13640118057226e-12
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.5625580122 lkt1=-8.95778784101337e-08 wkt1=-5.33497427626284e-08 pkt1=5.58134121183247e-14
+  kt2=-0.019032
+  at=216004.826571429 lat=-0.153246990486486 wat=-0.0682073740584937 pat=5.07394655621135e-8
+  ute=-1.338215 lute=-1.05325081499998e-7
+  ua1=5.524e-10
+  ub1=-4.41272757142857e-18 wub1=5.02215541589713e-25
+  uc1=-1.092e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=2.41e-6
+  sbref=2.41e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.86 pmos
* DC IV MOS Parameters
+  lmin=6e-07 lmax=8.0e-07 wmin=4.2e-07 wmax=7.0e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.558064692647251+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-2.48347583226624e-07 wvth0=-1.64131446703275e-07 pvth0=8.33614377803191e-14
+  k1=0.564196931124118 lk1=2.68226361940559e-08 wk1=-2.06938531384244e-08 pk1=-2.97768445522544e-15
+  k2=0.0432275006139837 lk2=-4.04192757297796e-09 wk2=2.72151525991801e-09 pk2=-1.82948149366351e-15
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=178069.579908598 lvsat=-0.0722122785041206 wvsat=-0.0354016126899425 pvsat=2.76015692364067e-8
+  ua=7.76241359106236e-09 lua=-3.8399318202734e-15 wua=-1.55476323241103e-15 pua=9.29326576489011e-22
+  ub=-9.37541582062067e-18 lub=6.5214392239268e-24 wub=2.70066421255633e-24 pub=-1.83666366447628e-30
+  uc=-1.65088913334329e-12 luc=5.18239142330895e-19 wuc=-6.20450188555919e-19 puc=-3.76158046389388e-25
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.0155163722732274 lu0=2.2822699685499e-10 wu0=2.0252896038454e-09 pu0=-1.13124087567951e-15
+  a0=-0.136546606731021 la0=6.28751715085507e-07 wa0=4.17307492482059e-07 pa0=-2.96489630260267e-13
+  keta=0.238488722765272 lketa=-2.04314606426845e-07 wketa=-9.83022425500867e-08 pketa=7.47374838200612e-14
+  a1=0.0
+  a2=0.5
+  ags=-2.54578392195299 lags=2.23876946352456e-06 wags=9.53476980045442e-07 pags=-7.23519169402832e-13
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={0.148074940307873+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=-1.36283519081466e-07 wvoff=-8.43143236864248e-08 pvoff=4.42614133489617e-14
+  nfactor={4.18612445575105+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.67731200157812e-06 wnfactor=-1.17157145111472e-06 pnfactor=6.85789865121739e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=6.16676275714286e-05 lcit=-3.40372925361e-11 wcit=-2.32645026783897e-11 pcit=1.46187071295866e-17
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=-1.68220605289058 leta0=8.78992087142794e-07 weta0=1.07536371896364e-06 peta0=-5.55974456441041e-13
+  etab=-0.150642763778943 letab=1.05021301435688e-07 wetab=8.21909026716768e-08 petab=-5.88118233407096e-14
+  dsub=-0.276965855507108 ldsub=3.06274679281639e-07 wdsub=4.04618188262091e-07 pdsub=-2.18619929093784e-13
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=1.4281061536073 lpclm=-3.66341801389834e-08 wpclm=-2.37996910216652e-07 ppclm=8.24447132749296e-14
+  pdiblc1=0.251125162132853 lpdiblc1=3.47328832291802e-07 wpdiblc1=9.26468803860956e-08 ppdiblc1=-1.46841083015429e-13
+  pdiblc2=-0.0286274445435638 lpdiblc2=1.88823853620314e-08 wpdiblc2=1.4555768200336e-08 ppdiblc2=-8.42998856845028e-15
+  pdiblcb=-0.025
+  drout=-2.4111417497724 ldrout=2.03567704222215e-06 wdrout=7.80939500778828e-07 pdrout=-5.3525852339076e-13
+  pscbe1=-236837638.804957 lpscbe1=356.017455176338 wpscbe1=112.176776207311 ppscbe1=-6.69048083155723e-5
+  pscbe2=1.27579085301273e-08 lpscbe2=1.370747867814e-15 wpscbe2=1.12982350122195e-15 ppscbe2=-8.79840045430584e-22
+  pvag=0.0
+  delta=0.01
+  alpha0=-0.000139558185443906 lalpha0=1.03817408541722e-10 walpha0=2.83352951981558e-11 palpha0=-2.10786260979081e-17
+  alpha1=3.7195e-10 lalpha1=-2.02303605e-16
+  beta0=-137.638708925486 lbeta0=0.000104621135569669 wbeta0=8.66714827986379e-06 pbeta0=-6.44749160539066e-12
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-2.91487613193114e-06 lagidl=1.56849208057535e-12 wagidl=1.73345407875067e-12 pagidl=-9.22820506262281e-19
+  bgidl=-3912089969.86831 lbgidl=3177.24350997462 wbgidl=1835.58698584824 pbgidl=-0.00106112984866016
+  cgidl=-15824.4005729203 lcgidl=0.00832926823097534 wcgidl=0.0106001975557716 pcgidl=-5.32989290720448e-9
+  egidl=-2.76384024294766 legidl=1.77362085256149e-06 wegidl=2.172426945465e-06 pegidl=-1.02996229726125e-12
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.899160058428571 lkt1=1.60820383779299e-07 wkt1=8.06326923860261e-08 pkt1=-4.38561213887596e-14
+  kt2=-0.019032
+  at=10000.0
+  ute=-1.53514571 lute=4.11716736690008e-08 wute=-1.9651441228104e-07 pute=1.46187071295865e-13
+  ua1=5.534878e-10 lua1=-8.09214420000127e-19
+  ub1=-1.13287630019286e-17 lub1=5.14483875674895e-24 wub1=1.86799070694294e-24 pub1=-1.01600014550627e-30
+  uc1=-5.369667722328e-10 luc1=3.1821570186398e-16 wuc1=1.41631867219191e-16 puc1=-1.05359946024356e-22
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=2.02e-6
+  sbref=2.01e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.87 pmos
* DC IV MOS Parameters
+  lmin=5e-07 lmax=6e-07 wmin=4.2e-07 wmax=7.0e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.175e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=2.805e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=4.4452e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.7338e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.577
+  rnoib=0.37
+  tnoia=1.5
+  tnoib=3.5
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.2455e-08+sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre*(1.2455e-08*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.920292953769325+sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-5.1331632002327e-08 wvth0=-7.77074967101001e-08 pvth0=3.63554513790317e-14
+  k1=0.828146444578352 lk1=-1.16739504173702e-07 wk1=-5.30290131692519e-08 pk1=1.4609409085542e-14
+  k2=-0.0494505190039934 lk2=4.63656472972399e-08 wk2=1.4869847569683e-08 pk2=-8.43695943694473e-15
+  k3=-2.2405
+  dvt0=4.657
+  dvt1=0.34864
+  dvt2=-0.030206
+  dvt0w=-2.2
+  dvt1w=1016300.0
+  dvt2w=0.0
+  w0=0.0
+  k3b=-0.172
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=-52527.7740062673 lvsat=0.0532096222901746 wvsat=0.0359664138582915 pvsat=-1.12155004031778e-8
+  ua=-1.51573773101998e-09 lua=1.20645468380719e-15 wua=-1.17202586810064e-15 pua=7.21155724040593e-22
+  ub=1.04192549331706e-18 lub=8.55447283276071e-25 wub=3.389780516984e-24 pub=-2.21147402245449e-30
+  uc=8.51631544345192e-12 luc=-5.01170342698803e-18 wuc=-8.56541821242558e-19 puc=-2.47747807371126e-25
+  rdsw=788.47
+  prwb=0.053538
+  prwg=0.0
+  wr=1.0
+  u0=0.00431292418352153 lu0=6.32178241284603e-09 wu0=3.39200082417777e-09 pu0=-1.87459510841829e-15
+  a0=-0.943454382667118 la0=1.06762885441715e-06 wa0=1.41863986555651e-06 pa0=-8.41114307975458e-13
+  keta=-0.328539821302111 lketa=1.04092218691405e-07 wketa=8.72891318757471e-08 pketa=-2.62056647301498e-14
+  a1=0.0
+  a2=0.5
+  ags=-0.912758372614142 lags=1.35056686723916e-06 wags=1.04562196961746e-06 pags=-7.73636829231052e-13
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.0235597028644077+sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))} lvoff=-4.29314366600625e-08 wvoff=-7.29492542403743e-08 pvoff=3.80799520772549e-14
+  nfactor={2.28808070781284+sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-6.44966007074519e-07 wnfactor=-6.76034548981595e-07 pnfactor=4.16267344051534e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-4.9352699e-05 lcit=2.63466630861e-11 wcit=1.9651441228104e-11 pcit=-8.72327476115537e-18
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=-0.997872740200232 leta0=5.06783198370516e-07 weta0=4.94210992330185e-07 peta0=-2.39885488425108e-13
+  etab=0.161195539690774 letab=-6.45875518214914e-08 wetab=-8.6645407436762e-08 petab=3.30182457272702e-14
+  dsub=0.413067179091799 ldsub=-6.90342882367067e-08 wdsub=-1.83596435248499e-08 pdsub=1.14377136151336e-14
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=3.06631863462312 lpclm=-9.27657948563489e-07 wpclm=-6.40024887563947e-07 ppclm=3.01107730154123e-13
+  pdiblc1=5.13040353250036 lpdiblc1=-2.30651067335109e-06 wpdiblc1=-1.63196930443172e-06 ppdiblc1=7.91177659906981e-13
+  pdiblc2=0.0338523313189721 lpdiblc2=-1.51003647296019e-08 wpdiblc2=-1.56299969105129e-08 ppdiblc2=7.98804907534046e-15
+  pdiblcb=-0.025
+  drout=1.89321025064145 ldrout=-3.05460010802943e-07 wdrout=-5.48737815711846e-07 pdrout=1.87952969048518e-13
+  pscbe1=298531226.702907 lpscbe1=64.830329226611 wpscbe1=62.0071614867607 ppscbe1=-3.96175548690651e-5
+  pscbe2=1.74445723072803e-08 lpscbe2=-1.17832856057953e-15 wpscbe2=-2.5212592811527e-15 ppscbe2=1.10598387990299e-21
+  pvag=0.0
+  delta=0.01
+  alpha0=0.000148449607267885 lalpha0=-5.28300299142215e-11 walpha0=-2.95445771565477e-11 palpha0=1.04022364758151e-17
+  alpha1=0.0
+  beta0=73.8823375132637 lbeta0=-1.04251615883669e-05 wbeta0=-7.09260102381109e-06 pbeta0=2.12423604087809e-12
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-2.73213070153714e-07 lagidl=1.31691541274605e-13 wagidl=1.73620421828254e-13 pagidl=-7.44269802621776e-20
+  bgidl=1980321031.12957 lbgidl=-27.6388334681269 wbgidl=-264.431952403152 pbgidl=8.10704518547783e-5
+  cgidl=-6883.18675323571 lcgidl=0.0034661420344489 wcgidl=0.00458665848639533 pcgidl=-2.05912900737072e-9
+  egidl=-0.248833943597596 legidl=4.05708926344994e-07 wegidl=7.99680506336034e-07 pegidl=-2.83325509019003e-13
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.175e-8
* Temperature Effects Parameters
+  kt1=-0.408974054085715 lkt1=-1.0579178398278e-07 wkt1=3.20767595556394e-09 pkt1=-1.74465495223118e-15
+  kt2=-0.019032
+  at=100432.703114286 lat=-0.04918634722386 wat=-0.0416997874223275 pat=2.26805143790039e-8
+  ute=-1.82049319058286 lute=1.96372168358016e-07 wute=3.69933557682022e-07 pute=-1.61903979567043e-13
+  ua1=5.52e-10
+  ub1=5.88967139119998e-19 lub1=-1.33721466696737e-24 wub1=6.91574936019525e-25 pub1=-3.7614760770102e-31
+  uc1=1.1017155022848e-09 luc1=-5.73063587246143e-16 wuc1=-5.00436227333864e-16 puc1=2.4386089060305e-22
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+40
+  noib=8.5300000000000003e+24
+  noic=84000000.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=4.02e-12
+  xtis=10.0
+  bvs=12.69
+  xjbvs=1.0
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.00096
+  tcjsw=3.0e-5
+  tcjswg=0.0
+  cgdo=2.5544132e-10
+  cgso=2.5544132e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=1.292646e-11
+  cgdl=1.292646e-11
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=2.7658e-8
+  dwc=3.2175e-8
+  vfbcv=-0.1446893
+  acde=0.401
+  moin=15.773
+  noff=4.0
+  voffcv=0.0
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000835724019
+  mjs=0.33956
+  pbs=0.6587
+  cjsws=1.059825712e-10
+  mjsws=0.24676
+  pbsws=1.0
+  cjswgs=1.567456e-10
+  mjswgs=0.81
+  pbswgs=3.0
* Stress Parameters
+  saref=1.81e-6
+  sbref=1.81e-6
+  wlod={0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.ends sky130_fd_pr__pfet_g5v0d10v5
