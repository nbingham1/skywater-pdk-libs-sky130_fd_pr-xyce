* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* statistics {
*   mismatch {
*   }
* }
* 4-terminal Vertical Parallel Plate Capacitor /w LI-M4 fingers and M5 Shield
* 4-terminal Vertical Parallel Plate Capacitor /w M1-M4 fingers and LI/M5 Shield
* Layout: sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3m4_shieldl1m5
.subckt sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3m4_shieldl1m5 c0 c1 b m5
.param mult=1.0
+  ctot_a={116.75e-15*sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3m4_shieldl1m5__cor+1.4*0.00244/sqrt(mult/0.27882)*116.75e-15*sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3m4_shieldl1m5__cor*sky130_fd_pr__model__cap_vpp_only_p__slope}
+  cm5_c0={5.41e-15*c0m5m4_vpp}
+  cm5_c1={3.88e-15*c1m5m4_vpp}
+  cli2s={(7.59-0.58)*1e-15*cli2s_vpp}
+  rat_m4=0.1376
+  rat_m3=0.1376
+  rat_m2=0.3485
+  rat_m1=0.3442
+  rat_m12li=0.0321
+  cap_m4={rat_m4*ctot_a}
+  cap_m3={rat_m3*ctot_a}
+  cap_m2={rat_m2*ctot_a}
+  cap_m1={rat_m1*ctot_a}
+  cap_m12li={rat_m12li*ctot_a}
+  lm1=5.215
+  lm2=5.095
+  lm3=5.050
+  lm4=4.910
+  wm1=0.140
+  wm2=0.140
+  wm3=0.300
+  wm4=0.300
+  nfm1=72.0
+  nfm2=72.0
+  nfm3=34.0
+  nfm4=34.0
+  nvia3_c0=103.0
+  nvia3_c1=49.0
+  nvia2_c0=104.0
+  nvia2_c1=49.0
+  nvia_c0=124.0
+  nvia_c1=62.0
+  nmcon=116.0
ccmvpp11p5x11p7_lim5shield m5 a0 c={cm5_c0}
cm5_1 m5 a1 c={cm5_c1}
rsm4 a0 a2 r={rm4*lm4/wm4*(1/3)*(1/nfm4)}
cm4 a2 a1 c={cap_m4}
rvia3_0 a0 b0 r={rcvia3/nvia3_c0}
rvia3_1 a1 b1 r={rcvia3/nvia3_c1}
rsm3 b0 b2 r={rm3*lm3/wm3*(1/3)*(1/nfm3)}
cm3 b2 b1 c={cap_m3}
rvia2_0 b0 c0 r={rcvia2/nvia2_c0}
rvia2_1 b1 c1 r={rcvia2/nvia2_c1}
rsm2 c0 c2 r={rm2*lm2/wm2*(1/3)*(1/nfm2)}
cm2 c2 c1 c={cap_m2}
rvia_0 c0 d0 r={rcvia/nvia_c0}
rvia_1 c1 d1 r={rcvia/nvia_c1}
rsm1 d0 d2 r={rm1*lm1/wm1*(1/3)*(1/nfm1)}
cm1 d2 d1 c={cap_m1}
rmcon d0 e0 r={rcl1/nmcon}
rliw e0 f0 r={rl1}
cli2b f0 b c={cli2s}
cm12li d1 f0 c={cap_m12li}
.ends sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3m4_shieldl1m5
