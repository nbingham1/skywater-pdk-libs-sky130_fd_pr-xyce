* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 11
.param
+  sky130_fd_pr__esd_nfet_g5v0d10v5__toxe_mult=0.94
+  sky130_fd_pr__esd_nfet_g5v0d10v5__rshn_mult=1.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__overlap_mult=0.76246
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ajunction_mult=8.1753e-1
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pjunction_mult=7.7786e-1
+  sky130_fd_pr__esd_nfet_g5v0d10v5__lint_diff=1.7325e-8
+  sky130_fd_pr__esd_nfet_g5v0d10v5__wint_diff=-3.2175e-8
+  sky130_fd_pr__esd_nfet_g5v0d10v5__dlc_diff=1.7325e-8
+  sky130_fd_pr__esd_nfet_g5v0d10v5__dwc_diff=-3.2175e-8
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 000, W = 17.5, L = 0.55
* -----------------------------------
+  sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_0=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_0=0.14328
+  sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_0=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_0=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_0=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_0=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_0=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_0=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_0=-0.00045472
+  sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_0=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_0=-0.0011699
+  sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_0=-0.0040664
+  sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_0=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_0=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_0=-7090.1
+  sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_0=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_0=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_0=-8.363e-19
+  sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_0=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_0=-2.0608e-12
+  sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_0=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_0=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_0=0.0
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 001, W = 19.5, L = 0.55
* -----------------------------------
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_1=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_1=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_1=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_1=0.15647
+  sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_1=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_1=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_1=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_1=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_1=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_1=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_1=0.00040364
+  sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_1=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_1=0.00057999
+  sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_1=-0.0025892
+  sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_1=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_1=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_1=-6925.9
+  sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_1=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_1=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_1=-7.4921e-19
+  sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_1=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_1=-1.8631e-11
+  sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_1=0.0
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 002, W = 21.5, L = 0.55
* -----------------------------------
+  sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_2=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_2=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_2=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_2=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_2=0.1669
+  sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_2=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_2=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_2=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_2=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_2=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_2=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_2=2.8343e-5
+  sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_2=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_2=-0.0010571
+  sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_2=-0.0034839
+  sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_2=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_2=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_2=-5424.6
+  sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_2=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_2=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_2=-7.5872e-19
+  sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_2=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_2=1.2923e-12
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 003, W = 23.5, L = 0.55
* -----------------------------------
+  sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_3=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_3=-1.6825e-12
+  sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_3=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_3=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_3=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_3=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_3=0.15401
+  sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_3=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_3=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_3=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_3=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_3=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_3=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_3=0.0001604
+  sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_3=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_3=-0.0013049
+  sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_3=-0.0016799
+  sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_3=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_3=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_3=-5330.1
+  sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_3=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_3=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_3=-7.6166e-19
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 004, W = 26.5, L = 0.55
* -----------------------------------
+  sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_4=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_4=-8.2209e-19
+  sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_4=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_4=-5.2787e-12
+  sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_4=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_4=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_4=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_4=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_4=0.14553
+  sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_4=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_4=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_4=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_4=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_4=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_4=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_4=-0.0026632
+  sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_4=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_4=-0.00096576
+  sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_4=-0.0043485
+  sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_4=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_4=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_4=-6212.8
+  sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_4=0.0
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 005, W = 30.25, L = 1.0
* -----------------------------------
+  sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_5=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_5=-1.0249e-18
+  sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_5=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_5=1.3027e-10
+  sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_5=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_5=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_5=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_5=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_5=0.17146
+  sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_5=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_5=0.24441
+  sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_5=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_5=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_5=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_5=-0.4
+  sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_5=0.054151
+  sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_5=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_5=-0.0059635
+  sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_5=-3.7876e-5
+  sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_5=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_5=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_5=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_5=0.0
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 006, W = 30.25, L = 0.55
* ------------------------------------
+  sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_6=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_6=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_6=-5.3272e-19
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_6=-1.7366e-12
+  sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_6=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_6=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_6=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_6=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_6=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_6=0.14152
+  sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_6=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_6=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_6=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_6=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_6=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_6=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_6=-0.0011048
+  sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_6=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_6=-0.00069586
+  sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_6=-0.0038289
+  sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_6=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_6=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_6=-4075.0
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 007, W = 40.31, L = 0.55
* ------------------------------------
+  sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_7=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_7=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_7=-2741.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_7=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_7=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_7=-2.1212e-19
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_7=2.6239e-12
+  sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_7=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_7=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_7=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_7=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_7=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_7=0.12367
+  sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_7=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_7=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_7=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_7=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_7=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_7=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_7=-0.0014188
+  sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_7=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_7=-0.00098518
+  sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_7=-0.0023054
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 008, W = 50.99, L = 1.0
* -----------------------------------
+  sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_8=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_8=-0.0085839
+  sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_8=-0.00047254
+  sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_8=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_8=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_8=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_8=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_8=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_8=-1.1983e-18
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_8=1.2035e-10
+  sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_8=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_8=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_8=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_8=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_8=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_8=0.17047
+  sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_8=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_8=0.16645
+  sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_8=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_8=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_8=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_8=-0.39993
+  sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_8=0.015735
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 009, W = 50.99, L = 0.55
* ------------------------------------
+  sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_9=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_9=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_9=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_9=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_9=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_9=-0.0059114
+  sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_9=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_9=0.0013661
+  sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_9=-0.010512
+  sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_9=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_9=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_9=-5727.6
+  sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_9=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_9=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_9=7.8668e-20
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_9=-1.2856e-11
+  sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_9=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_9=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_9=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_9=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_9=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_9=0.12716
+  sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_9=0.0
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 010, W = 5.4, L = 0.6
* ---------------------------------
+  sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_10=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_10=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_10=6.7679e-12
+  sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_10=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_10=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_10=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_10=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_10=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_10=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_10=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_10=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_10=-7615.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_10=-5.6629e-19
+  sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_10=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_10=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_10=-0.0031534
+  sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_10=0.28192
+  sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_10=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_10=-0.00288
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_10=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_10=-0.0017519
+  sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_10=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_10=0.0
.include "sky130_fd_pr__esd_nfet_g5v0d10v5.pm3.spice"
