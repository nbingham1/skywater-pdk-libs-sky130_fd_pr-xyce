* Transistor Vth and I-V characteristic
.options parser scale=1E-6

* Include SkyWater sky130 device models
.include "../sky130_fd_pr__rf_nfet_01v8_lvt_aM02W5p00L0p25.spice"
.lib "../../../models/sky130.lib.spice" tt

* Gate bias
Rg 1 2 680
X1 3 2 0 0 sky130_fd_pr__rf_nfet_01v8_lvt_aM02W5p00L0p25
Rd 3 4 100

* DC source for current measure
Vid 5 4 DC 0V
Vgb 1 0 DC 0V
Vdd 5 0 DC 3.3V

.control
* Sweep Vds from 0 to 1.8V
dc Vdd 0 1.8 0.01 Vgb 0 1.2 0.01
wrdata sky130_fd_pr__rf_nfet_01v8_lvt_aM02W5p00L0p25__iv.data Vid#branch V ( 1 ) V ( 3 )

* Sweep Vgs from 0 to 1.2V
dc Vgb 0 1.2 0.01
+ # Find threshold
let ih=Vid#branch[98]
let il=Vid#branch[85]
let vh=V(2)[98]
let vl=V(2)[85]
let vth=((vl - vh ) / ( ih - il ) ) * ih vh
echo threshold voltage
print vth
quit
.endc
.end
