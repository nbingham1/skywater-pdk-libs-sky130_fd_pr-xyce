* SKY130 Spice File.
* Fast    Varactor Parameters
.param
+  cnwvc_tox='41.6503*1.024*0.952'
+  cnwvc_cdepmult=1.1
+  cnwvc_cintmult=1.05
+  cnwvc_vt1='0.3333-0.112'
+  cnwvc_vt2='0.2380952-0.112'
+  cnwvc_vtr='0.16-0.112'
+  cnwvc_dwc=0.02
+  cnwvc_dlc=0.01
+  cnwvc_dld=0.0008
+  cnwvc2_tox='41.7642*1.017*0.95'
+  cnwvc2_cdepmult=1.05
+  cnwvc2_cintmult=1.05
+  cnwvc2_vt1='0.2-0.074'
+  cnwvc2_vt2='0.33-0.074'
+  cnwvc2_vtr='0.14-0.074'
+  cnwvc2_dwc=0.02
+  cnwvc2_dlc=0.01
+  cnwvc2_dld=0.0006
* sky130_fd_pr__model__parasitic__diode_ps2nw Parameters
.param
+  sky130_fd_pr__model__parasitic__diode_ps2nw__ajunction_mult=8.4794e-01 ; Units: farad/meter^2
+  sky130_fd_pr__model__parasitic__diode_ps2nw__pjunction_mult=9.3896e-01 ; Units: farad/meter^2
* sky130_fd_pr__model__parasitic__diode_ps2dn Parameters
+  sky130_fd_pr__model__parasitic__diode_ps2dn__ajunction_mult=7.9605e-01 ; Units: farad/meter
+  sky130_fd_pr__model__parasitic__diode_ps2dn__pjunction_mult=7.9633e-01 ; Units: farad/meter
* sky130_fd_pr__model__parasitic__diode_pw2dn Parameters
+  sky130_fd_pr__model__parasitic__diode_pw2dn__ajunction_mult=7.7428e-01 ; Units: farad/meter
+  sky130_fd_pr__model__parasitic__diode_pw2dn__pjunction_mult=9.1799e-01 ; Units: farad/meter
* sky130_fd_pr__diode_pw2nd_05v5  Parameters
+  sky130_fd_pr__nfet_01v8__ajunction_mult=7.7394e-1
+  sky130_fd_pr__nfet_01v8__pjunction_mult=7.9336e-1
* sky130_fd_pr__diode_pd2nw_05v5_hvt  Parameters
+  sky130_fd_pr__pfet_01v8_hvt__ajunction_mult=0.8902
+  sky130_fd_pr__pfet_01v8_hvt__pjunction_mult=0.93088
+  dkispp=1.1857e+00 dkbfpp=1.4174e+00 dknfpp=1.000
+  dkispp5x=1.2104e+00 dkbfpp5x=1.7922e+00 dknfpp5x=1.0009e+00 dkisepp5x=6.4618e-01
+  cvpp2_nhvnative10x4_cor=1.136
+  cvpp2_nhvnative10x4_sub=1.23e-14
+  cvpp2_phv5x4_cor=1.136
+  cvpp2_phv5x4_sub=1.23e-14
