* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param sky130_fd_pr__pfet_01v8__toxe_slope_spectre=0.0
.param sky130_fd_pr__pfet_01v8__vth0_slope_spectre=0.0
.param sky130_fd_pr__pfet_01v8__voff_slope_spectre=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_slope_spectre=0.0
* statistics {
*   process {
*   }
*   mismatch {
*     vary sky130_fd_pr__pfet_01v8__toxe_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_01v8__vth0_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_01v8__voff_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_01v8__nfactor_slope_spectre dist=gauss std = 1.0
*   }
* }
.subckt sky130_fd_pr__pfet_01v8 d g s b
.param l=1 w=1 ad=0 as=0 pd=0 ps=0 nrd=0 nrs=0 sa=0 sb=0 sd=0 mult=1 nf=1.0
msky130_fd_pr__pfet_01v8 d g s b sky130_fd_pr__pfet_01v8__model l={l} w={w} ad={ad} as={as} pd={pd} ps={ps} nrd={nrd} nrs={nrs} sa={sa} sb={sb} sd={sd} nf={nf}
.model sky130_fd_pr__pfet_01v8__model.0 pmos
* DC IV MOS Parameters
+  lmin=2.0e-05 lmax=1.0e-04 wmin=7e-06 wmax=1.0e-4
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.05956087+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+  k1=0.43448553
+  k2=0.019777346
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=160312.5
+  ua=-5.6585471e-10
+  ub=9.3302446e-19
+  uc=-6.6549964e-11
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0104767
+  a0=1.236661
+  keta=0.0051290095
+  a1=0.0
+  a2=0.9995
+  ags=0.2260578
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.25706245+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.3376708+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.0015228006
+  pdiblc1=0.39
+  pdiblc2=0.0029632464
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=800000000.0
+  pscbe2=9.3760948e-9
+  pvag=0.0
+  delta=0.01
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=4.6464006
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=3.2358e-10
+  bgidl=1181082000.0
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.4485
+  kt2=-0.0075706
+  at=90900.0
+  ute=-0.33954
+  ua1=1.6104e-9
+  ub1=-5.609e-19
+  uc1=-1.0858e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.1 pmos
* DC IV MOS Parameters
+  lmin=8e-06 lmax=2.0e-05 wmin=7e-06 wmax=1.0e-4
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.05956087+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+  k1=0.43448553
+  k2=0.019777346
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=160312.5
+  ua=-5.6585471e-10
+  ub=9.3302446e-19
+  uc=-6.6549964e-11
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0104767
+  a0=1.236661
+  keta=0.0051290095
+  a1=0.0
+  a2=0.9995
+  ags=0.2260578
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.25706245+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.3376708+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.0015228006
+  pdiblc1=0.39
+  pdiblc2=0.0029632464
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=800000000.0
+  pscbe2=9.3760948e-9
+  pvag=0.0
+  delta=0.01
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=4.6464006
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=3.2358e-10
+  bgidl=1181082000.0
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.4485
+  kt2=-0.0075706
+  at=90900.0
+  ute=-0.33954
+  ua1=1.6104e-9
+  ub1=-5.609e-19
+  uc1=-1.0858e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.2 pmos
* DC IV MOS Parameters
+  lmin=4e-06 lmax=8e-06 wmin=7e-06 wmax=1.0e-4
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.06315259668969+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0=2.88343387641138e-8
+  k1=0.43813350754211 lk1=-2.92859199323285e-8
+  k2=0.018505134186116 lk2=1.0213301175319e-8
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=267935.304375 lvsat=-0.863994582048848
+  ua=-5.7735106104059e-10 lua=9.22925681976438e-17
+  ub=9.2801494195413e-19 lub=4.02163507580296e-26
+  uc=-7.3225399476844e-11 luc=5.3590315902878e-17
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.010287384564 lu0=1.51982204842276e-9
+  a0=1.328364188802 la0=-7.3619209926419e-7
+  keta=0.0214568259084065 lketa=-1.31079514192891e-07 wketa=-1.32348898008484e-23 pketa=1.0097419586829e-28
+  a1=0.0
+  a2=1.2003959015 la2=-1.61278988649118e-6
+  ags=0.15348247893312 lags=5.8263380662106e-7
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.26700524634887+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff=7.98206497751723e-8
+  nfactor={1.1833079277709+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.23922328590075e-6
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-0.433600672985592 lpclm=3.49316602446345e-06 wpclm=1.95214624562515e-22 ppclm=-3.78653234506086e-28
+  pdiblc1=0.39
+  pdiblc2=0.00578918120501261 lpdiblc2=-2.26865707034236e-8
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=800000000.0
+  pscbe2=1.01417218694784e-08 lpscbe2=-6.14644492624777e-15
+  pvag=0.0
+  delta=0.01
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=3.2444736759574 lbeta0=1.12546525230909e-5
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=6.3172955084477e-10 lagidl=-2.4738208963872e-15
+  bgidl=1363431030.754 lbgidl=-1463.89583070474
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.43157364924622 lkt1=-1.35884540735137e-7
+  kt2=0.00980381507592701 lkt2=-1.39481595736561e-7
+  at=87860.10766631 lat=0.0244042191761553
+  ute=-0.47442366324068 lute=1.08284442989222e-6
+  ua1=1.2238699414329e-09 lua1=3.10305867181598e-15
+  ub1=-2.9939625202016e-19 lub1=-2.09934895073718e-24
+  uc1=-8.830298756836e-11 luc1=-1.62783612477057e-16
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.3 pmos
* DC IV MOS Parameters
+  lmin=2e-06 lmax=4e-06 wmin=7e-06 wmax=1.0e-4
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.064659692724+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0=3.49049035051586e-8
+  k1=0.4242721924985 lk1=2.65472907275519e-8
+  k2=0.023299152360404 lk2=-9.09694650249498e-9
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=53437.5
+  ua=-2.310026979311e-10 lua=-1.30279448222702e-15
+  ub=7.5275815268718e-19 lub=7.46148594843831e-25
+  uc=-8.0891709259708e-11 luc=8.44701197125367e-17
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0121662223152 lu0=-6.04811386735782e-9
+  a0=1.171560344358 la0=-1.04588095489892e-7
+  keta=-0.005464761922144 lketa=-2.2639681470487e-8
+  a1=0.0
+  a2=0.8
+  ags=0.0945043548257399 lags=8.20196982788097e-7
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.25410325634546+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff=2.78515888653169e-8
+  nfactor={1.514261668126+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor=-9.38544088047108e-8
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.160612523 leta0=-3.24706275293724e-7
+  etab=-0.140472582563983 letab=2.83862716896731e-7
+  dsub=0.8641982 ldsub=-1.2253066992216e-6
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.46461195637154 lpclm=-1.24823668035527e-7
+  pdiblc1=0.39
+  pdiblc2=-2.158869170794e-05 lpdiblc2=7.19140711328042e-10
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=800446289.17922 lpscbe1=-1.79764745842795
+  pscbe2=8.2864339326498e-09 lpscbe2=1.3266326198426e-15
+  pvag=0.0
+  delta=0.01
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=3.8949963916396 lbeta0=8.6343548305956e-6
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-1.249374783754e-11 lagidl=1.21102820025557e-16 pagidl=9.4039548065783e-38
+  bgidl=917252411.2336 lbgidl=333.306294579995
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.46636744099546 lkt1=4.26443490530082e-9
+  kt2=-0.005478318739886 lkt2=-7.79253441120721e-8
+  at=107038.244165516 lat=-0.0528450845050085
+  ute=-0.17571011240618 lute=-1.20370168306536e-7
+  ua1=2.345249984031e-09 lua1=-1.41384668320866e-15
+  ub1=-1.03151249939108e-18 lub1=8.49606508277918e-25 wub1=1.46936793852786e-39
+  uc1=-2.42518521215026e-10 luc1=4.5839470646531e-16
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.4 pmos
* DC IV MOS Parameters
+  lmin=1e-06 lmax=2e-06 wmin=7e-06 wmax=1.0e-4
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.0639605684452+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0=3.34870878572444e-8
+  k1=0.354542539783 lk1=1.67958189678753e-7
+  k2=0.051575195178736 lk2=-6.64404220255585e-08 pk2=5.04870979341448e-29
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=35126.46375 lvsat=0.037134561782565
+  ua=-7.4823552751872e-10 lua=-2.53852510617286e-16
+  ub=1.05727653665008e-18 lub=1.28588966387678e-25
+  uc=-4.298706539394e-11 luc=7.59995680848559e-18
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0097856841752 lu0=-1.2204110858955e-9
+  a0=1.293571997704 la0=-3.52026264335739e-7
+  keta=-0.006680825932652 lketa=-2.01735182499449e-8
+  a1=0.0
+  a2=0.6972012 la2=2.084747328144e-7
+  ags=0.3705824317914 lags=2.60313955638662e-7
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.2479929006116+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff=1.54598607613175e-8
+  nfactor={1.2665691307516+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor=4.08463084680124e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=-0.502700126 leta0=1.02048381712649e-06 weta0=-1.96868985787621e-22 peta0=7.13130258319795e-28
+  etab=7.64532070406077 letab=-1.55056326388588e-05 wetab=2.59238403974119e-21 petab=4.23144989560551e-27
+  dsub=0.26
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.18260436541916 lpclm=4.47084342324809e-7
+  pdiblc1=0.40860196713388 lpdiblc1=-3.77245661239032e-8
+  pdiblc2=0.00023332426360864 lpdiblc2=2.02180296901481e-10
+  pdiblcb=-0.0499342085713219 lpdiblcb=5.0566275772138e-8
+  drout=0.40005836936472 ldrout=3.2435970762878e-7
+  pscbe1=799107421.64156 lpscbe1=0.917559841535876
+  pscbe2=8.9458121167096e-09 lpscbe2=-1.05784248924693e-17
+  pvag=0.0
+  delta=0.01
+  alpha0=-4.5896723869156e-05 lalpha0=9.3078208044762e-11 walpha0=8.66662311998434e-27 palpha0=3.01759744206368e-32
+  alpha1=2.027988e-10 lalpha1=-2.084747328144e-16
+  beta0=-14.198337403152 lbeta0=4.53274186464274e-05 pbeta0=-2.58493941422821e-26
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-7.724678704e-11 lagidl=2.52421206491676e-16
+  bgidl=797814915.1704 lbgidl=575.524103346211
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.45620503904216 lkt1=-1.63447943071678e-8
+  kt2=-0.040349144324356 lkt2=-7.20772827667392e-9
+  at=70857.671813008 lat=0.0205286820590095
+  ute=-0.16467132300088 lute=-1.42756700755011e-7
+  ua1=1.4159172613352e-09 lua1=4.7082892642575e-16
+  ub1=-8.95996213599985e-21 lub1=-1.22411776664494e-24
+  uc1=-2.1606649321236e-11 luc1=1.03880812071668e-17
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=2.745e-6
+  sbref=2.74e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.5 pmos
* DC IV MOS Parameters
+  lmin=5e-07 lmax=1e-06 wmin=7e-06 wmax=1.0e-4
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.0624003766936+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0=3.18832294589003e-8
+  k1=0.56285163226288 lk1=-4.61810576814534e-8
+  k2=-0.036139298542928 lk2=2.37290249463875e-08 pk2=1.26217744835362e-29
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=59746.9366392 lvsat=0.0118250110981421
+  ua=-6.448941519468e-10 lua=-3.60086204608713e-16
+  ub=1.00672124302384e-18 lub=1.80559201571929e-25
+  uc=-5.9342542976688e-11 luc=2.44131914978195e-17
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0102386419232 lu0=-1.68604621534652e-9
+  a0=0.99456229288 la0=-4.46478758931254e-8
+  keta=-0.0433129398494 lketa=1.7483855271105e-8
+  a1=0.0
+  a2=1.0055976 la2=-1.085530656288e-7
+  ags=0.39664972986984 lags=2.33517086021603e-7
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.22937597595944+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff=-3.67811437800722e-9
+  nfactor={1.6385354519392+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor=2.60861700951257e-8
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.49
+  etab=-15.2926033993656 letab=8.07427808437425e-6
+  dsub=0.21844986818264 ldsub=4.27130369066643e-8
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.61161503644472 lpclm=6.06652063858516e-9
+  pdiblc1=0.723599095127128 lpdiblc1=-3.61537833735426e-7
+  pdiblc2=0.00043
+  pdiblcb=0.236063617142644 lpdiblcb=-2.4343605708791e-07 wpdiblcb=2.31610571514848e-23 ppdiblcb=9.93964740578475e-29
+  drout=0.41525382127056 ldrout=3.08738965415e-7
+  pscbe1=800000000.0
+  pscbe2=8.7131987305096e-09 lpscbe2=2.28545344760497e-16
+  pvag=0.0
+  delta=0.01
+  alpha0=9.1793747738312e-05 lalpha0=-4.84659444820559e-11
+  alpha1=-1.055976e-10 lalpha1=1.085530656288e-16
+  beta0=51.5327469369792 lbeta0=-2.22433472822154e-05 wbeta0=5.42101086242752e-20
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=3.2711551052e-10 lagidl=-1.63258383052434e-16
+  bgidl=1718213903.2296 lbgidl=-370.63501159079
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.43371464300408 lkt1=-3.94646515495619e-8
+  kt2=-0.03909512541676 lkt2=-8.49684466545573e-9
+  at=107540.83678144 lat=-0.017181171330559
+  ute=-0.23309857548808 lute=-7.24143063251996e-8
+  ua1=3.3723123594224e-09 lua1=-1.54032175766671e-15
+  ub1=-2.9027539688824e-18 lub1=1.75066774676228e-24 pub1=1.40129846432482e-45
+  uc1=-4.9327926350544e-11 luc1=3.8885221337971e-17 wuc1=2.46519032881566e-32 puc1=1.17549435082229e-38
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.745e-6
+  sbref=1.74e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.6 pmos
* DC IV MOS Parameters
+  lmin=2.5e-07 lmax=5e-07 wmin=7e-06 wmax=1.0e-4
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.0124465448592+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0=5.50820569631932e-9
+  k1=0.0870956844758403 lk1=2.0501237367873e-7
+  k2=0.14027851671536 lk2=-6.94174644962055e-08 wk2=5.29395592033938e-23 pk2=1.26217744835362e-29
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=61648.1343216 lvsat=0.0108212015362071
+  ua=-5.18986362291201e-10 lua=-4.26564006653394e-16
+  ub=7.784653081888e-19 lub=3.01075596093612e-25
+  uc=-2.77829419541042e-11 luc=7.75010087310758e-18
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.01008388675232 lu0=-1.60433734218393e-9
+  a0=1.19308860166064 la0=-1.49467384613598e-7
+  keta=0.069579111951392 lketa=-4.21217933750916e-08 pketa=-6.31088724176809e-30
+  a1=0.0
+  a2=0.8
+  ags=-0.50603033730192 lags=7.10121329327486e-7
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20612908974192+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff=-1.59521913382231e-8
+  nfactor={1.3360896749344+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor=1.85773911004336e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=1.03299080334588 leta0=-2.86692628276985e-7
+  etab=0.0054650329623552 letab=-2.918471073728e-09 wetab=8.27180612553028e-25 petab=9.86076131526265e-31
+  dsub=0.1689577833808 ldsub=6.88442637770182e-8
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.45686117965856 lpclm=8.77746999753961e-8
+  pdiblc1=-0.387531337591376 lpdiblc1=2.25125701174751e-07 wpdiblc1=-1.05879118406788e-22 ppdiblc1=-2.52435489670724e-29
+  pdiblc2=-0.010312532689536 lpdiblc2=5.67192834968273e-09 wpdiblc2=-3.30872245021211e-24 ppdiblc2=-3.15544362088405e-30
+  pdiblcb=-0.3917928 lpdiblcb=8.80645968864e-8
+  drout=1.59065746041392 ldrout=-3.11860051209025e-7
+  pscbe1=800003936.31008 lpscbe1=-0.00207832448649015
+  pscbe2=9.44025152052e-09 lpscbe2=-1.55329803731514e-16
+  pvag=0.0
+  delta=0.01
+  alpha0=-8.83801750964e-09 lalpha0=4.7191659888798e-15 walpha0=3.74708929979981e-30 palpha0=-9.4039548065783e-38
+  alpha1=2.111952e-10 lalpha1=-5.87097312576e-17
+  beta0=2.5236342748896 lbeta0=3.63287609401599e-6
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-2.83257415536e-10 lagidl=1.59011197430022e-16 wagidl=-9.86076131526265e-32 pagidl=-1.17549435082229e-38
+  bgidl=408956901.8912 lbgidl=320.636974031869
+  cgidl=560.212159639584 lcgidl=-0.000137388897743785
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.45237314112 lkt1=-2.96131884463334e-8
+  kt2=0.019059258944 lkt2=-3.92016617553247e-8
+  at=61656.576 lat=0.007045167750912
+  ute=-0.378311652 lute=4.25645551617605e-9
+  ua1=8.111838232e-10 lua1=-1.88076624083722e-16
+  ub1=4.3553038656e-19 lub1=-1.19063334990412e-26
+  uc1=9.12517592000001e-12 luc1=8.02268477635104e-18
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.245e-6
+  sbref=1.24e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.7 pmos
* DC IV MOS Parameters
+  lmin=1.8e-07 lmax=2.5e-07 wmin=7e-06 wmax=1.0e-4
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.898146022857143+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0=-2.62659678139886e-8
+  k1=0.237429301868572 lk1=1.6322143204696e-7
+  k2=0.109518224818628 lk2=-6.08664724724169e-8
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=133265.365337143 lvsat=-0.00908752927934167
+  ua=-1.39996641489714e-09 lua=-1.81662123789573e-16
+  ub=1.25608315379429e-18 lub=1.68303566429434e-25
+  uc=-7.82622461557714e-14 luc=4.85323704544066e-20
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.00603840557371429 lu0=-4.79742120305688e-10
+  a0=1.02350097064057 la0=-1.02324058241591e-7
+  keta=-0.255963735087943 lketa=4.8375211587679e-8
+  a1=0.0
+  a2=0.884075316078286 la2=-2.33719289659705e-8
+  ags=4.42094239888 lags=-6.59517967658253e-7
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.113778264501143+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff=-4.16246125452564e-8
+  nfactor={1.98383861314286+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor=5.70747916964326e-9
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=-0.500893996689577 leta0=1.39708939515272e-07 weta0=2.64697796016969e-23 peta0=7.25752032803331e-29
+  etab=0.150037252567531 letab=-4.31078132573317e-08 wetab=-7.94093388050907e-23 petab=-1.26217744835362e-29
+  dsub=0.813536297068 ldsub=-1.10340828085859e-7
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=1.17740760672457 lpclm=-1.1252856019183e-7
+  pdiblc1=1.12264261148057 lpdiblc1=-1.94684534579861e-7
+  pdiblc2=0.0276727296547886 lpdiblc2=-4.88751875889137e-9
+  pdiblcb=-0.075
+  drout=-0.96013260794457 ldrout=3.97228978313815e-7
+  pscbe1=799985941.749714 lpscbe1=0.00292394736050028
+  pscbe2=7.93289394397143e-09 lpscbe2=2.6369751425807e-16
+  pvag=0.0
+  delta=0.01
+  alpha0=3.20214911058571e-08 lalpha0=-6.63928709212501e-15
+  alpha1=-2.97125714285714e-10 lalpha1=8.25973830628571e-17
+  beta0=36.35176297792 lbeta0=-5.77093774788203e-06 wbeta0=5.42101086242752e-20
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=8.10931774104571e-10 lagidl=-1.45160267019782e-16
+  bgidl=3233344075.35429 lbgidl=-464.508767544787
+  cgidl=-629.329141569943 lcgidl=0.000193289309496849 pcgidl=5.16987882845642e-26
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=0.132422399428571 lkt1=-1.9217933117235e-7
+  kt2=-0.12196
+  at=232591.6 lat=-0.0404727177008
+  ute=-0.5501892 lute=5.20363513296e-8
+  ua1=1.3462e-10
+  ub1=3.927e-19
+  uc1=3.7985e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.1e-6
+  sbref=1.1e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.8 pmos
* DC IV MOS Parameters
+  lmin=1.5e-07 lmax=1.8e-07 wmin=7e-06 wmax=1.0e-4
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.864818294533334+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0=-3.3197735372601e-8
+  k1=-0.556924842106668 lk1=3.28437561744082e-7
+  k2=0.480439082930667 lk2=-1.38013559909424e-7
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=276959.752986667 lvsat=-0.0389742375777909
+  ua=-8.68544388573337e-10 lua=-2.92191528200609e-16
+  ub=7.07058731760001e-19 lub=2.82494057919502e-25
+  uc=2.97575570237334e-13 luc=-2.96373853015625e-20
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.00695832713466667 lu0=-6.71074765925051e-10
+  a0=-1.110903038712 la0=3.41606362855632e-7
+  keta=-0.108048302823173 lketa=1.76105766617942e-8
+  a1=0.0
+  a2=-0.579795937516 la2=2.81095725326598e-7
+  ags=1.25
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.562279240085334+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff=5.16582083645482e-8
+  nfactor={2.58027797133334+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor=-1.18344750061677e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=-0.807748139174667 leta0=2.03530918902461e-7
+  etab=-0.292823200157334 letab=4.90018465840075e-8
+  dsub=0.419602642290667 ldsub=-2.84073550960312e-8
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=2.47623844447867 lpclm=-3.82669788474629e-7
+  pdiblc1=1.17802969655867 lpdiblc1=-2.06204383631084e-7
+  pdiblc2=0.0263847365516267 lpdiblc2=-4.61963164935093e-9
+  pdiblcb=-0.501673309421254 lpdiblcb=8.87429282799077e-8
+  drout=0.651497248421334 ldrout=6.20293077479838e-8
+  pscbe1=883573612.777333 lpscbe1=-17.382308574332
+  pscbe2=1.035851282288e-08 lpscbe2=-2.40802105128364e-16
+  pvag=0.0
+  delta=0.01
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=15.8918131392 lbeta0=-1.51551370082633e-6
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=1.90167027089333e-10 lagidl=-1.60486488175762e-17
+  bgidl=728006451.213334 lbgidl=56.5713942250411
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-2.06952384 lkt1=2.6579906327392e-7
+  kt2=-0.12196
+  at=38000.0
+  ute=-0.3
+  ua1=1.3462e-10
+  ub1=3.927e-19
+  uc1=3.7985e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.04e-6
+  sbref=1.04e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.9 pmos
* DC IV MOS Parameters
+  lmin=2.0e-05 lmax=1.0e-04 wmin=5.0e-06 wmax=7.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.07086482305516+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} wvth0=7.8962545500707e-8
+  k1=0.444261859177239 wk1=-6.82914935793182e-8
+  k2=0.0156234349599887 wk2=2.90166977783888e-8
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=160312.5
+  ua=-5.9084498548094e-10 wua=1.74566875420409e-16
+  ub=9.43061924020675e-19 wub=-7.01156228778009e-26
+  uc=-7.48309447284178e-11 wuc=5.78458981886402e-17
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.01077283229668 wu0=-2.06860023539657e-9
+  a0=1.3417730091448 wa0=-7.34248608806413e-7
+  keta=0.0300324686133604 wketa=-1.73960429043486e-7
+  a1=0.0
+  a2=1.22315994939213 wa2=-1.56235246593619e-6
+  ags=0.221448331298841 wags=3.2198946711221e-8
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.269379060845788+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} wvoff=8.60363573326029e-8
+  nfactor={0.77913338195144+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} wnfactor=3.90160292344455e-6
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-0.561230562720794 wpclm=3.93105295466484e-6
+  pdiblc1=0.39
+  pdiblc2=0.00992920113806031 wpdiblc2=-4.86599258927995e-8
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=800000000.0
+  pscbe2=1.01214877089399e-08 wpscbe2=-5.20686181204394e-15
+  pvag=0.0
+  delta=0.01
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=0.396943770666869 wbeta0=2.96841225898604e-5
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-2.303023734492e-09 wagidl=1.83478572394113e-14
+  bgidl=280422540.76566 wbgidl=6291.45956139177
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.479524993031196 wkt1=2.16721744325171e-7
+  kt2=0.0995282524544426 wkt2=-7.48127488564214e-7
+  at=93143.42649 wat=-0.0156712139045194
+  ute=-0.775332799574229 wute=3.04418362296198e-6
+  ua1=7.4055649630191e-10 wua1=6.07619802595331e-15
+  ub1=-8.34809952239245e-20 wub1=-3.33495899209456e-24
+  uc1=-6.58246062190426e-10 wuc1=3.83963302342972e-15
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.10 pmos
* DC IV MOS Parameters
+  lmin=8e-06 lmax=2.0e-05 wmin=5.0e-06 wmax=7.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.07086482305516+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} wvth0=7.89625455007036e-8
+  k1=0.444261859177239 wk1=-6.82914935793165e-8
+  k2=0.0156234349599887 wk2=2.90166977783888e-8
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=160312.5
+  ua=-5.9084498548094e-10 wua=1.74566875420409e-16
+  ub=9.43061924020676e-19 wub=-7.01156228778009e-26
+  uc=-7.48309447284178e-11 wuc=5.78458981886404e-17
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.01077283229668 wu0=-2.06860023539657e-9
+  a0=1.3417730091448 wa0=-7.34248608806417e-7
+  keta=0.0300324686133604 wketa=-1.73960429043486e-7
+  a1=0.0
+  a2=1.22315994939213 wa2=-1.56235246593619e-6
+  ags=0.221448331298841 wags=3.21989467112193e-8
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.269379060845788+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} wvoff=8.60363573326021e-8
+  nfactor={0.77913338195144+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} wnfactor=3.90160292344455e-6
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-0.561230562720794 wpclm=3.93105295466484e-6
+  pdiblc1=0.39
+  pdiblc2=0.00992920113806031 wpdiblc2=-4.86599258927995e-8
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=800000000.0
+  pscbe2=1.01214877089399e-08 wpscbe2=-5.20686181204391e-15
+  pvag=0.0
+  delta=0.01
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=0.396943770666869 wbeta0=2.96841225898604e-5
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-2.303023734492e-09 wagidl=1.83478572394113e-14
+  bgidl=280422540.76566 wbgidl=6291.45956139178
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.479524993031196 wkt1=2.16721744325171e-7
+  kt2=0.0995282524544426 wkt2=-7.48127488564214e-7
+  at=93143.4264900001 wat=-0.0156712139045192
+  ute=-0.775332799574229 wute=3.04418362296198e-6
+  ua1=7.40556496301911e-10 wua1=6.07619802595332e-15
+  ub1=-8.34809952239249e-20 wub1=-3.33495899209456e-24
+  uc1=-6.58246062190426e-10 wuc1=3.83963302342972e-15
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.11 pmos
* DC IV MOS Parameters
+  lmin=4e-06 lmax=8e-06 wmin=5.0e-06 wmax=7.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.07223615742125+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0=1.10090558348923e-08 wvth0=6.34522342824343e-08 pvth0=1.24516592336558e-13
+  k1=0.417770816632546 lk1=2.12669771656287e-07 wk1=1.42241382250679e-07 pk1=-1.69015540076871e-12
+  k2=0.0238580777309972 lk2=-6.61076133499426e-08 wk2=-3.73924100854532e-08 pk2=5.33131521021628e-13
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=276284.616584665 lvsat=-0.93102276027629 wvsat=-0.0583232203847563 pvsat=4.68218113370182e-7
+  ua=-2.35694865293704e-10 lua=-2.85114090306169e-15 wua=-2.38660252485197e-15 pua=2.05610372113539e-20
+  ub=6.95634019930934e-19 lub=1.98634824489759e-24 wub=1.62327188012964e-24 pub=-1.35944945534938e-29
+  uc=-9.30449199971931e-11 luc=1.46221574890024e-16 wuc=1.38447124050586e-16 puc=-6.47065674004993e-22
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0119891938576625 lu0=-9.76493601522924e-09 wu0=-1.18878053658379e-08 pu0=7.88284609567216e-14
+  a0=1.62073496518233 la0=-2.2395032355258e-06 wa0=-2.04232454083508e-06 pa0=1.0501217885415e-11
+  keta=0.0730525366663151 lketa=-3.45364590088304e-07 wketa=-3.60416275481751e-07 pketa=1.49686529773623e-12
+  a1=0.0
+  a2=1.64928074895016 la2=-3.42089266540226e-06 wa2=-3.13563671207655e-06 pa2=1.26303070486038e-11
+  ags=0.178746859393834 lags=3.42806904035739e-07 wags=-1.76481606208101e-07 pags=1.67528497466966e-12
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.300303243065369+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff=2.4825896376861e-07 wvoff=2.32599566539056e-07 pvoff=-1.17660768475091e-12
+  nfactor={0.220392379615385+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor=4.48556606186184e-06 wnfactor=6.72634275934427e-06 pnfactor=-2.26769775057249e-11
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-1.54648460380339 lpclm=7.90960761876255e-06 wpclm=7.77393072983995e-06 ppclm=-3.08505766645725e-11
+  pdiblc1=0.39
+  pdiblc2=0.0196457120200023 lpdiblc2=-7.80040327620994e-08 wpdiblc2=-9.67933022740883e-08 ppdiblc2=3.8641416798847e-13
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=800000000.0
+  pscbe2=1.37702318462581e-08 lpscbe2=-2.92920741494609e-14 wpscbe2=-2.5346565289419e-14 ppscbe2=1.61681297839925e-19
+  pvag=0.0
+  delta=0.01
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=-3.69914660914365 lbeta0=3.28833644160343e-05 wbeta0=4.85039109793066e-05 pbeta0=-1.51085035353014e-10
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-2.47913390022633e-09 lagidl=1.41381029719326e-15 wagidl=2.17306012863772e-14 pagidl=-2.71566286161137e-20
+  bgidl=777327945.574429 lbgidl=-3989.15062693994 wbgidl=4094.15991960932 pbgidl=0.0176398951566339
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.48771334605363 lkt1=6.57359998038579e-08 wkt1=3.92157800188839e-07 pkt1=-1.40839855124088e-12
+  kt2=0.157972924743658 lkt2=-4.69193127801751e-07 wkt2=-1.03501934295391e-06 pkt2=2.30316436433822e-12
+  at=93374.1429062892 lat=-0.00185218862137315 wat=-0.038517698755876 pat=1.83411306228872e-7
+  ute=-1.3490524551764 lute=4.60581451053834e-06 wute=6.10962514108318e-06 pute=-2.46093277221788e-11
+  ua1=-5.22609029505498e-11 lua1=6.36472856738995e-15 wua1=8.91427444653555e-15 pua1=-2.27840434475172e-20
+  ub1=4.0123251243327e-19 lub1=-3.89127422290987e-24 wub1=-4.89416670630863e-24 pub1=1.25173008192179e-29
+  uc1=-1.19556152959347e-09 luc1=4.31356212452607e-15 wuc1=7.73463518284561e-15 puc1=-3.12690305957649e-20
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.12 pmos
* DC IV MOS Parameters
+  lmin=2e-06 lmax=4e-06 wmin=5.0e-06 wmax=7.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.07814560900045+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0=3.48122558825018e-08 wvth0=9.42044143673463e-08 pvth0=6.47179980677002e-16
+  k1=0.515778983259007 lk1=-1.82105947417098e-07 wk1=-6.39210822425474e-07 pk1=1.45752470224038e-12
+  k2=-0.00871027749946673 lk2=6.50773306981034e-08 wk2=2.23598421669588e-07 pk2=-5.18136417397698e-13
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=36738.8755806705 lvsat=0.0338646099389072 wvsat=0.116646440769514 pvsat=-2.36557582123284e-7
+  ua=-1.29668796248456e-09 lua=1.42252656050593e-15 wua=7.4442295346667e-15 pua=-1.90374363544026e-20
+  ub=1.41578715713785e-18 lub=-9.14419949934225e-25 wub=-4.63151763606348e-24 pub=1.1599722560258e-29
+  uc=-6.22940609826625e-11 luc=2.23574837898034e-17 wuc=-1.29911867212817e-16 puc=4.33881122496101e-22
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.00846000544531283 lu0=4.45059255945454e-09 wu0=2.58893784144182e-08 pu0=-7.3337581983945e-14
+  a0=1.09670762129305 la0=-1.28727382667908e-07 wa0=5.22875627846678e-07 pa0=1.68622388366885e-13
+  keta=-0.00898959240077878 lketa=-1.48998787115987e-08 wketa=2.46223233317775e-08 pketa=-5.40655578214769e-14
+  a1=0.0
+  a2=0.8
+  ags=-0.0697841063676887 lags=1.34388665175156e-06 wags=1.14761933537058e-06 pags=-3.65817772879797e-12
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.254605045408927+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff=6.41871719868327e-08 wvoff=3.50519340998654e-09 pvoff=-2.53818298919492e-13
+  nfactor={0.928009366123206+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.63529333161216e-06 wnfactor=4.09520225764236e-06 pnfactor=-1.20787751385556e-11
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.160612527827676 leta0=-3.24706294739544e-07 weta0=-3.37232077556222e-14 peta0=1.35836677596333e-19
+  etab=-0.140472582538707 letab=2.83862716794921e-07 wetab=-1.76561476756317e-16 petab=7.11186303100938e-22
+  dsub=0.8641982 ldsub=-1.2253066992216e-6
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=1.02803934334819 lpclm=-2.46054394607662e-06 wpclm=-3.93576127425305e-06 ppclm=1.63159222116101e-11
+  pdiblc1=0.39
+  pdiblc2=0.000471776621692122 lpdiblc2=-7.71651064930893e-10 wpdiblc2=-3.44635021197535e-09 ppdiblc2=1.04137652457033e-14
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=772367617.505149 lpscbe1=111.302905100674 wpscbe1=196.14053409842 ppscbe1=-0.000790051717662034
+  pscbe2=5.32147077870037e-09 lpscbe2=4.73943404552879e-15 wpscbe2=2.07114304888857e-14 ppscbe2=-2.3839756459137e-20
+  pvag=0.0
+  delta=0.01
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=0.927342922078175 lbeta0=1.42479201021472e-05 wbeta0=2.07302233985774e-05 pbeta0=-3.92129550620875e-11
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-3.90410346558025e-09 lagidl=7.15357060680406e-15 wagidl=2.71844201677642e-14 pagidl=-4.91245456245139e-20
+  bgidl=-859463748.071624 lbgidl=2603.82667356605 wbgidl=12411.0592008247 pbgidl=-0.0158604753453102
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.481217021021369 lkt1=3.95688805298159e-08 wkt1=1.03730140486261e-07 pkt1=-2.46615399090809e-13
+  kt2=0.125810850004869 lkt2=-3.39644676698805e-07 wkt2=-9.17106335294092e-07 pkt2=1.82821218444057e-12
+  at=101384.103772023 lat=-0.0341162148690159 wat=0.0394963882024144 pat=-1.30828499870078e-7
+  ute=-0.326588997179381 lute=4.87343971287855e-07 wute=1.05394818483942e-06 pute=-4.24512161055237e-12
+  ua1=1.03033322827696e-09 lua1=2.00405239793511e-15 wua1=9.18520924929356e-15 pua1=-2.38753655818088e-20
+  ub1=-3.55146725872715e-19 lub1=-8.44587727564221e-25 wub1=-4.72468019868216e-24 pub1=1.18346112003366e-29
+  uc1=9.56376815881239e-11 luc1=-8.87372803722882e-16 wuc1=-2.36215370144274e-15 puc1=9.40071386868202e-21
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.13 pmos
* DC IV MOS Parameters
+  lmin=1e-06 lmax=2e-06 wmin=5.0e-06 wmax=7.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.08398954705592+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0=4.66636921317415e-08 wvth0=1.39910270961289e-07 pvth0=-9.20437487215619e-14
+  k1=0.324438550909221 lk1=2.05930153303079e-07 wk1=2.10288169067784e-07 pk1=-2.65249058520049e-13
+  k2=0.0663841555451893 lk2=-8.72132783832624e-08 wk2=-1.03446396233932e-07 pk2=1.45106548772826e-13
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=-75792.7316435821 lvsat=0.262077359010405 wvsat=0.774814082332604 pvsat=-1.57131366120153e-6
+  ua=-5.35045536740578e-10 lua=-1.22075139193765e-16 wua=-1.48921569869969e-15 pua=-9.20516622478376e-22
+  ub=9.29006108501381e-19 lub=7.2766175327952e-26 wub=8.96019248280581e-25 pub=3.89944089250831e-31
+  uc=-5.36296885389152e-11 luc=4.78624044635334e-18 wuc=7.43428967044496e-17 puc=1.96549123290512e-23
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0110470217550709 lu0=-7.95845472539097e-10 wu0=-8.81093769199706e-09 pu0=-2.96575732392798e-15
+  a0=0.462190463499744 la0=1.15806579913102e-06 wa0=5.80752608425444e-06 pa0=-1.05485853214226e-11
+  keta=-0.0724434340750336 lketa=1.1378375075769e-07 wketa=4.59377609969449e-07 pketa=-9.35744062059234e-13
+  a1=0.0
+  a2=0.440955032155319 la2=7.28138886249397e-07 wa2=1.78997998214212e-06 pa2=-3.63005792402443e-12
+  ags=1.94258197034248 lags=-2.73716760342374e-06 wags=-1.09810333149983e-05 pags=2.09385843023183e-11
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.208292079609894+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff=-2.9734966898017e-08 wvoff=-2.77325805358916e-07 pvoff=3.15703596611859e-13
+  nfactor={2.0655144687291+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor=-6.71553366411369e-07 wnfactor=-5.58094653213443e-06 pnfactor=7.54433849332621e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=-0.502700135655352 leta0=1.02048382705207e-06 weta0=6.74464157296201e-14 peta0=-6.9334105233868e-20
+  etab=26.7021061400892 letab=-5.41525648217497e-05 wetab=-0.000133119120341906 petab=2.69963978624295e-10
+  dsub=0.26
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-1.51475066928458 lpclm=2.69620368606248e-06 wpclm=1.18566906200502e-05 ppclm=-1.57109807206142e-11
+  pdiblc1=0.432576358597428 lpdiblc1=-8.63443443192817e-08 wpdiblc1=-1.67470527129217e-07 ppdiblc1=3.39628219371727e-13
+  pdiblc2=-0.000256928577458731 lpdiblc2=7.06154334484646e-10 wpdiblc2=3.42460837201985e-09 ppdiblc2=-3.52045631113595e-15
+  pdiblcb=-0.0499802644894317 lpdiblcb=5.06596766213938e-08 wpdiblcb=3.21718651128339e-10 ppdiblcb=-6.52441563864533e-16
+  drout=0.646834960076699 ldrout=-1.76100257016025e-07 wdrout=-1.72383127190205e-06 pdrout=3.49590913344211e-12
+  pscbe1=855264764.989703 lpscbe1=-56.8115152322353 wpscbe1=-392.28106819684 ppscbe1=0.000403260230733532
+  pscbe2=1.92379287531711e-09 lpscbe2=1.16298840614551e-14 wpscbe2=4.90515584370729e-14 ppscbe2=-8.13131958565253e-20
+  pvag=0.0
+  delta=0.01
+  alpha0=-0.000160303557730188 lalpha0=3.25093894232929e-10 walpha0=7.99176604879549e-10 palpha0=-1.62072056457647e-15
+  alpha1=4.5904496784468e-10 lalpha1=-7.28138886249397e-16 walpha1=-1.78997998214212e-15 palpha1=3.63005792402443e-21
+  beta0=-68.323656004462 lbeta0=0.000154688114913184 wbeta0=0.000378086578380106 pbeta0=-7.63927354688367e-10
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-1.07716546111186e-09 lagidl=1.4205742569982e-15 wagidl=6.98482410649588e-15 pagidl=-8.16000720741452e-21
+  bgidl=-981367553.268816 lbgidl=2851.04612766028 wbgidl=12428.287337412 pbgidl=-0.0158954137995717
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.455903412914567 lkt1=-1.17668129474825e-08 wkt1=-2.1069767990056e-09 pkt1=-3.19789952816946e-14
+  kt2=-0.0367163772584209 lkt2=-1.00414101355812e-08 wkt2=-2.53763027268e-08 pkt2=1.9794379154492e-14
+  at=-89494.0497550208 lat=0.352982389945985 wat=1.12011966509788 pat=-2.32231953793476e-6
+  ute=0.300064203004743 lute=-7.83501198847148e-07 wute=-3.24635991842258e-06 pute=4.47585161916573e-12
+  ua1=2.24618137811119e-09 lua1=-4.61673059750918e-16 wua1=-5.79972048526692e-15 pua1=6.513892100723e-21
+  ub1=-4.27736023852957e-19 lub1=-6.97377502331863e-25 wub1=2.92531503506435e-24 pub1=-3.67948733375849e-30
+  uc1=-6.80795105722935e-10 luc1=6.87223571750498e-16 wuc1=4.60468990167847e-15 puc1=-4.72796135632456e-21
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=2.745e-6
+  sbref=2.74e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.14 pmos
* DC IV MOS Parameters
+  lmin=5e-07 lmax=1e-06 wmin=5.0e-06 wmax=7.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.06588452666826+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0=2.80519484334661e-08 wvth0=2.43381540565869e-08 pvth0=2.67630005910734e-14
+  k1=0.592920162830969 lk1=-7.00657219731344e-08 wk1=-2.10040478895788e-07 pk1=1.66843747642727e-13
+  k2=-0.0543909295533397 lk2=3.69420597970042e-08 wk2=1.27494800897408e-07 pk2=-9.2298230583826e-14
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=279632.478024475 lvsat=-0.103295491425842 wvsat=-1.53598674568547 pvsat=8.04161860391116e-7
+  ua=-3.55244762087223e-11 lua=-6.35576795167787e-16 wua=-4.2566861798173e-15 pua=1.92440982246474e-21
+  ub=7.17782078541963e-19 lub=2.89901943437875e-25 wub=2.01835338584623e-24 pub=-7.63801936157001e-31
+  uc=-8.36766426936607e-11 luc=3.56741487539818e-17 wuc=1.69983230356963e-16 puc=-7.86622029817287e-23
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0130430010549544 lu0=-2.84768824106778e-09 wu0=-1.95895484049561e-08 pu0=8.11452514566544e-15
+  a0=2.28523043331344 la0=-7.15997413357827e-07 wa0=-9.01582316097228e-06 pa0=4.68963982247954e-12
+  keta=0.0794843762667092 lketa=-4.23962151398977e-08 wketa=-8.57787414178404e-07 pketa=4.18285776784469e-13
+  a1=0.0
+  a2=1.52475384014655 la2=-3.85993282779889e-07 wa2=-3.62650995050102e-06 pa2=1.93802872885352e-12
+  ags=-2.24132075171841 lags=1.5638341880222e-06 wags=1.84272584259168e-05 pags=-9.29278670784154e-12
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.244832686193965+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff=7.82833818312952e-09 wvoff=1.07971183109911e-07 pvoff=-8.0377083970235e-14
+  nfactor={1.04003502020121+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor=3.82627200921925e-07 wnfactor=4.18076024755921e-06 pnfactor=-2.49057893571749e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.49
+  etab=-53.4060920144217 letab=2.81977015827096e-05 wetab=0.000266237666086402 petab=-1.40570005542569e-10
+  dsub=0.199057618246564 ldsub=6.2648037133952e-08 wdsub=1.35462471443922e-07 pdsub=-1.39253795094693e-13
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=1.62211710315261 lpclm=-5.28458741589685e-07 wpclm=-7.05875325486518e-06 ppclm=3.73386859747231e-12
+  pdiblc1=0.624709378761775 lpdiblc1=-2.83854783451988e-07 wpdiblc1=6.90783453358746e-07 ppdiblc1=-5.42646573522135e-13
+  pdiblc2=0.00043
+  pdiblcb=0.236155728978864 lpdiblcb=-2.43484691032092e-07 wpdiblcb=-6.43437302256969e-10 ppdiblcb=3.39727174344073e-16
+  drout=-0.078299360153399 ldrout=5.69329122568673e-07 wdrout=3.44766254380411e-06 pdrout=-1.82032445117804e-12
+  pscbe1=800000000.0
+  pscbe2=-3.88525944403607e-09 lpscbe2=1.76015201371224e-14 wpscbe2=8.80051714644976e-14 ppscbe2=-1.21357042605362e-19
+  pvag=0.0
+  delta=0.01
+  alpha0=0.000320607415460376 lalpha0=-1.69276815275293e-10 walpha0=-1.5983532097591e-09 palpha0=8.43911314514287e-16
+  alpha1=-6.1808993568936e-10 lalpha1=3.79142868964754e-16 walpha1=3.57995996428424e-15 palpha1=-1.89017590162251e-21
+  beta0=158.999009120538 lbeta0=-7.89968569633352e-05 wbeta0=-0.000750693989620188 pbeta0=3.96445523849119e-10
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=9.30173840431013e-10 lagidl=-6.42946456916246e-16 wagidl=-4.21259895390542e-15 pagidl=3.3508093296013e-21
+  bgidl=3146032936.68666 lbgidl=-1391.87204720806 wbgidl=-9973.87593932248 pbgidl=0.00713374122295202
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.423938544205404 lkt1=-4.46263144020773e-08 wkt1=-6.82898842947031e-08 pkt1=3.60562394289908e-14
+  kt2=-0.0372936072334215 lkt2=-9.44802464804029e-09 wkt2=-1.25843110660517e-08 pkt2=6.64436523114243e-15
+  at=431924.18515444 lat=-0.183029298522122 wat=-2.26594491153464 pat=1.15851421406855e-6
+  ute=-0.420594685599676 lute=-4.26725092684692e-08 wute=1.30973386510388e-06 pute=-2.07758117174068e-13
+  ua1=3.18798921225277e-09 lua1=-1.42984021155445e-15 wua1=1.28756947451818e-15 pua1=-7.71756930456557e-22
+  ub1=-2.62027112260764e-18 lub1=1.55652226876677e-24 wub1=-1.97325347100149e-24 pub1=1.35618230765514e-30
+  uc1=-5.0932591102821e-11 luc1=3.97324650711962e-17 wuc1=1.12092126441703e-17 puc1=-5.91832976557027e-24
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.745e-6
+  sbref=1.74e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.15 pmos
* DC IV MOS Parameters
+  lmin=2.5e-07 lmax=5e-07 wmin=5.0e-06 wmax=7.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.04105604595688+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0=1.4942808559632e-08 wvth0=1.99848585813647e-07 pvth0=-6.59044012514779e-14
+  k1=0.0514910163996825 lk1=2.15802370192828e-07 wk1=2.48712570662786e-07 pk1=-7.53723574876054e-14
+  k2=0.159319176640184 lk2=-7.58943117519023e-08 wk2=-1.33006477321721e-07 pk2=4.52433183005357e-14
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=19951.2006467036 lvsat=0.033813106854293 wvsat=0.291269435256539 pvsat=-1.60607476072096e-7
+  ua=-3.14511158059148e-10 lua=-4.88275174990943e-16 wua=-1.42833949673599e-15 pua=4.31076713958006e-22
+  ub=6.55772527240271e-19 lub=3.22642242410553e-25 wub=8.57057195034159e-25 pub=-1.5065148296252e-31
+  uc=-3.40688054573241e-11 luc=9.4818059872429e-18 wuc=4.39092218856572e-17 puc=-1.2096639396981e-23
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.011384104824662 lu0=-1.97181093822812e-09 wu0=-9.08253318083656e-09 pu0=2.566947191513e-15
+  a0=1.27052901763011 la0=-1.80247242294012e-07 wa0=-5.40951677677857e-07 pa0=2.15009377757876e-13
+  keta=0.0364728685250521 lketa=-1.96866551903955e-08 wketa=2.31260094601655e-07 pketa=-1.56718239281297e-13
+  a1=0.0
+  a2=0.786672191085628 la2=3.70497094448905e-09 wa2=9.30999724335609e-08 pa2=-2.58806751368595e-14
+  ags=-0.16130772847994 lags=4.65612271908561e-07 wags=-2.40802262282869e-06 pags=1.70799166252351e-12
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.198053973684804+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff=-1.68702606771574e-08 wvoff=-5.64078527194733e-08 pvoff=6.41307439925072e-15
+  nfactor={1.51612745620061+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor=1.31256107823473e-07 wnfactor=-1.25763451296229e-06 pnfactor=3.80828237100733e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=2.19585075491521 leta0=-9.00668728386175e-07 weta0=-8.1230328353848e-06 peta0=4.28886386068915e-12
+  etab=0.0153311551786357 letab=-8.16879376134646e-09 wetab=-6.89187331738524e-08 petab=3.6675563149573e-14
+  dsub=0.22030846578562 ldsub=5.14278446435005e-08 wdsub=-3.58704656335305e-07 pdsub=1.21660518367205e-13
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.228955171086374 lpclm=2.07114040598104e-07 wpclm=1.59201285461329e-06 ppclm=-8.33632099139008e-13
+  pdiblc1=-0.436001593357444 lpdiblc1=2.76187881295295e-07 wpdiblc1=3.38583746560303e-07 ppdiblc1=-3.56689354729037e-13
+  pdiblc2=-0.0199738913391894 lpdiblc2=1.07730097803959e-08 wpdiblc2=6.74883793526914e-08 ppdiblc2=-3.56330544376688e-14
+  pdiblcb=-0.25320487931064 lpdiblcb=1.48918378174662e-08 wpdiblcb=-9.68090980197671e-07 ppdiblcb=5.11140420452609e-13
+  drout=2.36484797423871 ldrout=-7.20623352222351e-07 wdrout=-5.40802437658572e-06 pdrout=2.85537197454474e-12
+  pscbe1=800013748.334866 lpscbe1=-0.00725895582877456 wpscbe1=-0.0685408413955884 ppscbe1=3.6188741768875e-8
+  pscbe2=6.57523595102706e-08 lpscbe2=-1.91663070193241e-14 wpscbe2=-3.93362159917161e-13 ppscbe2=1.32799131956178e-19
+  pvag=0.0
+  delta=0.01
+  alpha0=-7.80495931169914e-09 lalpha0=4.17372365706541e-15 walpha0=-7.21631667804203e-15 palpha0=3.81012861020606e-21
+  alpha1=2.111952e-10 lalpha1=-5.87097312576e-17
+  beta0=2.53564170559848 lbeta0=3.61392347134402e-06 wbeta0=-8.38766128157084e-08 pbeta0=1.32391502582281e-13
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=2.98733419932844e-10 lagidl=-3.09553492178258e-16 wagidl=-4.06543424255554e-15 pagidl=3.2731081279851e-21
+  bgidl=-99086310.5175924 lbgidl=321.511973884815 wbgidl=3548.88109322333 pbgidl=-6.11221714777108e-6
+  cgidl=485.525039274244 lcgidl=-9.79549944363295e-05 wcgidl=0.000521718828040507 pcgidl=-2.75461280579452e-10
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.477596142685464 lkt1=-1.62957462957877e-08 wkt1=1.76192558395976e-07 pkt1=-9.30275565223751e-14
+  kt2=0.0292038947384611 lkt2=-4.45579077191706e-08 wkt2=-7.08642597504696e-08 pkt2=3.74154787771309e-14
+  at=8508.65142454905 lat=0.0405290223008561 wat=0.371259097775544 pat=-2.33897856399114e-7
+  ute=-0.480706468446889 lute=-1.09342092665347e-08 wute=7.15267952128529e-07 pute=1.06112751285961e-13
+  ua1=9.57125756545949e-10 lua1=-2.51971077302714e-16 wua1=-1.01946164284771e-15 pua1=4.46327815139218e-22
+  ub1=2.99083011414212e-19 lub1=1.51383182528366e-26 wub1=9.53138430053858e-25 pub1=-1.88917499399284e-31
+  uc1=-5.43259176884165e-11 luc1=4.15241007884717e-17 wuc1=4.43230774373703e-16 puc1=-2.34020530100023e-22
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.245e-6
+  sbref=1.24e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.16 pmos
* DC IV MOS Parameters
+  lmin=1.8e-07 lmax=2.5e-07 wmin=5.0e-06 wmax=7.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.849074197505416+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0=-3.84258415276951e-08 wvth0=-3.42785946051707e-07 pvth0=8.49414869927084e-14
+  k1=0.345431055681784 lk1=1.34090566552874e-07 wk1=-7.54434608673133e-07 pk1=2.03490520601628e-13
+  k2=0.0698700846096645 lk2=-5.10285375565221e-08 wk2=2.76957809360206e-07 pk2=-6.87218338255993e-14
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=320137.666771546 lvsat=-0.0496351284908196 wvsat=-1.30537631683593 pvsat=2.83240883260584e-7
+  ua=-1.43135886191672e-09 lua=-1.77804915490984e-16 wua=2.19288554549476e-16 pua=-2.69441127627433e-23
+  ub=9.02727358177202e-19 lub=2.53991762868059e-25 wub=2.46832881852838e-24 pub=-5.9856565903443e-31
+  uc=1.7398130783619e-13 luc=-3.72778200304898e-20 wuc=-1.76202015455572e-18 puc=5.99417835293709e-25
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.00479080498808037 lu0=-1.38952703256473e-10 wu0=8.71497939960255e-09 pu0=-2.38054773569812e-15
+  a0=0.801114070626047 la0=-4.97555200062483e-08 wa0=1.55345971674365e-06 pa0=-3.67211856954569e-13
+  keta=-0.257871825644216 lketa=6.21376376523308e-08 wketa=1.33287608886821e-08 pketa=-9.61359436850955e-14
+  a1=0.0
+  a2=0.806834430701738 la2=-1.89988972191417e-09 wa2=5.39557878230444e-07 pa2=-1.49990615453524e-13
+  ags=2.29693798691255 lags=-2.17750538021968e-07 wags=1.4837003852123e-05 pags=-3.08591875719536e-12
+  b0=0.0
+  b1=1.56079073464786e-23 lb1=-4.3388109474329e-30 wb1=-1.09027354236414e-28 pb1=3.03082961494724e-35
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.302375506852193+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff=1.21298736849788e-08 wvoff=1.31742570566053e-06 pvoff=-3.75496168827691e-13
+  nfactor={4.25138870522417+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor=-6.29113696270089e-07 wnfactor=-1.58397267263341e-05 pnfactor=4.43447488731154e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=-4.45493573811138 leta0=9.48170107237301e-07 weta0=2.76205323390022e-05 peta0=-5.64741833500835e-12
+  etab=0.124971191967595 letab=-3.86474083082358e-08 wetab=1.75096264199521e-07 petab=-3.11576779402562e-14
+  dsub=0.917448105477036 ldsub=-1.42368609515037e-07 wdsub=-7.25864735948375e-07 pdsub=2.23726614578682e-13
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=1.9870776373425 lpclm=-2.81622907551503e-07 wpclm=-5.65586271645222e-06 ppclm=1.18119033511035e-12
+  pdiblc1=1.69036691024854 lpdiblc1=-3.14917046285125e-07 wpdiblc1=-3.96577688836422e-06 ppdiblc1=8.39871249452359e-13
+  pdiblc2=0.0625102378327662 lpdiblc2=-1.21565883198577e-08 wpdiblc2=-2.43353657893881e-07 ppdiblc2=5.07773018124314e-14
+  pdiblcb=-0.569956859604857 lpdiblcb=1.02945087315495e-07 wpdiblcb=3.45746778642026e-06 ppdiblcb=-7.19111809961978e-13
+  drout=-4.00933949582378 ldrout=1.05132427420538e-06 wdrout=2.12999060107777e-05 pdrout=-4.56911217797765e-12
+  pscbe1=799950898.804054 lpscbe1=0.0102124595423447 wpscbe1=0.244788719282951 ppscbe1=-5.09131161448989e-8
+  pscbe2=-3.88124220327636e-08 lpscbe2=9.90144747226091e-15 wpscbe2=3.2653436561042e-13 ppscbe2=-6.73234633821834e-20
+  pvag=0.0
+  delta=0.01
+  alpha0=2.83319975417827e-08 lalpha0=-5.8719167047203e-15 walpha0=2.57725595644359e-14 palpha0=-5.36038311868789e-21
+  alpha1=-2.97125714285714e-10 lalpha1=8.25973830628571e-17
+  beta0=35.9652186307162 lbeta0=-5.6790977589156e-06 wbeta0=2.70016386791144e-06 pbeta0=-6.41538342574117e-13
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-3.66793952791247e-09 lagidl=7.93133987247363e-16 wagidl=3.12866726579137e-14 pagidl=-6.55435336506253e-21
+  bgidl=1918143089.39785 lbgidl=-239.253592538879 wbgidl=9187.19470873238 pbgidl=-0.00157349574249591
+  cgidl=-362.589425979443 lcgidl=0.000137810649530612 wcgidl=-0.0018632815287161 pcgidl=3.87540198594604e-10
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=1.08254048749098 lkt1=-4.49995007845275e-07 wkt1=-6.63694748143003e-06 pkt1=1.80094361686878e-12
+  kt2=-0.131083267726 wkt2=6.37296032117115e-8
+  at=612742.466430184 lat=-0.12744072746493 wat=-2.65550289718465 pat=6.07505657055879e-7
+  ute=-1.17383484310212 lute=1.81747161347124e-07 wute=4.35640941088953e-06 pute=-9.06080880552092e-13
+  ua1=-1.9858495788599e-10 lua1=6.93026327807913e-17 wua1=2.32756731381812e-15 pua1=-4.84106070466404e-22
+  ub1=2.37184554712153e-19 lub1=3.23453464345286e-26 wub1=1.08633637849325e-24 pub1=-2.25944930690054e-31
+  uc1=9.50477991212e-11 wuc1=-3.98606031891397e-16
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.1e-6
+  sbref=1.1e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.17 pmos
* DC IV MOS Parameters
+  lmin=1.5e-07 lmax=1.8e-07 wmin=5.0e-06 wmax=7.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.850030758795288+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0=-3.82268882581376e-08 wvth0=-1.03296736801792e-07 pvth0=3.51306053392352e-14
+  k1=-0.724663606244714 lk1=3.56657415097643e-07 wk1=1.17172105464756e-06 pk1=-1.97126743501111e-13
+  k2=0.545043873773805 lk2=-1.49858983617193e-07 wk2=-4.5128980203829e-07 pk2=8.2744930373951e-14
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=332002.835255001 lvsat=-0.0521029411533566 wvsat=-0.384497517541181 pvsat=9.17091435528689e-8
+  ua=-1.1356720783473e-09 lua=-2.39304218232022e-16 wua=1.86599168055105e-15 pua=-3.6943860253356e-22
+  ub=1.4486747753705e-18 lub=1.40441251460858e-25 wub=-5.18047892643157e-24 pub=9.92294566224307e-31
+  uc=-6.91624311790405e-13 luc=1.42757761584407e-19 wuc=6.90994914015749e-18 puc=-1.2042477143751e-24
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.00802035654715585 lu0=-8.10660672925468e-10 wu0=-7.41869197417261e-09 pu0=9.7506230599063e-16
+  a0=1.28721176685324 la0=-1.50858007649149e-07 wa0=-1.67517724574999e-05 pa0=3.440056772502e-12
+  keta=0.326538314613292 lketa=-5.94126585995476e-08 wketa=-3.03575796766507e-06 pketa=5.38037506813342e-13
+  a1=0.0
+  a2=-2.88995283712663 la2=7.66987500539173e-07 wa2=1.61373519873163e-05 pa2=-3.39414461661407e-12
+  ags=1.25
+  b0=0.0
+  b1=-3.64184504751168e-23 lb1=6.48204716316508e-30 wb1=2.54397159884967e-28 pb1=-4.52796416936055e-35
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.4652600366511+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff=4.60079012687937e-08 wvoff=-6.77717186919716e-07 pvoff=3.94696111142877e-14
+  nfactor={-1.71714486913948+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor=6.1226966479466e-07 wnfactor=3.00191839899407e-05 pnfactor=-5.10362823474502e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=-1.89752005415794 leta0=4.16258333963195e-07 weta0=7.61248423470325e-06 peta0=-1.48598442589141e-12
+  etab=-0.272547274226358 letab=4.40316624385122e-08 wetab=-1.41635294846011e-07 petab=3.4718685562506e-14
+  dsub=0.0724235682306968 ldsub=3.33863539377547e-08 wdsub=2.42518199594174e-06 pdsub=-4.31653293093678e-13
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=4.43919083163356 lpclm=-7.91633026605712e-07 wpclm=-1.37119922942032e-05 ppclm=2.85676861372761e-12
+  pdiblc1=1.10627484963891 lpdiblc1=-1.9343290678305e-07 wpdiblc1=5.01235747985451e-07 ppdiblc1=-8.92137747567353e-14
+  pdiblc2=0.0410297202686464 lpdiblc2=-7.6888984327315e-09 wpdiblc2=-1.02300955025996e-07 ppdiblc2=2.14400322483457e-14
+  pdiblcb=-1.5652402037897 lpdiblcb=3.09952079505813e-07 wpdiblcb=7.42943188809961e-06 ppdiblcb=-1.54523267954206e-12
+  drout=1.31472570493286 ldrout=-5.60173987695902e-08 wdrout=-4.63291088693368e-06 pdrout=8.24602542943548e-13
+  pscbe1=1091897231.41031 lpscbe1=-60.7111213665657 wpscbe1=-1455.22218067451 ppscbe1=0.000302668750914132
+  pscbe2=1.20890865910322e-08 lpscbe2=-6.85455503385118e-16 wpscbe2=-1.20887365015751e-14 ppscbe2=3.10607837988624e-21
+  pvag=0.0
+  delta=0.01
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=21.0250054753212 lbeta0=-2.57171270515131e-06 wbeta0=-3.58573617058407e-05 pbeta0=7.37796428645949e-12
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=9.94797529148553e-10 lagidl=-1.76659367776644e-16 wagidl=-5.62065963296656e-15 pagidl=1.12192886345306e-21
+  bgidl=-1559685729.11232 lbgidl=484.093067765413 wbgidl=15980.4271124478 pbgidl=-0.00298640656367986
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-4.18807920411534 lkt1=6.46230640572539e-07 wkt1=1.47989401157595e-05 pkt1=-2.65746377269547e-12
+  kt2=-0.18521100692651 lkt2=1.12579202208355e-08 wkt2=4.41833090426586e-07 pkt2=-7.86409880988472e-14
+  at=-225373.045234974 lat=0.0468772415752826 wat=1.83976401587464 pat=-3.27455917657495e-7
+  ute=-0.3
+  ua1=1.3462e-10
+  ub1=3.927e-19
+  uc1=4.33597582120671e-10 luc1=-7.04142922664941e-17 wuc1=-2.7635090453676e-15 puc1=4.91871447966888e-22
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.04e-6
+  sbref=1.04e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.18 pmos
* DC IV MOS Parameters
+  lmin=2.0e-05 lmax=1.0e-04 wmin=3.0e-06 wmax=5.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.06585217671231+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} wvth0=5.39725375217025e-8
+  k1=0.44180966168701 wk1=-5.60663273386714e-8
+  k2=0.0215768006129515 wk2=-6.63164911639826e-10
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=319843.64933945 wvsat=-0.795325347573929
+  ua=-1.09626656057568e-09 wua=2.69429165360946e-15
+  ub=1.23472887415245e-18 wub=-1.52418976106254e-24
+  uc=-1.04160361652318e-11 wuc=-2.63287684525981e-16
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.00855994754755 wu0=8.9634981324151e-9
+  a0=1.3212184208017 wa0=-6.31775924406513e-7
+  keta=-0.0121258169575241 wketa=3.62151590069734e-8
+  a1=0.0
+  a2=1.07363292255787 wa2=-8.16901592667464e-7
+  ags=0.296043879899246 wags=-3.3968911943596e-7
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.251471733730319+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} wvoff=-3.2386915917047e-9
+  nfactor={1.28816711935094+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} wnfactor=1.36387009947623e-6
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.344479425579197 wpclm=-5.84266556468025e-7
+  pdiblc1=0.39
+  pdiblc2=0.000134084551929727 wpdiblc2=1.72571933786498e-10
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=863994449.244292 wpscbe1=-319.037428105788
+  pscbe2=7.8886136971903e-09 wpscbe2=5.92489086971511e-15
+  pvag=0.0
+  delta=0.01
+  alpha0=2.22675988548041e-10 walpha0=-6.11587916434692e-16
+  alpha1=2.49269515875774e-10 walpha1=-7.4416708014486e-16
+  beta0=1.38266462622756 wbeta0=2.47699175251708e-5
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=2.044997892491e-09 wagidl=-3.32873586518107e-15
+  bgidl=1825806024.97249 wbgidl=-1412.88320678178
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.423714028857974 wkt1=-6.15178011384897e-8
+  kt2=-0.0473577876525128 wkt2=-1.58429699261117e-8
+  at=90000.0
+  ute=-0.154965580668972 wute=-4.85902713039783e-8
+  ua1=1.73469673296457e-09 wua1=1.12001904438913e-15
+  ub1=-7.7325504722252e-19 wub1=1.03835186501631e-25
+  uc1=1.1392027463169e-10 wuc1=-9.91900926583334e-18
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.19 pmos
* DC IV MOS Parameters
+  lmin=8e-06 lmax=2.0e-05 wmin=3.0e-06 wmax=5.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.06585217671231+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} wvth0=5.39725375217025e-8
+  k1=0.44180966168701 wk1=-5.60663273386706e-8
+  k2=0.0215768006129515 wk2=-6.63164911639853e-10
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=319843.64933945 wvsat=-0.795325347573929
+  ua=-1.09626656057568e-09 wua=2.69429165360946e-15
+  ub=1.23472887415245e-18 wub=-1.52418976106254e-24
+  uc=-1.04160361652318e-11 wuc=-2.63287684525981e-16
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.00855994754755 wu0=8.9634981324151e-9
+  a0=1.3212184208017 wa0=-6.31775924406515e-7
+  keta=-0.0121258169575241 wketa=3.62151590069734e-8
+  a1=0.0
+  a2=1.07363292255787 wa2=-8.16901592667464e-7
+  ags=0.296043879899246 wags=-3.3968911943596e-7
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.251471733730319+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} wvoff=-3.23869159170427e-9
+  nfactor={1.28816711935094+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} wnfactor=1.36387009947623e-6
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.344479425579197 wpclm=-5.84266556468025e-7
+  pdiblc1=0.39
+  pdiblc2=0.000134084551929727 wpdiblc2=1.72571933786498e-10
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=863994449.244292 wpscbe1=-319.037428105788
+  pscbe2=7.8886136971903e-09 wpscbe2=5.9248908697151e-15
+  pvag=0.0
+  delta=0.01
+  alpha0=2.22675988548041e-10 walpha0=-6.11587916434693e-16
+  alpha1=2.49269515875774e-10 walpha1=-7.4416708014486e-16
+  beta0=1.38266462622756 wbeta0=2.47699175251708e-5
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=2.044997892491e-09 wagidl=-3.32873586518107e-15
+  bgidl=1825806024.97249 wbgidl=-1412.88320678178
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.423714028857974 wkt1=-6.15178011384897e-8
+  kt2=-0.0473577876525128 wkt2=-1.58429699261117e-8
+  at=90000.0
+  ute=-0.154965580668972 wute=-4.85902713039783e-8
+  ua1=1.73469673296457e-09 wua1=1.12001904438913e-15
+  ub1=-7.7325504722252e-19 wub1=1.03835186501632e-25
+  uc1=1.1392027463169e-10 wuc1=-9.91900926583314e-18
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.20 pmos
* DC IV MOS Parameters
+  lmin=4e-06 lmax=8e-06 wmin=3.0e-06 wmax=5.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.06963048651078+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0=3.0332225722391e-08 wvth0=5.04619428496452e-08 pvth0=2.81830119001467e-14
+  k1=0.52976404061942 lk1=-7.06096698616839e-07 wk1=-4.16088763066334e-07 pk1=2.89025579375245e-12
+  k2=-0.0102118934657894 lk2=2.55199254599803e-07 wk2=1.32459758573231e-07 pk2=-1.06870923226146e-12
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=544267.318869628 lvsat=-1.80167052590423 wvsat=-1.39432209409113 pvsat=4.80873869307915e-6
+  ua=-1.63066796214493e-09 lua=4.29016803898109e-15 wua=4.56788547139998e-15 pua=-1.50411886860965e-20
+  ub=1.54545602020819e-18 lub=-2.49451379980975e-24 wub=-2.613424091441e-24 pub=8.74436013346629e-30
+  uc=4.582367216758e-12 luc=-1.20407002369773e-16 wuc=-3.48263192133005e-16 puc=6.82182355363101e-22
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.00629440413992117 lu0=1.81877552899234e-08 wu0=1.65029548736302e-08 pu0=-6.0526668244994e-14
+  a0=1.33793090277023 la0=-1.34167604693537e-07 wa0=-6.3243537395748e-07 pa0=5.29405308173668e-15
+  keta=-0.0126902903205591 lketa=4.53158538476451e-09 wketa=6.70453453845611e-08 pketa=-2.47504366277037e-13
+  a1=0.0
+  a2=1.34918045467487 la2=-2.21209228126493e-06 wa2=-1.63951904577882e-06 pa2=6.60396304216854e-12
+  ags=0.334419598534634 lags=-3.08079808696275e-07 wags=-9.52571265673284e-07 pags=4.92021051540748e-12
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.253832649645215+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff=1.89534046337942e-08 wvoff=9.25432572850707e-10 pvoff=-3.34295388235551e-14
+  nfactor={1.22318305266557+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor=5.21691307541333e-07 wnfactor=1.72703795968711e-06 pnfactor=-2.91550722375856e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.206725750144198 lpclm=1.10588485334806e-06 wpclm=-9.6651049368957e-07 ppclm=3.06864974108731e-12
+  pdiblc1=0.39
+  pdiblc2=0.000322442719140064 lpdiblc2=-1.51213710606658e-09 wpdiblc2=-4.5922622307049e-10 ppdiblc2=5.07206802167003e-15
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=928436667.649947 lpscbe1=-517.341356053972 wpscbe1=-640.307161096034 ppscbe1=0.0025791495612089
+  pscbe2=6.36982365594844e-09 lpscbe2=1.21928282256092e-14 wpscbe2=1.15473719793668e-14 ppscbe2=-4.51372108785108e-20
+  pvag=0.0
+  delta=0.01
+  alpha0=2.1778265896932e-10 lalpha0=3.92835911380165e-17 walpha0=-5.87192749320908e-16 palpha0=-1.95844108847456e-22
+  alpha1=2.50600308015112e-10 lalpha1=-1.06835833250958e-17 walpha1=-7.50801600896135e-16 palpha1=5.3261852976983e-23
+  beta0=-9.4582837194124 lbeta0=8.70310032274175e-05 wbeta0=7.72154682075711e-05 pbeta0=-4.21032251531701e-10
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=1.96968488748295e-09 lagidl=6.04611900448605e-16 wagidl=-4.48505197082119e-16 pagidl=-2.31224572407303e-20
+  bgidl=1435872467.17634 lbgidl=3130.38192278479 wbgidl=811.057198262406 pbgidl=-0.0178537668844098
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.36925500460282 lkt1=-4.37196393212085e-07 wkt1=-1.98403491304958e-07 pkt1=1.09891667802813e-12
+  kt2=-0.0432594978210332 lkt2=-3.290102158764e-08 wkt2=-3.17967931127962e-08 pkt2=1.28077101096826e-13
+  at=13497.2871138284 lat=0.614162861017631 wat=0.359699755072383 pat=-2.88766531732403e-6
+  ute=-0.0288287594987497 lute=-1.01262488671269e-06 wute=-4.72207773603336e-07 pute=3.40079622504922e-12
+  ua1=1.28492568479749e-09 lua1=3.61075657743271e-15 wua1=2.24787486203185e-15 pua1=-9.05441296976595e-21
+  ub1=-6.22270435662136e-19 lub1=-1.21210264979143e-24 wub1=2.08396907803213e-25 pub1=-8.3942024386845e-31
+  uc1=3.59891340229908e-10 luc1=-1.97465276296971e-15 wuc1=-1.99074218394996e-17 puc1=8.0186856280442e-23
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.21 pmos
* DC IV MOS Parameters
+  lmin=2e-06 lmax=4e-06 wmin=3.0e-06 wmax=5.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.07224101358323+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0=4.08473974438931e-08 wvth0=6.4767690430209e-08 pvth0=-2.9440367685387e-14
+  k1=0.37366012860566 lk1=-7.73120142723565e-08 wk1=6.93074070362553e-08 pk1=9.35085845333262e-13
+  k2=0.0449017933247142 lk2=3.32019855718958e-08 wk2=-4.3678778043131e-08 pk2=-3.59225320433194e-13
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=97503.5788322117 lvsat=-0.00211154219840071 wvsat=-0.186289436856035 pvsat=-5.72023538719362e-8
+  ua=1.3507363128952e-10 lua=-2.82221791047376e-15 wua=3.06336452805816e-16 pua=2.1242796222126e-21
+  ub=4.63252491038355e-19 lub=1.86458902924401e-24 wub=1.17241258538553e-25 pub=-2.25472712826714e-30
+  uc=-6.16313473490057e-11 luc=1.46301045336548e-16 wuc=-1.33215754592883e-16 puc=-1.84026142479259e-22
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0136568945468041 lu0=-1.14682677191161e-08 wu0=-1.91519764212138e-11 pu0=6.02417988173103e-15
+  a0=1.1172682009854 la0=7.54659110143325e-07 wa0=4.20373074220957e-07 pa0=-4.23540574247959e-12
+  keta=-0.0139430117354255 lketa=9.57753221118941e-09 wketa=4.93170614460544e-08 pketa=-1.76095051312139e-13
+  a1=0.0
+  a2=0.8
+  ags=0.254098822546019 lags=1.54513131365553e-08 wags=-4.67064092148974e-07 pags=2.96459344653765e-12
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.245204931884238+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff=-1.57989389748084e-08 wvoff=-4.33580592351117e-08 pvoff=1.44943834777012e-13
+  nfactor={1.67455573885579+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.29643245596062e-06 wnfactor=3.73375794083068e-07 pnfactor=2.53702773534853e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.280942516865585 leta0=-8.09394046624373e-07 weta0=-5.99892222498885e-07 peta0=2.41635867351884e-12
+  etab=-0.245666731739443 letab=7.07583487445697e-07 wetab=5.24434090734426e-07 petab=-2.11241422426918e-12
+  dsub=1.31827366676702 ldsub=-3.05431723045356e-06 wdsub=-2.26374429023166e-06 pdsub=9.11833483612165e-12
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-0.0167107524854462 lpclm=2.00588440470224e-06 wpclm=1.2727277044652e-06 ppclm=-5.9509748502217e-12
+  pdiblc1=0.39
+  pdiblc2=-0.000868109022524547 lpdiblc2=3.28339102273757e-09 wpdiblc2=3.23350522759441e-09 ppdiblc2=-9.80220994883077e-15
+  pdiblcb=0.0108149534565344 lpdiblcb=-1.44262202743479e-07 wpdiblcb=-1.7855158960557e-07 ppdiblcb=7.1920366031216e-13
+  drout=0.56
+  pscbe1=829191134.970585 lpscbe1=-117.581541367899 wpscbe1=-87.1469866503321 ppscbe1=0.000351027016463702
+  pscbe2=8.69970203313866e-09 lpscbe2=2.80810608082749e-15 wpscbe2=3.86962274321286e-15 ppscbe2=-1.42113290882733e-20
+  pvag=0.0
+  delta=0.01
+  alpha0=2.81831355015394e-10 lalpha0=-2.18703787951219e-16 walpha0=-9.06500619009178e-16 palpha0=1.09032415856246e-21
+  alpha1=3.97966325078039e-10 lalpha1=-6.04272131662362e-16 walpha1=-1.48547899290672e-15 palpha1=3.01253357186691e-21
+  beta0=13.5215377181067 lbeta0=-5.53144176505219e-06 wbeta0=-4.20567771028238e-05 pbeta0=5.93949213116258e-11
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=3.77980778446279e-09 lagidl=-6.68654140711146e-15 wagidl=-1.11228910436927e-14 pagidl=1.98738408567869e-20
+  bgidl=2570451567.50282 lbgidl=-1439.68907838105 wbgidl=-4688.41386010068 pbgidl=0.00429803654502397
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.50460799020204 lkt1=1.08003808545747e-07 wkt1=2.20343295790019e-07 pkt1=-5.87790355428998e-13
+  kt2=-0.0754041176538033 lkt2=9.65771213633199e-08 wkt2=8.60291949947027e-08 pkt2=-3.46524565088322e-13
+  at=174420.68008278 lat=-0.0340346347805908 wat=-0.324619589651941 pat=-1.31235208606589e-7
+  ute=-1.40423704832166 lute=4.52750319576653e-06 wute=6.42644637334934e-06 pute=-2.43868998950264e-11
+  ua1=3.36989280642313e-10 lua1=7.42903303813294e-15 wua1=1.26418007577486e-14 pua1=-5.09210217506021e-20
+  ub1=4.58142767663473e-19 lub1=-5.56399406782854e-24 wub1=-8.77924729609942e-24 pub1=3.53627027577209e-29
+  uc1=-5.35545681927539e-10 luc1=1.63215681703623e-15 wuc1=7.8454291579801e-16 puc1=-3.16012945031939e-21
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.22 pmos
* DC IV MOS Parameters
+  lmin=1e-06 lmax=2e-06 wmin=3.0e-06 wmax=5.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.05431745609063+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0=4.49863793159452e-09 wvth0=-8.01673989473574e-09 pvth0=1.18165583600433e-13
+  k1=0.0980653419667101 lk1=4.81590905893993e-07 wk1=1.33884739921875e-06 pk1=-1.63952602433292e-12
+  k2=0.154627916744053 lk2=-1.89321276009043e-07 wk2=-5.43376155013411e-07 pk2=6.54154963694011e-13
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=244870.871758392 lvsat=-0.300970643845179 wvsat=-0.823819744891491 pvsat=1.23570146046027e-6
+  ua=-1.72978311402204e-09 lua=9.59689190737141e-16 wua=4.46701970012618e-15 pua=-6.31353607515413e-21
+  ub=1.68939709549884e-18 lub=-6.22017514866594e-25 wub=-2.89482804724683e-24 pub=3.85371327903394e-30
+  uc=5.25843552313134e-11 luc=-8.5327028907908e-17 wuc=-4.55175768638106e-16 puc=4.68904902484284e-22
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.00611174655753136 lu0=3.8332018613531e-09 wu0=1.57933447826701e-08 pu0=-2.60433737957449e-14
+  a0=2.85342139564645 la0=-2.76623873479096e-06 wa0=-6.1136979532685e-06 pa0=9.01561189241668e-12
+  keta=0.102921143491894 lketa=-2.27421572219952e-07 wketa=-4.14883587189008e-07 pketa=7.65298293711983e-13
+  a1=0.0
+  a2=0.8
+  ags=-1.46540800495429 lags=3.50259052522526e-06 wags=6.0091333255244e-06 pags=-1.01690572021349e-11
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.306431699428405+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff=1.08368210883552e-07 wvoff=2.11938689795257e-07 pvoff=-3.72794908695587e-13
+  nfactor={-0.352535582831902+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor=2.81448441932616e-06 wnfactor=6.47398133412741e-06 pnfactor=-9.83492709259492e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=-0.743360113731169 leta0=1.26787939659428e-06 weta0=1.19978444499777e-06 peta0=-1.23336401204437e-12
+  etab=-34.7328784543308 letab=7.06472350143202e-05 wetab=0.000173158372662235 petab=-3.52211970040009e-10
+  dsub=-0.648150933534041 ldsub=9.33568261861792e-07 wdsub=4.52748858046332e-06 pdsub=-4.65420393085333e-12
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=1.85601505614594 lpclm=-1.79198106249251e-06 wpclm=-4.94789853553843e-06 ppclm=6.66438051699077e-12
+  pdiblc1=0.391067255322459 lpdiblc1=-2.16438098688287e-09 wpdiblc1=3.94686325668098e-08 ppdiblc1=-8.00419132218985e-14
+  pdiblc2=0.00108084150236606 lpdiblc2=-6.69057254334284e-10 wpdiblc2=-3.24470014933205e-09 ppdiblc2=3.33551281711155e-15
+  pdiblcb=-0.121567847713041 lpdiblcb=1.24208529434806e-07 wpdiblcb=3.57213897670962e-07 ppdiblcb=-3.673223186988e-13
+  drout=0.220528215552783 ldrout=6.88444705197542e-07 wdrout=4.0147504705487e-07 pdrout=-8.14186577726708e-13
+  pscbe1=741617730.058828 lpscbe1=60.0162729122849 wpscbe1=174.293973300666 ppscbe1=-0.000179172113025405
+  pscbe2=1.32811339333389e-08 lpscbe2=-6.48298283559588e-15 wpscbe2=-7.56924108632876e-15 ppscbe2=8.98654949167113e-21
+  pvag=0.0
+  delta=0.01
+  alpha0=2.50048018043741e-10 lalpha0=-1.54247561972749e-16 walpha0=-7.48048218780726e-16 palpha0=7.68984592327961e-22
+  alpha1=1.0e-10
+  beta0=12.6274591926958 lbeta0=-3.71826124446125e-06 wbeta0=-2.54864799051063e-05 pbeta0=2.5790557438221e-11
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=1.09713481351658e-09 lagidl=-1.2461128141082e-15 wagidl=-3.85491552309459e-15 pagidl=5.13447371672018e-21
+  bgidl=2579670906.36265 lbgidl=-1458.38578695672 wbgidl=-5324.88602313467 pbgidl=0.00558879445399096
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.390580576897025 lkt1=-1.23242417307863e-07 wkt1=-3.27766933962736e-07 pkt1=5.23770613186833e-13
+  kt2=-0.0111038593327429 lkt2=-3.38230309086907e-08 wkt2=-1.53064749815835e-07 pkt2=1.3835508586011e-13
+  at=353983.792411005 lat=-0.398186471824883 wat=-1.09079131010945 pat=1.4225518464206e-6
+  ute=1.67023776830381 lute=-1.70749483865212e-06 wute=-1.00772125235107e-05 pute=9.08232230389904e-12
+  ua1=3.61852389490631e-09 lua1=7.7412021882092e-16 wua1=-1.26413861642257e-14 pua1=3.52977928918536e-22
+  ub1=-6.77880942391506e-19 lub1=-3.26015161612156e-24 wub1=4.17238556081607e-24 pub1=9.09694674349057e-30
+  uc1=7.19692533299023e-10 luc1=-9.13451220584661e-16 wuc1=-2.37729025009802e-15 puc1=3.25203026811976e-21
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=2.745e-6
+  sbref=2.74e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.23 pmos
* DC IV MOS Parameters
+  lmin=5e-07 lmax=1e-06 wmin=3.0e-06 wmax=5.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.09311938443813+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0=4.43865546496828e-08 wvth0=1.6011460155065e-07 pvth0=-5.4671417829325e-14
+  k1=0.607856353255918 lk1=-4.2468136219177e-08 wk1=-2.84503246138047e-07 pk1=2.92589588861162e-14
+  k2=-0.0503231996028657 lk2=2.13660121821936e-08 wk2=1.07215571730609e-07 pk2=-1.46455242981209e-14
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=-171328.91580929 lvsat=0.126877743376947 wvsat=0.712232669634504 pvsat=-3.43341989043476e-7
+  ua=3.94608610900403e-11 lua=-8.59072384750374e-16 wua=-4.63051749550091e-15 pua=3.03862299150418e-21
+  ub=6.11580293647775e-19 lub=4.85965223634673e-25 wub=2.54781093588378e-24 pub=-1.74125428395653e-30
+  uc=-4.25031695544227e-11 luc=1.24218055215313e-17 wuc=-3.52826814783031e-17 puc=3.72598476010526e-23
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0134637613764527 lu0=-3.72458114832024e-09 wu0=-2.16872036298233e-08 pu0=1.24861802057172e-14
+  a0=-0.456732722382784 la0=6.36559976693679e-07 wa0=4.65393856812308e-06 pa0=-2.0533892399356e-12
+  keta=-0.226023486691235 lketa=1.10729560272743e-07 wketa=6.65289102850801e-07 pketa=-3.4510626957666e-13
+  a1=0.0
+  a2=0.858265210704412 la2=-5.98959374216073e-08 wa2=-3.03802735891509e-07 pa2=3.1230556686364e-13
+  ags=3.23940229355105 lags=-1.33389800391465e-06 wags=-8.8962954943298e-06 pags=5.15354475952933e-12
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.187819540799715+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff=-1.35636648408379e-08 wvoff=-1.76261707236047e-07 pvoff=2.62704410478296e-14
+  nfactor={2.93720749969435+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor=-5.67331992593843e-07 wnfactor=-5.27738863376058e-06 pnfactor=2.24534021795432e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.49
+  etab=69.8838533918854 letab=-3.68975099228079e-05 wetab=-0.000348411066080627 petab=1.83955154154389e-10
+  dsub=0.222046819523638 ldsub=3.9015414091535e-08 wdsub=2.08522867129654e-08 pdsub=-2.14359005134877e-14
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-0.428421300191785 lpclm=5.56392098586396e-07 wpclm=3.16398490696842e-06 ppclm=-1.67453831930497e-12
+  pdiblc1=1.04647985794606 lpdiblc1=-6.75920671532716e-07 wpdiblc1=-1.41190780375686e-06 ppdiblc1=1.4119556468016e-12
+  pdiblc2=0.000678123889252548 lpdiblc2=-2.55068380664949e-10 wpdiblc2=-1.23699490211332e-09 ppdiblc2=1.27161591543367e-15
+  pdiblcb=0.236071081599945 lpdiblcb=-2.43439998231792e-07 wpdiblcb=-2.21436919645206e-10 ppdiblcb=1.16916036329595e-16
+  drout=0.774314128894433 ldrout=1.19159431713286e-07 wdrout=-8.02950094109737e-07 pdrout=4.23948014288812e-13
+  pscbe1=800000000.0
+  pscbe2=2.64032820157266e-08 lpscbe2=-1.99723935985134e-14 wpscbe2=-6.29950868783798e-14 ppscbe2=6.59636538557501e-20
+  pvag=0.0
+  delta=0.01
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=8.54089891363691 lbeta0=4.82673683687974e-07 wbeta0=-6.01300567961907e-07 pbeta0=2.08891701788605e-13
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-5.38320026446754e-10 lagidl=4.35115135916034e-16 wagidl=3.10841891577484e-15 pagidl=-2.02375052642433e-21
+  bgidl=753521141.376451 lbgidl=418.874257651909 wbgidl=1953.73370342503 pbgidl=-0.00189353928147571
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.512587569822165 lkt1=2.17930733526492e-09 wkt1=3.73660276552699e-07 pkt1=-1.97288142096507e-13
+  kt2=-0.0321981266248769 lkt2=-1.21383772635845e-08 wkt2=-3.79872803471408e-08 pkt2=2.00568281759261e-14
+  at=-138709.587173076 lat=0.108296410066998 wat=0.578888246083538 pat=-2.93858701191119e-7
+  ute=0.354388745501949 lute=-3.54817833400083e-07 wute=-2.5538624874394e-06 pute=1.34840874701815e-12
+  ua1=8.69330327009257e-09 lua1=-4.44269208151806e-15 wua1=-2.61585802879867e-14 pua1=1.42484912818154e-20
+  ub1=-8.43319901854543e-18 lub1=4.71222230234777e-24 wub1=2.70064719205692e-23 pub1=-1.43762200252993e-29
+  uc1=-3.72913201647328e-10 luc1=2.0973436367137e-16 wuc1=1.616408837004e-15 puc1=-8.53444469032066e-22
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.745e-6
+  sbref=1.74e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.24 pmos
* DC IV MOS Parameters
+  lmin=2.5e-07 lmax=5e-07 wmin=3.0e-06 wmax=5.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.69237414749775+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0=-1.67202121511997e-07 wvth0=-1.53846743104571e-06 pvth0=8.42159512397162e-13
+  k1=0.111235728789203 lk1=2.19741594051755e-07 wk1=-4.91382524751791e-08 pk1=-9.50109333879541e-14
+  k2=0.127938719360873 lk2=-7.27541418876327e-08 wk2=2.34374096309928e-08 pk2=2.95883399525312e-14
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=8143.60268097318 lvsat=0.0321184072843101 wvsat=0.350134942055627 pvsat=-1.5215873405456e-7
+  ua=-9.35894198245189e-10 lua=-3.44096617682085e-16 wua=1.66949866501979e-15 pua=-2.87709941056827e-22
+  ub=1.02366082295916e-18 lub=2.68391649124614e-25 wub=-9.77010244914083e-25 pub=1.19809001650575e-31
+  uc=-5.10855973052019e-11 luc=1.69532243848097e-17 wuc=1.28744603233091e-16 puc=-4.93445903991469e-23
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.00709506696259313 lu0=-3.61986922135346e-10 wu0=1.2300002722226e-08 pu0=-5.45865690168857e-15
+  a0=0.559400242467097 la0=1.0005396484852e-07 wa0=3.00430417121536e-06 pa0=-1.18240207398109e-12
+  keta=0.117680960981484 lketa=-7.07422636450811e-08 wketa=-1.7359409610752e-07 pketa=9.78139928749459e-14
+  a1=0.0
+  a2=0.683469578591175 la2=3.23940587865962e-08 wa2=6.07605471783016e-07 pa2=-1.68907029890017e-13
+  ags=-3.26526362487771 lags=2.10048754502471e-06 wags=1.30664148922167e-05 pags=-6.44250277204261e-12
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.205339729331252+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff=-4.31321553844871e-09 wvoff=-2.00855033485626e-08 pvoff=-5.61887204903156e-14
+  nfactor={1.38500884853079+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor=2.52210268836702e-07 wnfactor=-6.03956829010318e-07 pnfactor=-2.22175693772163e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.353485933730394 leta0=7.20777888215568e-08 weta0=1.0618783737044e-06 peta0=-5.60659038775439e-13
+  etab=0.00514231527341621 letab=-2.38901888966769e-09 wetab=-1.81233701833225e-08 petab=7.86111858654968e-15
+  dsub=0.290725058975033 ldsub=2.75412780007136e-09 wdsub=-7.09758990772381e-07 pdsub=3.64318086663445e-13
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.812502089886035 lpclm=-9.88005602940122e-08 wpclm=-1.31719740270458e-06 ppclm=6.91472166014662e-13
+  pdiblc1=-0.87109547305574 lpdiblc1=3.36536092332264e-07 wpdiblc1=2.50769738067592e-06 ppdiblc1=-6.57548855316698e-13
+  pdiblc2=-0.00500165762792038 lpdiblc2=2.74378810302415e-09 wpdiblc2=-7.15407780804622e-09 ppdiblc2=4.39576468477137e-15
+  pdiblcb=-0.612965135720228 lpdiblcb=2.04840936078652e-07 wpdiblcb=8.25454995976688e-07 ppdiblcb=-4.3583033241574e-13
+  drout=1.01083301632419 ldrout=-5.71970262297527e-09 wdrout=1.34227123328469e-06 pdrout=-7.0870310391952e-13
+  pscbe1=800000000.0
+  pscbe2=-4.68577695333453e-08 lpscbe2=1.8708562486778e-14 wpscbe2=1.68043499057875e-13 ppscbe2=-5.6021947055561e-20
+  pvag=0.0
+  delta=0.01
+  alpha0=-2.32128195859522e-08 lalpha0=1.23088889875477e-14 walpha0=6.95979097519089e-14 palpha0=-3.67468611740909e-20
+  alpha1=3.7717584137872e-10 lalpha1=-1.46345518137868e-16 walpha1=-8.27478594880468e-16 palpha1=4.36898768353749e-22
+  beta0=-8.50151007830923 lbeta0=9.48086112252763e-06 wbeta0=5.49406538008938e-05 pbeta0=-2.91165937015148e-11
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=2.8304705487095e-09 lagidl=-1.34356586227957e-15 wagidl=-1.66871367768091e-14 pagidl=8.42806533259166e-21
+  bgidl=34752386.8210707 lbgidl=798.375534832095 wbgidl=2881.642695453 pbgidl=-0.00238346409435857
+  cgidl=626.255574195907 lcgidl=-0.000172259028108549 wcgidl=-0.000179878083059782 pcgidl=9.49734693185679e-11
+  egidl=2.20111972662033 legidl=-1.10936600221882e-06 wegidl=-1.04749058963591e-05 pegidl=5.53062461440687e-12
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.386136323069855 lkt1=-6.45854335349934e-08 wkt1=-2.79770512929085e-07 pkt1=1.47715473580402e-13
+  kt2=0.11033875387042 lkt2=-8.73961397225351e-08 wkt2=-4.75353353615034e-07 pkt2=2.50980866468495e-13
+  at=67228.2041039711 lat=-0.000436272473787899 wat=0.0785190978600638 pat=-2.9669795358903e-8
+  ute=-0.33723371376 lute=1.03505256207149e-8
+  ua1=4.57804105070251e-10 lua1=-9.44473483762536e-17 wua1=1.46985262371035e-15 pua1=-3.38989754365674e-22
+  ub1=5.581698006954e-19 lub1=-3.51125377855634e-26 wub1=-3.38510828351616e-25 pub1=6.16027263378787e-32
+  uc1=1.05251536618683e-11 luc1=7.28351332837748e-18 wuc1=1.19922749102349e-16 puc1=-6.33177724530512e-23
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.245e-6
+  sbref=1.24e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.25 pmos
* DC IV MOS Parameters
+  lmin=1.8e-07 lmax=2.5e-07 wmin=3.0e-06 wmax=5.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-2.05698104162996+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0=2.12142219774028e-07 wvth0=5.67910341297341e-06 pvth0=-1.16423857139003e-12
+  k1=0.517108815050108 lk1=1.06913746548259e-07 wk1=-1.61031557114145e-06 pk1=3.38977627073446e-13
+  k2=0.00989741452749859 lk2=-3.99400756396127e-08 wk2=5.75945091001007e-07 pk2=-1.24002165376156e-13
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=234047.757030305 lvsat=-0.0306802367749521 wvsat=-0.876184352313243 pvsat=1.88743313948454e-7
+  ua=-1.7683141663095e-09 lua=-1.12693855599822e-16 wua=1.89914290081789e-15 pua=-3.51548282877873e-22
+  ub=1.86129873909603e-18 lub=3.55383600935579e-26 wub=-2.31052546704758e-24 pub=4.90510231221019e-31
+  uc=3.88090964234418e-11 luc=-8.03642173542856e-18 wuc=-1.94373221697998e-16 puc=4.04782875177967e-23
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0122696634293582 lu0=-1.80046264473842e-09 wu0=-2.85700631384478e-08 pu0=5.90273096678843e-15
+  a0=3.75554605911061 la0=-7.88436218428578e-07 wa0=-1.31755424740778e-05 pa0=3.31540113525067e-12
+  keta=-0.073204668515808 lketa=-1.76783492723879e-08 wketa=-9.07309443855457e-07 pketa=3.01778054964699e-13
+  a1=0.0
+  a2=0.518565270761412 la2=7.82354775115763e-08 wa2=1.97669269969749e-06 pa2=-5.49496850203505e-13
+  ags=13.3256920067458 lags=-2.51159902909904e-06 wags=-4.01456604140722e-05 pags=8.34981561820205e-12
+  b0=0.0
+  b1=-1.56079073464786e-23 lb1=4.3388109474329e-30 wb1=4.65957248504999e-29 pb1=-1.29530523597408e-35
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={0.305855280067916+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff=-1.46419293811305e-07 wvoff=-1.71484331525084e-06 pvoff=4.14933614124775e-13
+  nfactor={1.16590864714949+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor=3.13117495618288e-07 wnfactor=-4.57398511553034e-07 pnfactor=-2.62917147325478e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=1.77650939199273 leta0=-3.23505656293872e-07 weta0=-3.44566560734673e-06 peta0=6.92384097429002e-13
+  etab=0.0518455394210459 letab=-1.53719547640189e-08 wetab=5.39656322024998e-07 petab=-1.47194942491057e-13
+  dsub=0.153984768260277 ldsub=4.07662877352853e-08 wdsub=3.08029943039803e-06 pdsub=-6.89272673720874e-13
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-0.109830324704986 lpclm=1.57596782973317e-07 wpclm=4.7980458816572e-06 ppclm=-1.0084920841185e-12
+  pdiblc1=0.737367328973287 lpdiblc1=-1.10597265078181e-07 wpdiblc1=7.85299790728681e-07 ppdiblc1=-1.78742994082445e-13
+  pdiblc2=0.00594861771443089 lpdiblc2=-3.00257038845393e-10 wpdiblc2=3.86282018634308e-08 ppdiblc2=-8.33115967654318e-15
+  pdiblcb=1.04668204256623 lpdiblcb=-2.56521063718845e-07 wpdiblcb=-4.60211118668005e-06 ppdiblcb=1.07296793556864e-12
+  drout=1.61785633007545 ldrout=-1.7446489956606e-07 wdrout=-6.75387216753285e-06 pdrout=1.54192760778695e-12
+  pscbe1=800000000.0
+  pscbe2=5.38579888049033e-08 lpscbe2=-9.28920974215507e-15 wpscbe2=-1.3546397775048e-13 ppscbe2=2.83494894074398e-20
+  pvag=0.0
+  delta=0.01
+  alpha0=8.33600699498292e-08 lalpha0=-1.73170954287251e-14 walpha0=-2.48563963399674e-13 palpha0=5.16983216195715e-20
+  alpha1=-8.89913719209714e-10 lalpha1=2.0589017463099e-16 walpha1=2.95528069600167e-15 palpha1=-6.14662921399995e-22
+  beta0=76.1650183581019 lbeta0=-1.40554177844534e-05 wbeta0=-0.000197711604134559 pbeta0=4.11177021774459e-11
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-7.35639591473438e-09 lagidl=1.48826077216027e-15 wagidl=4.96750743588158e-14 pagidl=-1.00198330165784e-20
+  bgidl=7882249052.55016 lbgidl=-1383.13436828061 wbgidl=-20546.2126399406 pbgidl=0.00412919855461685
+  cgidl=-865.198479271098 lcgidl=0.000242347301306637 wcgidl=0.000642421725213504 pcgidl=-1.33616009783706e-10
+  egidl=-7.40399902364405 legidl=1.56074174892968e-06 wegidl=3.74103782012826e-05 pegidl=-7.78090974132838e-12
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-1.00994470300671 lkt1=1.08825810386893e-07 wkt1=3.79491186589264e-06 pkt1=-9.84997331543492e-13
+  kt2=-0.475065770562859 lkt2=7.53392932156233e-08 wkt2=1.77861728979107e-06 pkt2=-3.75595924750681e-13
+  at=169427.559955075 lat=-0.0288464670081245 wat=-0.445404220299908 pat=1.15974600009751e-7
+  ute=-0.3
+  ua1=6.88193517716455e-11 lua1=1.36857452237189e-17 wua1=9.94451954204561e-16 pua1=-2.06834073051098e-22
+  ub1=5.48215445287846e-19 lub1=-3.23453464345286e-26 wub1=-4.64274597341862e-25 pub1=9.65635449519396e-32
+  uc1=3.6725972864055e-11 wuc1=-1.07848854179271e-16
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.1e-6
+  sbref=1.1e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.26 pmos
* DC IV MOS Parameters
+  lmin=1.5e-07 lmax=1.8e-07 wmin=3.0e-06 wmax=5.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.960264026003735+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0=-1.59617588720394e-08 wvth0=4.46259333719737e-07 pvth0=-7.58697970342118e-14
+  k1=-0.296887372665633 lk1=2.7621518563888e-07 wk1=-9.60911243582975e-07 pk1=2.03909319793214e-13
+  k2=0.396688359746296 lk2=-1.2038795075378e-07 wk2=2.88320620421442e-07 pk2=-6.41797269892537e-14
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=120859.556181338 lvsat=-0.00713844925677692 wvsat=0.668134539035084 pvsat=-1.32456483625302e-7
+  ua=-6.94613071502795e-10 lua=-3.36010798906481e-16 wua=-3.3286045191125e-16 pua=1.12681630449556e-22
+  ub=1.25646898917168e-19 lub=3.96533115028679e-25 wub=1.41533392922136e-24 pub=-2.84423812890165e-31
+  uc=8.64214249584742e-13 luc=-1.44341581852367e-19 wuc=-8.46516288181396e-19 puc=2.2705511301971e-25
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.00674518297616 lu0=-6.51437004238645e-10 wu0=-1.06145159968366e-09 pu0=1.8126987006396e-16
+  a0=-6.86077712125912 la0=1.41963160721016e-06 wa0=2.38691477909821e-05 pa0=-4.38944990359861e-12
+  keta=-0.825048860183211 lketa=1.38696220464132e-07 wketa=2.70535575118545e-06 pketa=-4.49612953621469e-13
+  a1=0.0
+  a2=2.76344646704595 la2=-3.88672872741253e-07 wa2=-1.20470608071911e-05 pa2=2.36727559418725e-12
+  ags=1.25
+  b0=0.0
+  b1=3.64184504751168e-23 lb1=-6.48204716316509e-30 wb1=-1.087233579845e-28 pb1=1.93514530409452e-35
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.764685300034826+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff=7.62403003631043e-08 wvoff=8.15035185636466e-07 pvoff=-1.11250755517775e-13
+  nfactor={4.53005986986764+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor=-3.86585588892415e-07 wnfactor=-1.12558178770849e-06 pnfactor=-1.23943044084458e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.121958650053124 leta0=2.06210434206614e-08 weta0=-2.45540914533672e-06 peta0=4.86422636408465e-13
+  etab=-0.0623581802556036 letab=8.381048484088e-09 wetab=-1.18951036445288e-06 petab=2.12450978296104e-13
+  dsub=0.883879723873455 ldsub=-1.11043104292788e-07 wdsub=-1.62024519304165e-06 pdsub=2.88384201419098e-13
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=1.60732549945199 lpclm=-1.99551022581445e-07 wpclm=4.05967044305216e-07 ppclm=-9.49923908953373e-14
+  pdiblc1=1.30985000315984 lpdiblc1=-2.29666791516893e-07 wpdiblc1=-5.13666234491565e-07 ppdiblc1=9.14263515710638e-14
+  pdiblc2=0.0132604600262662 lpdiblc2=-1.8210324975994e-09 wpdiblc2=3.61396983861358e-08 ppdiblc2=-7.81358081530755e-15
+  pdiblcb=-0.185381051168264 lpdiblcb=-2.66724979194323e-10 wpdiblcb=5.50292831522065e-07 ppdiblcb=1.32972863082054e-15
+  drout=-0.53193990621094 ldrout=2.72666920026673e-07 wdrout=4.57344144687087e-06 pdrout=-8.14017696245653e-13
+  pscbe1=800000000.0
+  pscbe2=1.06672940621216e-08 lpscbe2=-3.06063523993387e-16 wpscbe2=-5.00054311792556e-15 ppscbe2=1.21466056508415e-21
+  pvag=0.0
+  delta=0.01
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=11.0593811976463 lbeta0=-5.14226522724595e-07 wbeta0=1.38251838362102e-05 pbeta0=-2.87941127901845e-12
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-1.04627209499632e-09 lagidl=1.75830739140593e-16 wagidl=4.55487295090224e-15 pagidl=-6.35372566149298e-22
+  bgidl=2609694922.03997 lbgidl=-286.50637978405 wbgidl=-4805.57066463772 pbgidl=0.000855333911457538
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=0.120672169813581 lkt1=-1.26328931757253e-07 wkt1=-6.68187537556506e-06 pkt1=1.19404869323281e-12
+  kt2=-0.0587089930734905 lkt2=-1.12579202208356e-08 wkt2=-1.88829062720548e-07 pkt2=3.36093072155047e-14
+  at=-12370.3889396135 lat=0.00896532478658391 wat=0.777862234600464 pat=-1.38450143412067e-7
+  ute=-0.3
+  ua1=1.3462e-10
+  ub1=3.927e-19
+  uc1=2.92562488016356e-11 luc1=1.55361296829446e-18 wuc1=-7.47708916101277e-16 puc1=1.33083214559034e-22
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.04e-6
+  sbref=1.04e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.27 pmos
* DC IV MOS Parameters
+  lmin=2.0e-05 lmax=1.0e-04 wmin=2e-06 wmax=3.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.0477733+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+  k1=0.42302944
+  k2=0.021354664
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=53438.0
+  ua=-1.9377487e-10
+  ub=7.2417962e-19
+  uc=-9.8608028e-11
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0115624
+  a0=1.109596
+  keta=4.9707517e-6
+  a1=0.0
+  a2=0.8
+  ags=0.18226013
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.25255658+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.745015+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.14877095
+  pdiblc1=0.39
+  pdiblc2=0.00019189
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=757128280.0
+  pscbe2=9.873241e-9
+  pvag=0.0
+  delta=0.01
+  alpha0=1.7815831e-11
+  alpha1=6.3056523e-17
+  beta0=9.6797043
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=9.2999e-10
+  bgidl=1352540500.0
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.4443203
+  kt2=-0.052664618
+  at=90000.0
+  ute=-0.17124159
+  ua1=2.1098632e-9
+  ub1=-7.3847396e-19
+  uc1=1.1059776e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.28 pmos
* DC IV MOS Parameters
+  lmin=8e-06 lmax=2.0e-05 wmin=2e-06 wmax=3.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.0477733+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+  k1=0.42302944
+  k2=0.021354664
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=53438.0
+  ua=-1.9377487e-10
+  ub=7.2417962e-19
+  uc=-9.8608028e-11
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0115624
+  a0=1.109596
+  keta=4.9707517e-6
+  a1=0.0
+  a2=0.8
+  ags=0.18226013
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.25255658+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.745015+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.14877095
+  pdiblc1=0.39
+  pdiblc2=0.00019189
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=757128280.0
+  pscbe2=9.873241e-9
+  pvag=0.0
+  delta=0.01
+  alpha0=1.7815831e-11
+  alpha1=6.3056523e-17
+  beta0=9.6797043
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=9.2999e-10
+  bgidl=1352540500.0
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.4443203
+  kt2=-0.052664618
+  at=90000.0
+  ute=-0.17124159
+  ua1=2.1098632e-9
+  ub1=-7.3847396e-19
+  uc1=1.1059776e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.29 pmos
* DC IV MOS Parameters
+  lmin=4e-06 lmax=8e-06 wmin=2e-06 wmax=3.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.05272753391057+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0=3.97725303832486e-8
+  k1=0.39038913267053 lk1=2.62035995557297e-7
+  k2=0.034157405339651 lk2=-1.02780253841822e-7
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=77219.105207405 lvsat=-0.190914427231785
+  ua=-1.0058910972481e-10 lua=-7.48094165260102e-16
+  ub=6.7005208117432e-19 lub=4.34535232162094e-25
+  uc=-1.12073391491597e-10 luc=1.08099776526179e-16
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0118223059257 lu0=-2.08652165264849e-9
+  a0=1.126087589869 la0=-1.32394285569253e-7
+  keta=0.00976751116514225 lketa=-7.83735572886294e-08 wketa=2.14549971380942e-24 pketa=-4.92051989631606e-29
+  a1=0.0
+  a2=0.8
+  ags=0.0153421702244496 lags=1.3400153780626e-6
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.25352266271189+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff=7.75570041805986e-9
+  nfactor={1.8016792246885+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor=-4.54899715828586e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-0.11702082281515 lpclm=2.13377316265875e-06 ppclm=8.07793566946316e-28
+  pdiblc1=0.39
+  pdiblc2=0.00016861829933 lpdiblc2=1.86824933718352e-10
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=713956586.575161 lpscbe1=346.581836754292
+  pscbe2=1.02377817685766e-08 lpscbe2=-2.92652891564374e-15
+  pvag=0.0
+  delta=0.01
+  alpha0=2.1094013061788e-11 lalpha0=-2.63172062538493e-17 walpha0=-2.46519032881566e-32
+  alpha1=-8.91472829004879e-13 lalpha1=7.15723939058718e-18 walpha1=4.95588418306676e-35 palpha1=-2.12226091902608e-39
+  beta0=16.4061464909871 lbeta0=-5.39997971919381e-05 pbeta0=5.16987882845642e-26
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=1.81945162932607e-09 lagidl=-7.14058728669014e-15
+  bgidl=1707547725.8785 lbgidl=-2849.99374926589
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.43571310391217 lkt1=-6.90984669067463e-8
+  kt2=-0.053910290407949 lkt2=1.00002431429455e-8
+  at=133983.88685519 lat=-0.353102115866823
+  ute=-0.18700153612868 lute=1.2652065840169e-7
+  ua1=2.0378836586382e-09 lua1=5.77850894298032e-16
+  ub1=-5.52464897949799e-19 lub1=-1.49327851803026e-24
+  uc1=3.5322306333165e-10 luc1=-1.94779302364285e-15
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.30 pmos
* DC IV MOS Parameters
+  lmin=2e-06 lmax=4e-06 wmin=2e-06 wmax=3.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.05054614534106+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0=3.09859234019265e-8
+  k1=0.39687564013418 lk1=2.35908421331804e-7
+  k2=0.0302709592108142 lk2=-8.71256954722211e-8
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=35103.256068578 lvsat=-0.0212722922907794
+  ua=2.3768542641842e-10 lua=-2.1106599375506e-15
+  ub=5.0252413465642e-19 lub=1.10933579040084e-24
+  uc=-1.06253877880466e-10 luc=8.46588455347066e-17
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0136504793172 lu0=-9.4503821355298e-9
+  a0=1.258078200496 la0=-6.64050881287482e-7
+  keta=0.00257644639341079 lketa=-4.94080346808724e-8
+  a1=0.0
+  a2=0.8
+  ags=0.0976489959038203 lags=1.008484471908e-6
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.25972833662654+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff=3.27520804781837e-8
+  nfactor={1.7996233243084+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor=-4.46618573768344e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.40960767377198 lpclm=1.25198979477494e-8
+  pdiblc1=0.39
+  pdiblc2=0.000215
+  pdiblcb=-0.048993466222987 lpdiblcb=9.6645394024597e-8
+  drout=0.56
+  pscbe1=800000000.0
+  pscbe2=9.9958877548046e-09 lpscbe2=-1.95218273089826e-15 wpscbe2=1.26217744835362e-29
+  pvag=0.0
+  delta=0.01
+  alpha0=-2.1814048429144e-11 lalpha0=1.46515950534887e-16 palpha0=9.4039548065783e-38
+  alpha1=-9.96162012334853e-11 lalpha1=4.04819260707093e-16 walpha1=4.62223186652937e-33 palpha1=7.93458686805044e-38
+  beta0=-0.565983882178802 lbeta0=1.43637402856096e-5
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.40356585449e-11 lagidl=-2.95129413752347e-17
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.43080083823386 lkt1=-8.88850141117907e-8
+  kt2=-0.046587403054394 lkt2=-1.94962592425256e-8
+  at=65684.68564562 lat=-0.0779937529850897
+  ute=0.748393474846899 lute=-3.64123922106781e-06 wute=-2.11758236813575e-22 pute=-1.61558713389263e-27
+  ua1=4.5715420331244e-09 lua1=-9.62769463423188e-15
+  ub1=-2.48259222055664e-18 lub1=6.28125117590222e-24 pub1=2.80259692864963e-45
+  uc1=-2.7275176299186e-10 luc1=5.73626065090336e-16 puc1=3.76158192263132e-37
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.31 pmos
* DC IV MOS Parameters
+  lmin=1e-06 lmax=2e-06 wmin=2e-06 wmax=3.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.057002778272+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0=4.40798975062762e-8
+  k1=0.5465315097348 lk1=-6.75918863478171e-8
+  k2=-0.0273837315122164 lk2=2.97973254577963e-8
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=-31079.385260264 lvsat=0.112945310132416
+  ua=-2.3349070054076e-10 lua=-1.15512040619091e-15
+  ub=7.19732859340241e-19 lub=6.68839103246746e-25
+  uc=-9.9883306685304e-11 luc=7.17394035977723e-17
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0114019542504 lu0=-4.89040028236019e-9
+  a0=0.805550448148 la0=2.53669970141233e-7
+  keta=-0.0360500734855628 lketa=2.89260841154475e-8
+  a1=0.0
+  a2=0.8
+  ags=0.54743751849968 lags=9.63187455458712e-8
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.23543979096316+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff=-1.6504798664603e-8
+  nfactor={1.8160174582484+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor=-4.79865680669056e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=-0.34147508 leta0=8.5474640453904e-07 weta0=-2.11758236813575e-22 peta0=2.01948391736579e-28
+  etab=23.269005741064 letab=-4.73312235748089e-05 wetab=5.29395592033938e-21 petab=1.66607423182678e-26
+  dsub=0.8683964 ldsub=-6.254241984432e-7
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.19864536932944 lpclm=4.40348919809567e-7
+  pdiblc1=0.40428784073392 lpdiblc1=-2.89755695543012e-8
+  pdiblc2=-6.01742000000014e-06 lpdiblc2=4.4822067555096e-10
+  pdiblcb=-0.00191392161550472 lpdiblcb=1.16864251515819e-9
+  drout=0.35500804941008 ldrout=4.1572121589295e-7
+  pscbe1=800000000.0
+  pscbe2=1.07457079057876e-08 lpscbe2=-3.47280899924998e-15
+  pvag=0.0
+  delta=0.01
+  alpha0=-5.21477910835981e-13 lalpha0=1.03334873034605e-16
+  alpha1=1.0e-10
+  beta0=4.0903966569572 lbeta0=4.92065642880828e-6
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-1.9412451351408e-10 lagidl=4.73752909638312e-16 pagidl=-1.88079096131566e-37
+  bgidl=796023845.4724 lbgidl=413.661193668118
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.50037081952 lkt1=5.22020730967256e-8
+  kt2=-0.062375095928 lkt2=1.25209924528329e-8
+  at=-11392.425196 lat=0.0783177028763856
+  ute=-1.705269317 lute=1.3347594768442e-06 wute=-1.6940658945086e-21
+  ua1=-6.1588998352e-10 lua1=8.92355246338758e-16 pua1=-3.76158192263132e-37
+  ub1=7.1971953396e-19 lub1=-2.12998634516472e-25
+  uc1=-7.6614983716e-11 luc1=1.75863030360243e-16 wuc1=2.46519032881566e-32 puc1=-4.70197740328915e-38
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=2.745e-6
+  sbref=2.74e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.32 pmos
* DC IV MOS Parameters
+  lmin=5e-07 lmax=1e-06 wmin=2e-06 wmax=3.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.0394866987392+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0=2.60735779395127e-8
+  k1=0.51255790431576 lk1=-3.26674276603094e-8
+  k2=-0.014409803791552 lk2=1.64602834480859e-08 pk2=1.57772181044202e-30
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=67243.647498976 lvsat=0.0118704123323107
+  ua=-1.51159748745824e-09 lua=1.58758033478822e-16
+  ub=1.4650061637508e-18 lub=-9.72929104076568e-26
+  uc=-5.43216105211752e-11 luc=2.49025266814019e-17
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.00619932100248 lu0=4.57844264902592e-10
+  a0=1.102170850864 la0=-5.12522444059819e-8
+  keta=-0.0031753453814264 lketa=-4.86874187886744e-9
+  a1=0.0
+  a2=0.75650212045064 la2=4.47152982021872e-8
+  ags=0.25946033003624 lags=3.92355839560026e-7
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.24686093148736+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff=-4.76400325941179e-9
+  nfactor={1.1694703716344+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.84776965805096e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.49
+  etab=-46.8214378193087 letab=2.47209113199315e-5
+  dsub=0.22903159248344 ldsub=3.18351513061334e-8
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.63140089233904 lpclm=-4.5185647780253e-9
+  pdiblc1=0.5735410582276 lpdiblc1=-2.02965846099194e-7
+  pdiblc2=0.00026377467841408 lpdiblc2=1.70877635886467e-10
+  pdiblcb=0.235996908122958 lpdiblcb=-2.43400835526024e-07 wpdiblcb=1.05879118406788e-22 ppdiblcb=5.60091242706918e-29
+  drout=0.50535446117984 ldrout=2.61166908750579e-7
+  pscbe1=800000000.0
+  pscbe2=5.302172795176e-09 lpscbe2=2.12307977203741e-15
+  pvag=0.0
+  delta=0.01
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=8.3394846512288 lbeta0=5.52644959753011e-7
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.0288953917576e-10 lagidl=-2.42769172358211e-16
+  bgidl=1407952309.0552 lbgidl=-215.393923753437 wbgidl=1.81898940354586e-12
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.38742469288 lkt1=-6.39051897356744e-8
+  kt2=-0.044922511832 lkt2=-5.42005456684598e-9
+  at=55197.3460879999 lat=0.00986421707368904
+  ute=-0.50106417872 lute=9.68510451540152e-8
+  ua1=-6.88889430400002e-11 lua1=3.30044740737804e-16 pua1=-1.88079096131566e-37
+  ub1=6.1300667616e-19 lub1=-1.03299097252366e-25
+  uc1=1.6852615664e-10 luc1=-7.61391202320403e-17
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.745e-6
+  sbref=1.74e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.33 pmos
* DC IV MOS Parameters
+  lmin=2.5e-07 lmax=5e-07 wmin=2e-06 wmax=3.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.2077059122976+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0=1.14891304067785e-7
+  k1=0.0947761652936001 lk1=1.87916317162523e-7
+  k2=0.135789416375152 lk2=-6.28431024092917e-08 wk2=2.64697796016969e-23 pk2=1.26217744835362e-29
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=125426.330912 lvsat=-0.018849346317565
+  ua=-3.76671639473921e-10 lua=-4.40469195146724e-16
+  ub=6.96397207507201e-19 lub=3.08523395181488e-25
+  uc=-7.96074314597599e-12 luc=4.24545037705176e-19
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.01121512955344 lu0=-2.19044246030168e-9
+  a0=1.56573507888 la0=-2.96008594027694e-7
+  keta=0.059533124959296 lketa=-3.79780617171248e-08 wketa=-2.64697796016969e-23
+  a1=0.0
+  a2=0.88699575909872 la2=-2.41837770803352e-8
+  ags=1.111519731164 lags=-5.7521299522618e-8
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.21206765718896+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff=-2.31344345696753e-8
+  nfactor={1.1827048333296+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor=1.77789328843571e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.70917734797888 leta0=-1.15723009604673e-7
+  etab=-0.000928367896226464 letab=2.44175699153738e-10
+  dsub=0.0529810899339203 ldsub=1.24787704046249e-7
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.37128789943408 lpclm=1.32817974119879e-7
+  pdiblc1=-0.0311062144665597 lpdiblc1=1.1628065811605e-7
+  pdiblc2=-0.00739801875194496 lpdiblc2=4.21621262559488e-09 wpdiblc2=1.65436122510606e-24 ppdiblc2=-7.88860905221012e-31
+  pdiblcb=-0.3364671278616 lpdiblcb=5.88533059053904e-8
+  drout=1.46044604649312 ldrout=-2.4310998719581e-7
+  pscbe1=800000000.0
+  pscbe2=9.4308142774768e-09 lpscbe2=-5.67933869196181e-17
+  pvag=0.0
+  delta=0.01
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=9.9016510878832 lbeta0=-2.72160172803277e-7
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-2.75912561115488e-09 lagidl=1.47953568283456e-15 wagidl=-5.91645678915759e-31 pagidl=-2.35098870164458e-38
+  bgidl=1000000000.0
+  cgidl=566.002826479952 lcgidl=-0.000140446300347497
+  egidl=-1.3076004664448 legidl=7.43196155077257e-07 wegidl=2.11758236813575e-22 pegidl=-3.53409685539013e-28
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.47984947504 lkt1=-1.51060138525803e-8
+  kt2=-0.048887679968 lkt2=-3.32649337305561e-9
+  at=93529.3037919999 lat=-0.0103745966105305
+  ute=-0.33723371376 lute=1.0350525620715e-8
+  ua1=9.5015235456e-10 lua1=-2.07996835899425e-16
+  ub1=4.4478073632e-19 lub1=-1.44778197281242e-26
+  uc1=5.06950010616e-11 luc1=-1.39256840605121e-17
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.245e-6
+  sbref=1.24e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.34 pmos
* DC IV MOS Parameters
+  lmin=1.8e-07 lmax=2.5e-07 wmin=2e-06 wmax=3.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.154683777982859+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0=-1.77836213006102e-7
+  k1=-0.0222895163119983 lk1=2.204591718607e-7
+  k2=0.202818495717771 lk2=-8.14763821175879e-8
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=-59442.7774171428 lvsat=0.0325420473686367
+  ua=-1.13216897211429e-09 lua=-2.30450002640694e-16
+  ub=1.08735504518285e-18 lub=1.99841807801707e-25
+  uc=-2.62990061896749e-11 luc=5.52236210469693e-18
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.00269971039657143 lu0=1.76741880277903e-10
+  a0=-0.657791148 la0=3.22105014730224e-7
+  keta=-0.377120999460686 lketa=8.34065450221371e-08 wketa=-2.11758236813575e-22
+  a1=0.0
+  a2=1.180686884028 la2=-1.05826385517176e-7
+  ags=-0.121673607082855 lags=2.85291650189949e-7
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.268556120635429+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff=-7.43131959311844e-9
+  nfactor={1.01269644556572+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor=2.25049620541278e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.622334202767429 leta0=-9.15816573536319e-8
+  etab=0.232611176185622 letab=-6.46770150810711e-08 wetab=-3.94978742494071e-23 petab=3.94430452610506e-30
+  dsub=1.18577530834343 ldsub=-1.90115495140973e-7
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=1.49734406318857 lpclm=-1.80212126729905e-7
+  pdiblc1=1.00041477403886 lpdiblc1=-1.70469798436594e-7
+  pdiblc2=0.0188876887897257 lpdiblc2=-3.09089864249907e-9
+  pdiblcb=-0.494861204810126 lpdiblcb=1.02884958568157e-7
+  drout=-0.644450166046856 ldrout=3.42025901135754e-7
+  pscbe1=800000000.0
+  pscbe2=8.48238363300001e-09 lpscbe2=2.06858951077195e-16
+  pvag=0.0
+  delta=0.01
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=9.93867659484572 lbeta0=-2.8245281943277e-7
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=9.28298378178114e-09 lagidl=-1.86802622308894e-15
+  bgidl=1000000000.0
+  cgidl=-650.010094571257 lcgidl=0.000197590699549687 pcgidl=5.16987882845642e-26
+  egidl=5.12714452301714 legidl=-1.04558573505329e-06 pegidl=8.07793566946316e-28
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=0.261215537142856 lkt1=-2.21113194459268e-7
+  kt2=0.120707638971428 lkt2=-5.04719568943895e-8
+  at=20233.0185142858 lat=0.0100008911412507
+  ute=-0.3
+  ua1=4.01925318285714e-10 lua1=-5.55962985396092e-17
+  ub1=3.927e-19
+  uc1=6.0045e-13
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.1e-6
+  sbref=1.1e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.35 pmos
* DC IV MOS Parameters
+  lmin=1.5e-07 lmax=1.8e-07 wmin=2e-06 wmax=3.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.655380072203755+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0=-7.36973921636854e-08 wvth0=-4.63938843859879e-07 pvth0=9.6493712256728e-14
+  k1=1.13537408832746 lk1=-2.03209659410525e-08 wk1=-5.23677343759238e-06 pk1=1.08918603373796e-12
+  k2=-0.168045627012562 lk2=-4.34109495915141e-09 wk2=1.97427305956624e-06 pk2=-4.10625105113063e-13
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=431917.593817058 lvsat=-0.0696550135236222 wvsat=-0.260495700269901 pvsat=5.41799797077362e-8
+  ua=-2.38057911553099e-09 lua=2.92043262682609e-17 wua=4.70040942539538e-15 pua=-9.77628755569136e-22
+  ub=2.00636057944279e-18 lub=8.69968474205221e-27 wub=-4.19933402305312e-24 pub=8.73411084786774e-31
+  uc=-5.15107532176243e-13 luc=1.59620590721112e-19 wuc=3.27130020037795e-18 puc=-6.80391186076209e-25
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.000950824701720573 lu0=5.40489118178539e-10 wu0=1.62369803968332e-08 pu0=-3.37709707877655e-15
+  a0=-2.15964664451502 la0=6.3447293573939e-07 wa0=9.83442953452796e-06 pa0=-2.0454433300274e-12
+  keta=-0.5449792734476 lketa=1.18319051712127e-07 wketa=1.86923819148773e-06 pketa=-3.88779112971151e-13
+  a1=0.0
+  a2=-1.27188959606534 la2=4.04280091424477e-7
+  ags=-12.7193944818877 lags=2.90546641949885e-06 wags=4.17041213249505e-05 pags=-8.6739567861338e-12
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.859739614646242+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff=1.15527752959202e-07 wvoff=1.09880959505373e-06 pvoff=-2.28539210056036e-13
+  nfactor={6.85878289689938+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor=-9.9086620829871e-07 wnfactor=-8.07773334856944e-06 pnfactor=1.68007160370226e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=-1.28630528404293 leta0=3.05392452229081e-07 weta0=1.74881101905496e-06 peta0=-3.63731706231202e-13
+  etab=-0.297163827087051 letab=4.55098282996057e-08 wetab=-4.8852341788632e-07 petab=1.0160700863934e-13
+  dsub=0.344676596942732 ldsub=-1.51770563541649e-08 wdsub=-1.05123836870656e-08 pdsub=2.18644965830532e-15
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=2.83116724889235 lpclm=-4.57631343478062e-07 wpclm=-3.24768056850837e-06 ppclm=6.75478586082918e-13
+  pdiblc1=1.13779011954 lpdiblc1=-1.99042221796686e-7
+  pdiblc2=0.0253659711166133 lpdiblc2=-4.43830362710378e-9
+  pdiblcb=-0.294959646075795 lpdiblcb=6.13078331701212e-08 wpdiblcb=8.77427914045966e-07 ppdiblcb=-1.82494476986592e-13
+  drout=1.0
+  pscbe1=580945406.108536 lpscbe1=45.560726874297 wpscbe1=653.963875977737 ppscbe1=-0.000136016638636857
+  pscbe2=5.92861474346898e-09 lpscbe2=7.38012234872975e-16 wpscbe2=9.14627315828109e-15 ppscbe2=-1.90231506164457e-21
+  pvag=0.0
+  delta=0.01
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=16.4346727555795 lbeta0=-1.63354206891147e-06 wbeta0=-2.22216965356937e-06 pbeta0=4.62184621906578e-13
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-9.79791607908776e-10 lagidl=2.66507904661891e-16 wagidl=4.35640262329887e-15 pagidl=-9.06079468814686e-22
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-2.4779732524977 lkt1=3.48605203520492e-07 wkt1=1.07610039876875e-06 pkt1=-2.23815969739114e-13
+  kt2=-0.098872768856284 lkt2=-4.80186703111902e-09 wkt2=-6.89244397760454e-08 pkt2=1.433545638014e-14
+  at=105527.85395772 lat=-0.00773941109295823 wat=0.425889739861059 pat=-8.85799552142221e-8
+  ute=0.731504505742421 lute=-2.14540559140355e-07 wute=-3.07944550570828e-06 pute=6.40487711841254e-13
+  ua1=1.40038431799035e-10 lua1=-1.1269687930177e-18 wua1=-1.61761440290717e-17 pua1=3.3644438443184e-24
+  ub1=2.86333827945026e-19 lub1=2.21228873933699e-26 wub1=3.17544740396779e-25 pub1=-6.60454954656448e-32
+  uc1=-5.92675497788958e-10 luc1=1.2339427782873e-16 wuc1=1.10900126910266e-15 puc1=-2.30658955958124e-22
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.04e-6
+  sbref=1.04e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.36 pmos
* DC IV MOS Parameters
+  lmin=2.0e-05 lmax=1.0e-04 wmin=1.68e-06 wmax=2.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.0477733+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+  k1=0.42302944
+  k2=0.021354664
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=53438.0
+  ua=-1.9377487e-10
+  ub=7.2417962e-19
+  uc=-9.8608028e-11
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0115624
+  a0=1.109596
+  keta=4.9707517e-6
+  a1=0.0
+  a2=0.8
+  ags=0.18226013
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.25255658+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.745015+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.14877095
+  pdiblc1=0.39
+  pdiblc2=0.00019189
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=757128280.0
+  pscbe2=9.873241e-9
+  pvag=0.0
+  delta=0.01
+  alpha0=1.7815831e-11
+  alpha1=6.3056523e-17
+  beta0=9.6797043
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=9.2999e-10
+  bgidl=1352540500.0
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.4443203
+  kt2=-0.052664618
+  at=90000.0
+  ute=-0.17124159
+  ua1=2.1098632e-9
+  ub1=-7.3847396e-19
+  uc1=1.1059776e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.37 pmos
* DC IV MOS Parameters
+  lmin=8e-06 lmax=2.0e-05 wmin=1.68e-06 wmax=2.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.0477733+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+  k1=0.42302944
+  k2=0.021354664
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=53438.0
+  ua=-1.9377487e-10
+  ub=7.2417962e-19
+  uc=-9.8608028e-11
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0115624
+  a0=1.109596
+  keta=4.9707517e-6
+  a1=0.0
+  a2=0.8
+  ags=0.18226013
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.25255658+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.745015+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.14877095
+  pdiblc1=0.39
+  pdiblc2=0.00019189
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=757128280.0
+  pscbe2=9.873241e-9
+  pvag=0.0
+  delta=0.01
+  alpha0=1.7815831e-11
+  alpha1=6.3056523e-17
+  beta0=9.6797043
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=9.2999e-10
+  bgidl=1352540500.0
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.4443203
+  kt2=-0.052664618
+  at=90000.0
+  ute=-0.17124159
+  ua1=2.1098632e-9
+  ub1=-7.3847396e-19
+  uc1=1.1059776e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.38 pmos
* DC IV MOS Parameters
+  lmin=4e-06 lmax=8e-06 wmin=1.68e-06 wmax=2.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.05272753391057+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0=3.97725303832486e-8
+  k1=0.39038913267053 lk1=2.62035995557296e-7
+  k2=0.034157405339651 lk2=-1.02780253841822e-07 pk2=-2.01948391736579e-28
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=77219.1052074048 lvsat=-0.190914427231785
+  ua=-1.0058910972481e-10 lua=-7.48094165260102e-16
+  ub=6.7005208117432e-19 lub=4.34535232162091e-25
+  uc=-1.12073391491597e-10 luc=1.08099776526179e-16
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0118223059257 lu0=-2.08652165264849e-9
+  a0=1.126087589869 la0=-1.32394285569253e-7
+  keta=0.00976751116514225 lketa=-7.83735572886293e-08 wketa=-2.42984304937452e-24 pketa=2.89906382668722e-29
+  a1=0.0
+  a2=0.8
+  ags=0.0153421702244501 lags=1.3400153780626e-6
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.25352266271189+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff=7.75570041805986e-9
+  nfactor={1.8016792246885+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor=-4.54899715828579e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-0.11702082281515 lpclm=2.13377316265875e-06 ppclm=-1.61558713389263e-27
+  pdiblc1=0.39
+  pdiblc2=0.00016861829933 lpdiblc2=1.86824933718352e-10
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=713956586.575159 lpscbe1=346.581836754289
+  pscbe2=1.02377817685766e-08 lpscbe2=-2.92652891564369e-15
+  pvag=0.0
+  delta=0.01
+  alpha0=2.1094013061788e-11 lalpha0=-2.63172062538494e-17
+  alpha1=-8.91472829004879e-13 lalpha1=7.15723939058718e-18 walpha1=-1.97483050938144e-35 palpha1=-5.49147568432238e-39
+  beta0=16.4061464909871 lbeta0=-5.39997971919381e-5
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=1.81945162932607e-09 lagidl=-7.14058728669013e-15
+  bgidl=1707547725.8785 lbgidl=-2849.99374926589
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.43571310391217 lkt1=-6.90984669067463e-8
+  kt2=-0.0539102904079489 lkt2=1.00002431429453e-8
+  at=133983.88685519 lat=-0.353102115866823
+  ute=-0.18700153612868 lute=1.26520658401691e-7
+  ua1=2.0378836586382e-09 lua1=5.77850894298026e-16
+  ub1=-5.52464897949799e-19 lub1=-1.49327851803027e-24
+  uc1=3.5322306333165e-10 luc1=-1.94779302364285e-15 wuc1=-3.94430452610506e-31
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.39 pmos
* DC IV MOS Parameters
+  lmin=2e-06 lmax=4e-06 wmin=1.68e-06 wmax=2.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.05054614534106+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0=3.09859234019248e-8
+  k1=0.396875640134181 lk1=2.35908421331805e-7
+  k2=0.0302709592108142 lk2=-8.71256954722211e-08 pk2=5.04870979341448e-29
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=35103.256068578 lvsat=-0.0212722922907793
+  ua=2.3768542641842e-10 lua=-2.1106599375506e-15 pua=-1.50463276905253e-36
+  ub=5.0252413465642e-19 lub=1.10933579040084e-24
+  uc=-1.06253877880466e-10 luc=8.46588455347064e-17
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0136504793172 lu0=-9.4503821355298e-9
+  a0=1.258078200496 la0=-6.64050881287481e-7
+  keta=0.00257644639341079 lketa=-4.94080346808724e-08 pketa=-5.04870979341448e-29
+  a1=0.0
+  a2=0.8
+  ags=0.0976489959038203 lags=1.008484471908e-6
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.25972833662654+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff=3.27520804781846e-8
+  nfactor={1.7996233243084+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor=-4.46618573768347e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.409607673771981 lpclm=1.25198979477494e-8
+  pdiblc1=0.39
+  pdiblc2=0.000215
+  pdiblcb=-0.0489934662229869 lpdiblcb=9.66453940245971e-8
+  drout=0.56
+  pscbe1=800000000.0
+  pscbe2=9.9958877548046e-09 lpscbe2=-1.95218273089831e-15
+  pvag=0.0
+  delta=0.01
+  alpha0=-2.18140484291439e-11 lalpha0=1.46515950534887e-16
+  alpha1=-9.96162012334852e-11 lalpha1=4.04819260707094e-16 walpha1=-8.62816615085482e-32 palpha1=3.70280720509021e-37
+  beta0=-0.565983882178799 lbeta0=1.43637402856096e-5
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.40356585449001e-11 lagidl=-2.95129413752348e-17
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.43080083823386 lkt1=-8.88850141117899e-8
+  kt2=-0.046587403054394 lkt2=-1.94962592425257e-8
+  at=65684.68564562 lat=-0.0779937529850898 wat=1.11022302462516e-16
+  ute=0.748393474846899 lute=-3.64123922106781e-06 pute=-1.61558713389263e-27
+  ua1=4.5715420331244e-09 lua1=-9.62769463423188e-15
+  ub1=-2.48259222055664e-18 lub1=6.28125117590222e-24 pub1=-5.60519385729927e-45
+  uc1=-2.7275176299186e-10 luc1=5.73626065090336e-16
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.40 pmos
* DC IV MOS Parameters
+  lmin=1e-06 lmax=2e-06 wmin=1.68e-06 wmax=2.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.057002778272+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0=4.40798975062779e-8
+  k1=0.5465315097348 lk1=-6.75918863478176e-8
+  k2=-0.0273837315122164 lk2=2.97973254577963e-8
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=-31079.385260264 lvsat=0.112945310132416
+  ua=-2.33490700540761e-10 lua=-1.15512040619091e-15
+  ub=7.19732859340241e-19 lub=6.6883910324675e-25
+  uc=-9.9883306685304e-11 luc=7.17394035977723e-17
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0114019542504 lu0=-4.89040028236019e-9
+  a0=0.805550448148001 la0=2.53669970141232e-7
+  keta=-0.0360500734855628 lketa=2.89260841154475e-8
+  a1=0.0
+  a2=0.8
+  ags=0.54743751849968 lags=9.63187455458712e-8
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.23543979096316+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff=-1.65047986646032e-8
+  nfactor={1.8160174582484+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor=-4.79865680669059e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=-0.34147508 leta0=8.54746404539041e-07 weta0=2.11758236813575e-22 peta0=2.01948391736579e-28
+  etab=23.269005741064 letab=-4.73312235748089e-05 wetab=9.10560418298373e-21 petab=2.24162714827603e-26
+  dsub=0.868396400000001 ldsub=-6.254241984432e-7
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.19864536932944 lpclm=4.40348919809568e-7
+  pdiblc1=0.40428784073392 lpdiblc1=-2.89755695543016e-8
+  pdiblc2=-6.01742000000014e-06 lpdiblc2=4.4822067555096e-10
+  pdiblcb=-0.00191392161550472 lpdiblcb=1.16864251515819e-9
+  drout=0.355008049410081 ldrout=4.1572121589295e-7
+  pscbe1=800000000.0
+  pscbe2=1.07457079057876e-08 lpscbe2=-3.47280899924997e-15
+  pvag=0.0
+  delta=0.01
+  alpha0=-5.21477910836032e-13 lalpha0=1.03334873034605e-16
+  alpha1=1.0e-10
+  beta0=4.0903966569572 lbeta0=4.9206564288083e-6
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-1.9412451351408e-10 lagidl=4.73752909638312e-16 wagidl=9.86076131526265e-32 pagidl=-3.76158192263132e-37
+  bgidl=796023845.472403 lbgidl=413.661193668118
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.500370819520001 lkt1=5.22020730967264e-8
+  kt2=-0.0623750959280001 lkt2=1.25209924528329e-8
+  at=-11392.425196 lat=0.0783177028763857
+  ute=-1.705269317 lute=1.3347594768442e-6
+  ua1=-6.1588998352e-10 lua1=8.92355246338758e-16 pua1=7.52316384526264e-37
+  ub1=7.19719533960001e-19 lub1=-2.12998634516473e-25
+  uc1=-7.6614983716e-11 luc1=1.75863030360243e-16 wuc1=2.46519032881566e-32 puc1=-4.70197740328915e-38
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=2.745e-6
+  sbref=2.74e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.41 pmos
* DC IV MOS Parameters
+  lmin=5e-07 lmax=1e-06 wmin=1.68e-06 wmax=2.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.0394866987392+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0=2.60735779395135e-8
+  k1=0.512557904315759 lk1=-3.26674276603094e-8
+  k2=-0.014409803791552 lk2=1.6460283448086e-08 wk2=1.32348898008484e-23 pk2=9.46633086265214e-30
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=67243.6474989759 lvsat=0.0118704123323107
+  ua=-1.51159748745824e-09 lua=1.5875803347882e-16
+  ub=1.4650061637508e-18 lub=-9.72929104076575e-26
+  uc=-5.43216105211752e-11 luc=2.49025266814019e-17 puc=-4.70197740328915e-38
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.00619932100247998 lu0=4.57844264902599e-10
+  a0=1.102170850864 la0=-5.12522444059819e-8
+  keta=-0.0031753453814264 lketa=-4.86874187886743e-9
+  a1=0.0
+  a2=0.756502120450639 la2=4.47152982021876e-8
+  ags=0.25946033003624 lags=3.92355839560025e-7
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.24686093148736+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff=-4.76400325941179e-9
+  nfactor={1.1694703716344+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.84776965805098e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.49
+  etab=-46.8214378193087 letab=2.47209113199315e-5
+  dsub=0.22903159248344 ldsub=3.18351513061336e-8
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.63140089233904 lpclm=-4.51856477802572e-9
+  pdiblc1=0.5735410582276 lpdiblc1=-2.02965846099194e-7
+  pdiblc2=0.000263774678414079 lpdiblc2=1.70877635886466e-10
+  pdiblcb=0.235996908122957 lpdiblcb=-2.43400835526024e-07 wpdiblcb=-1.62127400060393e-22 ppdiblcb=-4.10207670714926e-29
+  drout=0.50535446117984 ldrout=2.61166908750579e-7
+  pscbe1=800000000.0
+  pscbe2=5.30217279517598e-09 lpscbe2=2.12307977203741e-15
+  pvag=0.0
+  delta=0.01
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=8.3394846512288 lbeta0=5.52644959753008e-7
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.0288953917576e-10 lagidl=-2.42769172358211e-16
+  bgidl=1407952309.0552 lbgidl=-215.393923753436
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.38742469288 lkt1=-6.39051897356744e-8
+  kt2=-0.0449225118319999 lkt2=-5.42005456684598e-9
+  at=55197.3460879999 lat=0.00986421707368906
+  ute=-0.501064178719999 lute=9.68510451540152e-8
+  ua1=-6.88889430400008e-11 lua1=3.30044740737803e-16 pua1=-3.76158192263132e-37
+  ub1=6.1300667616e-19 lub1=-1.03299097252366e-25
+  uc1=1.6852615664e-10 luc1=-7.61391202320403e-17
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.745e-6
+  sbref=1.74e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.42 pmos
* DC IV MOS Parameters
+  lmin=2.5e-07 lmax=5e-07 wmin=1.68e-06 wmax=2.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.2077059122976+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0=1.14891304067785e-7
+  k1=0.0947761652936006 lk1=1.87916317162523e-7
+  k2=0.135789416375152 lk2=-6.28431024092917e-08 wk2=-5.29395592033938e-23 pk2=-2.52435489670724e-29
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=125426.330912 lvsat=-0.0188493463175651
+  ua=-3.76671639473921e-10 lua=-4.40469195146724e-16
+  ub=6.96397207507204e-19 lub=3.08523395181489e-25
+  uc=-7.960743145976e-12 luc=4.24545037705176e-19
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.01121512955344 lu0=-2.19044246030168e-9
+  a0=1.56573507888 la0=-2.96008594027693e-7
+  keta=0.059533124959296 lketa=-3.79780617171248e-08 pketa=1.26217744835362e-29
+  a1=0.0
+  a2=0.886995759098721 la2=-2.41837770803352e-8
+  ags=1.111519731164 lags=-5.75212995226182e-8
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.21206765718896+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff=-2.31344345696753e-8
+  nfactor={1.1827048333296+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor=1.77789328843571e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.709177347978882 leta0=-1.15723009604673e-7
+  etab=-0.000928367896226465 letab=2.44175699153739e-10
+  dsub=0.0529810899339203 ldsub=1.24787704046249e-7
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.371287899434082 lpclm=1.32817974119879e-7
+  pdiblc1=-0.0311062144665599 lpdiblc1=1.1628065811605e-7
+  pdiblc2=-0.00739801875194495 lpdiblc2=4.21621262559487e-09 wpdiblc2=6.61744490042422e-24
+  pdiblcb=-0.3364671278616 lpdiblcb=5.88533059053906e-8
+  drout=1.46044604649312 ldrout=-2.4310998719581e-7
+  pscbe1=800000000.0
+  pscbe2=9.43081427747681e-09 lpscbe2=-5.67933869196181e-17
+  pvag=0.0
+  delta=0.01
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=9.90165108788321 lbeta0=-2.72160172803277e-7
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-2.75912561115488e-09 lagidl=1.47953568283456e-15 wagidl=1.77493703674728e-30 pagidl=-1.31655367292096e-36
+  bgidl=1000000000.0
+  cgidl=566.002826479952 lcgidl=-0.000140446300347497 pcgidl=2.06795153138257e-25
+  egidl=-1.3076004664448 legidl=7.43196155077258e-07 wegidl=-4.2351647362715e-22 pegidl=-4.03896783473158e-28
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.479849475040001 lkt1=-1.51060138525806e-8
+  kt2=-0.048887679968 lkt2=-3.32649337305563e-9
+  at=93529.3037919999 lat=-0.0103745966105305
+  ute=-0.337233713760001 lute=1.03505256207148e-8
+  ua1=9.5015235456e-10 lua1=-2.07996835899425e-16 wua1=-1.57772181044202e-30
+  ub1=4.44780736320002e-19 lub1=-1.4477819728124e-26
+  uc1=5.06950010616e-11 luc1=-1.39256840605121e-17
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.245e-6
+  sbref=1.24e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.43 pmos
* DC IV MOS Parameters
+  lmin=1.8e-07 lmax=2.5e-07 wmin=1.68e-06 wmax=2.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.154683777982864+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0=-1.77836213006101e-7
+  k1=-0.022289516312 lk1=2.20459171860702e-7
+  k2=0.202818495717771 lk2=-8.14763821175879e-8
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=-59442.7774171424 lvsat=0.0325420473686367
+  ua=-1.1321689721143e-09 lua=-2.30450002640695e-16
+  ub=1.08735504518286e-18 lub=1.99841807801708e-25
+  uc=-2.62990061896749e-11 luc=5.52236210469694e-18
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.00269971039657144 lu0=1.76741880277901e-10
+  a0=-0.657791147999998 la0=3.22105014730224e-7
+  keta=-0.377120999460686 lketa=8.34065450221371e-08 wketa=-4.2351647362715e-22 pketa=-1.0097419586829e-28
+  a1=0.0
+  a2=1.180686884028 la2=-1.05826385517176e-7
+  ags=-0.121673607082858 lags=2.8529165018995e-7
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.26855612063543+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff=-7.43131959311865e-9
+  nfactor={1.01269644556572+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor=2.25049620541278e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.62233420276743 leta0=-9.1581657353632e-8
+  etab=0.232611176185622 letab=-6.46770150810712e-08 wetab=-1.3648480107125e-23 petab=4.52115906304792e-29
+  dsub=1.18577530834343 ldsub=-1.90115495140973e-7
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=1.49734406318857 lpclm=-1.80212126729905e-7
+  pdiblc1=1.00041477403886 lpdiblc1=-1.70469798436594e-7
+  pdiblc2=0.0188876887897257 lpdiblc2=-3.09089864249907e-9
+  pdiblcb=-0.494861204810126 lpdiblcb=1.02884958568157e-7
+  drout=-0.644450166046855 ldrout=3.42025901135754e-7
+  pscbe1=800000000.0
+  pscbe2=8.48238363300005e-09 lpscbe2=2.06858951077198e-16
+  pvag=0.0
+  delta=0.01
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=9.93867659484576 lbeta0=-2.82452819432763e-7
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=9.28298378178115e-09 lagidl=-1.86802622308894e-15
+  bgidl=1000000000.0
+  cgidl=-650.010094571256 lcgidl=0.000197590699549687 wcgidl=-4.33680868994202e-19 pcgidl=1.03397576569128e-25
+  egidl=5.12714452301714 legidl=-1.04558573505329e-6
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=0.261215537142855 lkt1=-2.21113194459269e-7
+  kt2=0.120707638971428 lkt2=-5.04719568943896e-8
+  at=20233.0185142858 lat=0.0100008911412507
+  ute=-0.3
+  ua1=4.01925318285714e-10 lua1=-5.55962985396093e-17
+  ub1=3.927e-19
+  uc1=6.0045e-13
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.1e-6
+  sbref=1.1e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.44 pmos
* DC IV MOS Parameters
+  lmin=1.5e-07 lmax=1.8e-07 wmin=1.68e-06 wmax=2.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.06576568622668+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0=1.16578909257127e-08 wvth0=3.50837553213438e-07 pvth0=-7.29700010177535e-14
+  k1=-5.8336075143807 lk1=1.42914357964301e-06 wk1=8.5993882783679e-06 pk1=-1.78856956924118e-12
+  k2=2.57411961054937 lk2=-5.74678558389182e-07 wk2=-3.47000041420037e-06 pk2=7.21718446148706e-13
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=186963.406096112 lvsat=-0.018707481927918 wvsat=0.225834433388601 pvsat=-4.69708521316284e-8
+  ua=3.21091545248878e-09 lua=-1.13375944594503e-15 wua=-6.40090027629346e-15 pua=1.33131044666572e-21
+  ub=-3.40841716984992e-18 lub=1.13490847926194e-24 wub=6.55112348512614e-24 pub=-1.36255507142442e-30
+  uc=7.50245319750923e-13 luc=-1.03557618245515e-19 wuc=7.59078517914002e-19 puc=-1.57879222783897e-25
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.014534386875666 lu0=-2.28472881125602e-09 wu0=-1.0731717991533e-08 pu0=2.23206856162297e-15
+  a0=10.1659127171841 la0=-1.92909550478169e-06 wa0=-1.46366398828265e-05 pa0=3.04424545594931e-12
+  keta=2.45759646241143 lketa=-5.06180670437721e-07 wketa=-4.09205225439605e-06 pketa=8.51097764287326e-13
+  a1=0.0
+  a2=-1.27188959606533 la2=4.04280091424477e-7
+  ags=44.9043577558987 lags=-9.07958256093386e-06 wags=-7.27016269026832e-05 pags=1.51210659762353e-11
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.0505760503693384+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff=-5.27685584476216e-08 wvoff=-5.07697433985828e-07 pvoff=1.05594973899844e-13
+  nfactor={2.42294788309161+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor=-6.82657554468575e-08 wnfactor=7.29138888331404e-07 pnfactor=-1.5165213910627e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.211640034146233 leta0=-6.16219861044704e-09 weta0=-1.22519793170433e-06 peta0=2.5482646741932e-13
+  etab=-1.634369859887 letab=3.23632636649601e-07 wetab=2.16635500942764e-06 petab=-4.50575845700837e-13
+  dsub=0.330151342033462 ldsub=-1.21559776360958e-08 wdsub=1.83259441128108e-08 pdsub=-3.81157646413499e-15
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-0.526166193498042 lpclm=2.40653724537832e-07 wpclm=3.41794306081267e-06 ppclm=-7.10891141332306e-13
+  pdiblc1=1.13779011954 lpdiblc1=-1.99042221796686e-7
+  pdiblc2=0.0253659711166133 lpdiblc2=-4.43830362710378e-9
+  pdiblcb=0.918160911621315 lpdiblcb=-1.91006685384185e-07 wpdiblcb=-1.53109217886553e-06 ppdiblcb=3.18448800097883e-13
+  drout=1.0
+  pscbe1=1484545605.91082 lpscbe1=-142.377271482178 wpscbe1=-1140.03691262814 ppscbe1=0.000237113997383701
+  pscbe2=1.12801103999521e-08 lpscbe2=-3.75034643727644e-16 wpscbe2=-1.47854457643429e-15 ppscbe2=3.07519529363411e-22
+  pvag=0.0
+  delta=0.01
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=18.161524987624 lbeta0=-1.99270661094992e-06 wbeta0=-5.65064860562293e-06 pbeta0=1.17526710218632e-12
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.36463543920016e-09 lagidl=-1.0530567880122e-15 wagidl=-8.23977334950025e-15 pagidl=1.71377397941586e-21
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-2.5498929631214 lkt1=3.63563640293694e-07 wkt1=1.21888923126729e-06 pkt1=-2.53514333432821e-13
+  kt2=-0.133588549333332 lkt2=2.41859871874132e-9
+  at=731816.038326358 lat=-0.137999837983423 wat=-0.817537936336597 pat=1.70038080302776e-7
+  ute=-0.819546972000001 lute=1.08059535612336e-7
+  ua1=1.04739583685367e-09 lua1=-1.89846420755521e-16 wua1=-1.81763645863678e-15 pua1=3.78046571758947e-22
+  ub1=-9.47109584890814e-21 lub1=8.36467618834228e-26 wub1=9.04833528818852e-25 pub1=-1.88194515991975e-31
+  uc1=-3.40950474866667e-11 luc1=7.21624713125683e-18 wuc1=1.23259516440783e-32 puc1=5.87747175411144e-39
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.04e-6
+  sbref=1.04e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.45 pmos
* DC IV MOS Parameters
+  lmin=2.0e-05 lmax=1.0e-04 wmin=1.65e-06 wmax=1.68e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.0477733+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+  k1=0.42302944
+  k2=0.021354664
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=53438.0
+  ua=-1.9377487e-10
+  ub=7.2417962e-19
+  uc=-9.8608028e-11
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0115624
+  a0=1.109596
+  keta=4.9707517e-6
+  a1=0.0
+  a2=0.8
+  ags=0.18226013
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.25255658+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.745015+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.14877095
+  pdiblc1=0.39
+  pdiblc2=0.00019189
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=757128280.0
+  pscbe2=9.873241e-9
+  pvag=0.0
+  delta=0.01
+  alpha0=1.7815831e-11
+  alpha1=6.3056523e-17
+  beta0=9.6797043
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=9.2999e-10
+  bgidl=1352540500.0
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.4443203
+  kt2=-0.052664618
+  at=90000.0
+  ute=-0.17124159
+  ua1=2.1098632e-9
+  ub1=-7.3847396e-19
+  uc1=1.1059776e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.46 pmos
* DC IV MOS Parameters
+  lmin=8e-06 lmax=2.0e-05 wmin=1.65e-06 wmax=1.68e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.0477733+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+  k1=0.42302944
+  k2=0.021354664
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=53438.0
+  ua=-1.9377487e-10
+  ub=7.2417962e-19
+  uc=-9.8608028e-11
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0115624
+  a0=1.109596
+  keta=4.9707517e-6
+  a1=0.0
+  a2=0.8
+  ags=0.18226013
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.25255658+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.745015+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.14877095
+  pdiblc1=0.39
+  pdiblc2=0.00019189
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=757128280.0
+  pscbe2=9.873241e-9
+  pvag=0.0
+  delta=0.01
+  alpha0=1.7815831e-11
+  alpha1=6.3056523e-17
+  beta0=9.6797043
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=9.2999e-10
+  bgidl=1352540500.0
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.4443203
+  kt2=-0.052664618
+  at=90000.0
+  ute=-0.17124159
+  ua1=2.1098632e-9
+  ub1=-7.3847396e-19
+  uc1=1.1059776e-10
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.47 pmos
* DC IV MOS Parameters
+  lmin=4e-06 lmax=8e-06 wmin=1.65e-06 wmax=1.68e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.05272753391057+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0=3.9772530383269e-8
+  k1=0.390389132670528 lk1=2.62035995557316e-7
+  k2=0.0341574053396512 lk2=-1.02780253841821e-7
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=77219.1052074051 lvsat=-0.190914427231782
+  ua=-1.00589109724807e-10 lua=-7.48094165260124e-16
+  ub=6.70052081174317e-19 lub=4.34535232162091e-25
+  uc=-1.12073391491597e-10 luc=1.08099776526176e-16
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0118223059256999 lu0=-2.08652165264828e-9
+  a0=1.126087589869 la0=-1.32394285569273e-7
+  keta=0.00976751116514214 lketa=-7.83735572886297e-08 wketa=-3.6189151799195e-24 pketa=-3.7392006907476e-28
+  a1=0.0
+  a2=0.8
+  ags=0.0153421702244501 lags=1.3400153780626e-6
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.253522662711887+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff=7.75570041807003e-9
+  nfactor={1.80167922468848+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor=-4.54899715828525e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-0.117020822815149 lpclm=2.13377316265876e-6
+  pdiblc1=0.39
+  pdiblc2=0.000168618299329997 lpdiblc2=1.86824933718349e-10
+  pdiblcb=-0.025
+  drout=0.56
+  pscbe1=713956586.57515 lpscbe1=346.58183675434
+  pscbe2=1.02377817685768e-08 lpscbe2=-2.92652891564308e-15 wpscbe2=-2.01948391736579e-28
+  pvag=0.0
+  delta=0.01
+  alpha0=2.10940130617878e-11 lalpha0=-2.63172062538492e-17 walpha0=-3.94430452610506e-31
+  alpha1=-8.91472829004876e-13 lalpha1=7.15723939058718e-18 walpha1=-1.2172479101635e-33 palpha1=-3.5431282361455e-38
+  beta0=16.4061464909871 lbeta0=-5.39997971919382e-05 pbeta0=8.27180612553028e-25
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=1.81945162932607e-09 lagidl=-7.14058728669009e-15
+  bgidl=1707547725.87851 lbgidl=-2849.99374926591
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.435713103912178 lkt1=-6.90984669067768e-8
+  kt2=-0.0539102904079494 lkt2=1.0000243142947e-8
+  at=133983.886855191 lat=-0.353102115866825
+  ute=-0.187001536128683 lute=1.26520658401692e-7
+  ua1=2.03788365863822e-09 lua1=5.77850894298115e-16
+  ub1=-5.52464897949789e-19 lub1=-1.49327851803024e-24
+  uc1=3.53223063331649e-10 luc1=-1.94779302364286e-15 wuc1=3.15544362088405e-30
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.48 pmos
* DC IV MOS Parameters
+  lmin=2e-06 lmax=4e-06 wmin=1.65e-06 wmax=1.68e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.05054614534106+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0=3.09859234019316e-8
+  k1=0.396875640134176 lk1=2.35908421331797e-7
+  k2=0.030270959210814 lk2=-8.7125695472221e-08 pk2=-8.07793566946316e-28
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=35103.256068578 lvsat=-0.0212722922907789
+  ua=2.37685426418416e-10 lua=-2.1106599375506e-15 pua=-1.20370621524202e-35
+  ub=5.02524134656426e-19 lub=1.10933579040083e-24
+  uc=-1.06253877880465e-10 luc=8.46588455347068e-17
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0136504793171999 lu0=-9.4503821355298e-9
+  a0=1.258078200496 la0=-6.64050881287457e-7
+  keta=0.00257644639341081 lketa=-4.94080346808722e-08 pketa=4.03896783473158e-28
+  a1=0.0
+  a2=0.8
+  ags=0.0976489959038247 lags=1.00848447190801e-6
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.259728336626541+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff=3.27520804781854e-8
+  nfactor={1.79962332430839+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor=-4.46618573768354e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.409607673771973 lpclm=1.25198979477443e-8
+  pdiblc1=0.39
+  pdiblc2=0.000215
+  pdiblcb=-0.0489934662229872 lpdiblcb=9.66453940245963e-8
+  drout=0.56
+  pscbe1=800000000.0
+  pscbe2=9.99588775480453e-09 lpscbe2=-1.95218273089831e-15
+  pvag=0.0
+  delta=0.01
+  alpha0=-2.18140484291439e-11 lalpha0=1.46515950534886e-16
+  alpha1=-9.96162012334844e-11 lalpha1=4.04819260707093e-16 walpha1=-6.90253292068385e-31 palpha1=1.88079096131566e-36
+  beta0=-0.565983882178841 lbeta0=1.43637402856095e-5
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.40356585448996e-11 lagidl=-2.95129413752356e-17
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.430800838233857 lkt1=-8.88850141118034e-8
+  kt2=-0.046587403054394 lkt2=-1.94962592425255e-8
+  at=65684.6856456203 lat=-0.0779937529850887
+  ute=0.748393474846893 lute=-3.64123922106781e-06 pute=1.29246970711411e-26
+  ua1=4.57154203312436e-09 lua1=-9.62769463423185e-15
+  ub1=-2.48259222055661e-18 lub1=6.2812511759022e-24
+  uc1=-2.72751762991859e-10 luc1=5.73626065090341e-16
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.49 pmos
* DC IV MOS Parameters
+  lmin=1e-06 lmax=2e-06 wmin=1.65e-06 wmax=1.68e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.05700277827199+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0=4.40798975062694e-8
+  k1=0.546531509734791 lk1=-6.75918863478201e-8
+  k2=-0.0273837315122161 lk2=2.97973254577964e-8
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=-31079.3852602639 lvsat=0.112945310132417
+  ua=-2.3349070054076e-10 lua=-1.1551204061909e-15
+  ub=7.19732859340232e-19 lub=6.68839103246744e-25
+  uc=-9.98833066853036e-11 luc=7.17394035977729e-17
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0114019542504 lu0=-4.8904002823604e-9
+  a0=0.805550448147983 la0=2.53669970141227e-7
+  keta=-0.0360500734855624 lketa=2.89260841154472e-8
+  a1=0.0
+  a2=0.8
+  ags=0.547437518499663 lags=9.63187455458746e-8
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.235439790963159+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff=-1.65047986646045e-8
+  nfactor={1.81601745824841+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor=-4.79865680669056e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=-0.341475080000002 leta0=8.54746404539044e-07 weta0=-1.6940658945086e-21 peta0=-3.23117426778526e-27
+  etab=23.269005741064 letab=-4.73312235748095e-05 wetab=-5.59041745187838e-20 petab=-2.73034225627855e-25
+  dsub=0.868396400000002 ldsub=-6.25424198443206e-7
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.198645369329434 lpclm=4.40348919809558e-7
+  pdiblc1=0.404287840733915 lpdiblc1=-2.89755695542991e-8
+  pdiblc2=-6.01742000000058e-06 lpdiblc2=4.48220675550961e-10
+  pdiblcb=-0.00191392161550472 lpdiblcb=1.16864251515819e-9
+  drout=0.355008049410081 ldrout=4.15721215892958e-7
+  pscbe1=800000000.0
+  pscbe2=1.07457079057877e-08 lpscbe2=-3.47280899924986e-15
+  pvag=0.0
+  delta=0.01
+  alpha0=-5.21477910836549e-13 lalpha0=1.03334873034604e-16
+  alpha1=1.0e-10
+  beta0=4.09039665695707 lbeta0=4.92065642880839e-6
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-1.94124513514081e-10 lagidl=4.73752909638313e-16
+  bgidl=796023845.472382 lbgidl=413.661193668115
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.500370819520001 lkt1=5.22020730967256e-8
+  kt2=-0.0623750959280001 lkt2=1.25209924528334e-8
+  at=-11392.4251960004 lat=0.0783177028763866
+  ute=-1.70526931699999 lute=1.3347594768442e-06 pute=-2.58493941422821e-26
+  ua1=-6.1588998352e-10 lua1=8.92355246338761e-16 pua1=6.01853107621011e-36
+  ub1=7.19719533959987e-19 lub1=-2.12998634516469e-25
+  uc1=-7.66149837160004e-11 luc1=1.75863030360244e-16 wuc1=3.94430452610506e-31 puc1=1.1284745767894e-36
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=2.745e-6
+  sbref=2.74e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.50 pmos
* DC IV MOS Parameters
+  lmin=5e-07 lmax=1e-06 wmin=1.65e-06 wmax=1.68e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.0394866987392+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0=2.60735779395067e-8
+  k1=0.512557904315756 lk1=-3.26674276603115e-8
+  k2=-0.0144098037915521 lk2=1.64602834480861e-08 wk2=1.05879118406788e-22 pk2=2.52435489670724e-29
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=67243.6474989746 lvsat=0.0118704123323115
+  ua=-1.51159748745826e-09 lua=1.5875803347882e-16
+  ub=1.46500616375079e-18 lub=-9.7292910407656e-26
+  uc=-5.43216105211753e-11 luc=2.49025266814022e-17
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.00619932100248 lu0=4.57844264902573e-10
+  a0=1.102170850864 la0=-5.12522444059895e-8
+  keta=-0.00317534538142628 lketa=-4.86874187886741e-9
+  a1=0.0
+  a2=0.756502120450648 la2=4.47152982021884e-8
+  ags=0.259460330036234 lags=3.92355839560026e-7
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.246860931487362+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff=-4.76400325941179e-9
+  nfactor={1.16947037163436+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.84776965805099e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.49
+  etab=-46.8214378193088 letab=2.47209113199316e-5
+  dsub=0.229031592483441 ldsub=3.18351513061334e-8
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.63140089233903 lpclm=-4.51856477802742e-9
+  pdiblc1=0.573541058227605 lpdiblc1=-2.02965846099194e-7
+  pdiblc2=0.000263774678414083 lpdiblc2=1.70877635886466e-10
+  pdiblcb=0.235996908122957 lpdiblcb=-2.43400835526024e-07 wpdiblcb=-1.16467030247466e-21 ppdiblcb=-1.76704842769507e-28
+  drout=0.505354461179834 ldrout=2.61166908750577e-7
+  pscbe1=800000000.0
+  pscbe2=5.30217279517591e-09 lpscbe2=2.12307977203742e-15
+  pvag=0.0
+  delta=0.01
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=8.33948465122864 lbeta0=5.5264495975294e-7
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.02889539175754e-10 lagidl=-2.4276917235821e-16
+  bgidl=1407952309.05522 lbgidl=-215.393923753436
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.387424692880003 lkt1=-6.39051897356731e-8
+  kt2=-0.0449225118319996 lkt2=-5.4200545668464e-9
+  at=55197.3460880006 lat=0.00986421707368956
+  ute=-0.501064178720007 lute=9.68510451540169e-8
+  ua1=-6.88889430399988e-11 lua1=3.30044740737801e-16
+  ub1=6.13006676160004e-19 lub1=-1.03299097252362e-25
+  uc1=1.68526156640002e-10 luc1=-7.61391202320401e-17
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.745e-6
+  sbref=1.74e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.51 pmos
* DC IV MOS Parameters
+  lmin=2.5e-07 lmax=5e-07 wmin=1.65e-06 wmax=1.68e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.2077059122976+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0=1.14891304067776e-7
+  k1=0.0947761652936023 lk1=1.87916317162521e-7
+  k2=0.135789416375152 lk2=-6.28431024092917e-08 pk2=3.02922587604869e-28
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=125426.330912 lvsat=-0.0188493463175652
+  ua=-3.76671639473904e-10 lua=-4.40469195146719e-16
+  ub=6.96397207507188e-19 lub=3.08523395181492e-25
+  uc=-7.96074314597594e-12 luc=4.2454503770517e-19
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0112151295534401 lu0=-2.19044246030167e-9
+  a0=1.56573507888001 la0=-2.96008594027696e-7
+  keta=0.0595331249592963 lketa=-3.79780617171248e-08 pketa=-1.0097419586829e-28
+  a1=0.0
+  a2=0.88699575909871 la2=-2.41837770803373e-8
+  ags=1.11151973116399 lags=-5.7521299522622e-8
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.21206765718896+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff=-2.31344345696754e-8
+  nfactor={1.18270483332961+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor=1.77789328843567e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.709177347978887 leta0=-1.15723009604668e-7
+  etab=-0.000928367896226467 letab=2.44175699153738e-10
+  dsub=0.0529810899339225 ldsub=1.24787704046247e-7
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.371287899434066 lpclm=1.3281797411988e-7
+  pdiblc1=-0.0311062144665613 lpdiblc1=1.16280658116051e-7
+  pdiblc2=-0.00739801875194496 lpdiblc2=4.21621262559486e-09 wpdiblc2=3.97046694025453e-23 ppdiblc2=-6.31088724176809e-30
+  pdiblcb=-0.336467127861599 lpdiblcb=5.88533059053909e-8
+  drout=1.46044604649313 ldrout=-2.43109987195808e-7
+  pscbe1=800000000.0
+  pscbe2=9.4308142774766e-09 lpscbe2=-5.67933869196308e-17
+  pvag=0.0
+  delta=0.01
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=9.90165108788301 lbeta0=-2.72160172803244e-7
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-2.75912561115489e-09 lagidl=1.47953568283456e-15 wagidl=-1.10440526730942e-29 pagidl=-6.77084746073638e-36
+  bgidl=1000000000.0
+  cgidl=566.002826479955 lcgidl=-0.000140446300347498
+  egidl=-1.3076004664448 legidl=7.43196155077257e-07 wegidl=3.3881317890172e-21 pegidl=6.46234853557053e-27
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.479849475039998 lkt1=-1.51060138525791e-8
+  kt2=-0.0488876799679998 lkt2=-3.32649337305565e-9
+  at=93529.3037919998 lat=-0.0103745966105304
+  ute=-0.33723371376 lute=1.03505256207158e-8
+  ua1=9.50152354559999e-10 lua1=-2.07996835899423e-16
+  ub1=4.44780736319999e-19 lub1=-1.44778197281249e-26
+  uc1=5.06950010616002e-11 luc1=-1.3925684060512e-17
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.245e-6
+  sbref=1.24e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.52 pmos
* DC IV MOS Parameters
+  lmin=1.8e-07 lmax=2.5e-07 wmin=1.65e-06 wmax=1.68e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.15468377798291+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0=-1.77836213006108e-7
+  k1=-0.0222895163119858 lk1=2.20459171860698e-7
+  k2=0.202818495717768 lk2=-8.14763821175869e-08 pk2=8.07793566946316e-28
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=-59442.7774171401 lvsat=0.0325420473686364
+  ua=-1.13216897211434e-09 lua=-2.304500026407e-16
+  ub=1.08735504518291e-18 lub=1.99841807801707e-25
+  uc=-2.6299006189675e-11 luc=5.52236210469693e-18
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.00269971039657146 lu0=1.76741880277908e-10
+  a0=-0.657791147999973 la0=3.22105014730227e-7
+  keta=-0.377120999460683 lketa=8.3406545022137e-08 wketa=-3.3881317890172e-21
+  a1=0.0
+  a2=1.18068688402801 la2=-1.05826385517179e-7
+  ags=-0.121673607082812 lags=2.85291650189955e-7
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.268556120635438+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff=-7.4313195931178e-9
+  nfactor={1.01269644556584+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor=2.25049620541283e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.622334202767433 leta0=-9.15816573536328e-8
+  etab=0.232611176185621 letab=-6.46770150810708e-08 wetab=-2.18375681713999e-22 petab=7.09974814698911e-29
+  dsub=1.18577530834344 ldsub=-1.90115495140974e-7
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=1.49734406318856 lpclm=-1.802121267299e-7
+  pdiblc1=1.00041477403886 lpdiblc1=-1.70469798436593e-7
+  pdiblc2=0.0188876887897258 lpdiblc2=-3.09089864249909e-9
+  pdiblcb=-0.494861204810128 lpdiblcb=1.02884958568158e-7
+  drout=-0.644450166046852 ldrout=3.42025901135753e-7
+  pscbe1=800000000.0
+  pscbe2=8.48238363300058e-09 lpscbe2=2.06858951077166e-16
+  pvag=0.0
+  delta=0.01
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=9.93867659484613 lbeta0=-2.82452819432716e-7
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=9.28298378178108e-09 lagidl=-1.86802622308894e-15
+  bgidl=1000000000.0
+  cgidl=-650.010094571251 lcgidl=0.000197590699549686 pcgidl=1.65436122510606e-24
+  egidl=5.12714452301719 legidl=-1.04558573505328e-6
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=0.26121553714286 lkt1=-2.21113194459269e-7
+  kt2=0.120707638971425 lkt2=-5.04719568943894e-8
+  at=20233.0185142867 lat=0.0100008911412508
+  ute=-0.3
+  ua1=4.01925318285718e-10 lua1=-5.55962985396096e-17
+  ub1=3.927e-19
+  uc1=6.0045e-13
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.1e-6
+  sbref=1.1e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.53 pmos
* DC IV MOS Parameters
+  lmin=1.5e-07 lmax=1.8e-07 wmin=1.65e-06 wmax=1.68e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={4.94632011420754+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0=-1.23878381053499e-06 wvth0=-9.66164324456037e-06 pvth0=2.00950585514962e-12
+  k1=-0.670026059893303 lk1=3.55180600087097e-7
+  k2=-1.91120888457414 lk2=3.58215944654566e-07 wk2=3.99983067601606e-06 pk2=-8.31916782643231e-13
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=1227147.95420303 lvsat=-0.23505338571958 wvsat=-1.5064807995892 pvsat=3.13329928544957e-7
+  ua=6.73525794569108e-09 lua=-1.86678039242119e-15 wua=-1.2270312774601e-14 pua=2.5520778133637e-21
+  ub=1.09879805359291e-17 lub=-1.85936948676764e-24 wub=-1.7424524962176e-23 pub=3.62409209783309e-30
+  uc=1.20604096831587e-12 luc=-1.9835764359924e-19
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0783571856307834 lu0=-1.55591050787354e-08 wu0=-1.17021709220475e-07 pu0=2.43391112573483e-14
+  a0=1.3772082409493 la0=-1.01150438178568e-7
+  keta=0.000486206703467218 lketa=4.8687774264674e-9
+  a1=0.0
+  a2=-1.27188959606525 la2=4.04280091424478e-7
+  ags=1.25
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={5.80515516196859+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff=-1.27069038183936e-06 wvoff=-1.025978652031e-05 pvoff=2.13391247878623e-12
+  nfactor={-12.4261185639391+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor=3.02016187673818e-06 wnfactor=2.54586583264983e-05 pnfactor=-5.29509542801167e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=-0.524041285668005 leta0=1.46850687735076e-7
+  etab=-0.333562152592798 letab=5.30802432248948e-8
+  dsub=0.341155323025333 ldsub=-1.44446736346352e-8
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=1.52616902268267 lpclm=-1.86207372405165e-7
+  pdiblc1=1.13779011954 lpdiblc1=-1.99042221796684e-7
+  pdiblc2=0.0253659711166132 lpdiblc2=-4.4383036271038e-9
+  pdiblcb=-0.00119741061985267 lpdiblcb=2.08813342110715e-10
+  drout=1.0
+  pscbe1=800000000.0
+  pscbe2=1.03923047668799e-08 lpscbe2=-1.90381725716235e-16
+  pvag=0.0
+  delta=0.01
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=14.7685412774667 lbeta0=-1.28700671504171e-6
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=4.16988062503996e-10 lagidl=-2.40055054279194e-17
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=4.60711023176492 lkt1=-1.12500714020431e-06 wkt1=-1.07003280648715e-05 pkt1=2.22553983355647e-12
+  kt2=-0.133588549333332 lkt2=2.41859871874143e-9
+  at=240917.896533329 lat=-0.0358989152681755
+  ute=-0.819546971999998 lute=1.08059535612337e-7
+  ua1=-4.40206226666681e-11 lua1=3.71551058271973e-17
+  ub1=5.33844483999972e-19 lub1=-2.93563589381902e-26
+  uc1=-3.40950474866664e-11 luc1=7.21624713125679e-18 wuc1=-9.86076131526265e-32 puc1=2.35098870164458e-38
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.04e-6
+  sbref=1.04e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.54 pmos
* DC IV MOS Parameters
+  lmin=2.0e-05 lmax=1.0e-04 wmin=1.26e-06 wmax=1.65e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.137212577834+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} wvth0=1.46268297343356e-7
+  k1=0.203519229344934 wk1=3.58985286325653e-7
+  k2=0.0981375988951133 wk2=-1.25570212820576e-7
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=47690.62037634 wvsat=0.00939921980697256
+  ua=3.69523124728207e-09 wua=-6.36005026995538e-15
+  ub=-1.33842099521907e-18 wub=3.37316095784446e-24
+  uc=-2.8922147369136e-10 wuc=3.11727742298774e-16
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0285845955831707 wu0=-2.78379658835918e-8
+  a0=0.78132019602 wa0=5.36859689277621e-7
+  keta=-0.021183514387207 wketa=3.46514833259845e-8
+  a1=0.0
+  a2=0.8
+  ags=-0.1558799465992 wags=5.52991643777734e-7
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.252878050853266+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} wvoff=5.25730925959465e-10
+  nfactor={2.33929763662267+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} wnfactor=-9.71885188528142e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.618286094535021 wpclm=-7.67841405154446e-7
+  pdiblc1=0.39
+  pdiblc2=-0.00100863084676653 wpdiblc2=1.96332242873938e-9
+  pdiblcb=0.613662666666666 wpdiblcb=-1.04446394349787e-6
+  drout=0.56
+  pscbe1=620272418.5402 wpscbe1=223.813008355638
+  pscbe2=7.00331450793333e-09 wpscbe2=4.69345539969919e-15
+  pvag=0.0
+  delta=0.01
+  alpha0=7.47073616767133e-11 walpha0=-9.30399655147577e-17
+  alpha1=2.6441575864954e-16 walpha1=-3.2930132337922e-22
+  beta0=-55.209366896086 wbeta0=0.000106119080899324
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=3.52004831650547e-09 wagidl=-4.23576116835817e-15
+  bgidl=2478312779.19 wbgidl=-1841.07920436355
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.120870550460667 wkt1=-5.28967197488579e-7
+  kt2=-0.05324138786764 wkt2=9.43244942733505e-10
+  at=345465.066666667 wat=-0.417785577399147
+  ute=3.30390850076513 wute=-5.68323335226659e-6
+  ua1=9.66496536706933e-09 wua1=-1.23555551542283e-14
+  ub1=-4.67523521598747e-18 wub1=6.4381486513041e-24
+  uc1=4.376015395468e-10 wuc1=-5.34779430441356e-16
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.55 pmos
* DC IV MOS Parameters
+  lmin=8e-06 lmax=2.0e-05 wmin=1.26e-06 wmax=1.65e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.137212577834+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} wvth0=1.46268297343357e-7
+  k1=0.203519229344933 wk1=3.58985286325653e-7
+  k2=0.0981375988951133 wk2=-1.25570212820576e-7
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=47690.6203763401 wvsat=0.00939921980697256
+  ua=3.69523124728206e-09 wua=-6.36005026995538e-15
+  ub=-1.33842099521907e-18 wub=3.37316095784446e-24
+  uc=-2.8922147369136e-10 wuc=3.11727742298774e-16
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0285845955831707 wu0=-2.78379658835918e-8
+  a0=0.781320196020002 wa0=5.36859689277621e-7
+  keta=-0.021183514387207 wketa=3.46514833259845e-8
+  a1=0.0
+  a2=0.8
+  ags=-0.1558799465992 wags=5.52991643777734e-7
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.252878050853266+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} wvoff=5.25730925959677e-10
+  nfactor={2.33929763662267+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} wnfactor=-9.71885188528144e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.618286094535021 wpclm=-7.67841405154447e-7
+  pdiblc1=0.39
+  pdiblc2=-0.00100863084676653 wpdiblc2=1.96332242873938e-9
+  pdiblcb=0.613662666666666 wpdiblcb=-1.04446394349787e-6
+  drout=0.56
+  pscbe1=620272418.5402 wpscbe1=223.813008355638
+  pscbe2=7.00331450793334e-09 wpscbe2=4.6934553996992e-15
+  pvag=0.0
+  delta=0.01
+  alpha0=7.47073616767133e-11 walpha0=-9.30399655147577e-17
+  alpha1=2.6441575864954e-16 walpha1=-3.2930132337922e-22
+  beta0=-55.209366896086 wbeta0=0.000106119080899324
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=3.52004831650547e-09 wagidl=-4.23576116835817e-15
+  bgidl=2478312779.19 wbgidl=-1841.07920436355
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.120870550460667 wkt1=-5.28967197488579e-7
+  kt2=-0.0532413878676401 wkt2=9.43244942733452e-10
+  at=345465.066666667 wat=-0.417785577399147
+  ute=3.30390850076513 wute=-5.68323335226659e-6
+  ua1=9.66496536706933e-09 wua1=-1.23555551542283e-14
+  ub1=-4.67523521598747e-18 wub1=6.4381486513041e-24
+  uc1=4.376015395468e-10 wuc1=-5.34779430441356e-16
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.56 pmos
* DC IV MOS Parameters
+  lmin=4e-06 lmax=8e-06 wmin=1.26e-06 wmax=1.65e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.16848313722176+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0=2.5103967551823e-07 wvth0=1.89305810761418e-07 pvth0=-3.45504641270025e-13
+  k1=-0.0684463462446692 lk1=2.18333637724642e-06 wk1=7.50375963301182e-07 pk1=-3.14207965807141e-12
+  k2=0.190687381623033 lk2=-7.4298854514235e-07 wk2=-2.55987902280029e-07 pk2=1.04699164596821e-12
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=107242.108209568 lvsat=-0.478078629707302 wvsat=-0.0490993849303141 pvsat=4.6962609684768e-7
+  ua=5.94087624940628e-09 lua=-1.80280111293132e-14 wua=-9.88016532489318e-15 pua=2.82594414196601e-20
+  ub=-2.80617705308136e-18 lub=1.17831280194458e-23 wub=5.6849980115745e-24 pub=-1.85594001253001e-29
+  uc=-3.96023936194337e-10 luc=8.57408887344346e-16 wuc=4.64370505992611e-16 puc=-1.22541427522097e-21
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0367870931327305 lu0=-6.58495518978957e-08 wu0=-4.08272182730374e-08 pu0=1.04277562311441e-13
+  a0=0.602621409222692 la0=1.43459171602335e-06 wa0=8.56072508792763e-07 pa0=-2.56263668451372e-12
+  keta=0.00876325947860087 lketa=-2.40412341233419e-07 wketa=1.64234537500663e-09 pketa=2.64996963360795e-13
+  a1=0.0
+  a2=0.8
+  ags=-0.682951034216164 lags=4.23132036653594e-06 wags=1.14198325985519e-06 pags=-4.72841762597039e-12
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.220739138238022+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff=-2.58010804808232e-07 wvoff=-5.36139202130727e-08 pvoff=4.34632469668336e-13
+  nfactor={3.88350450622816+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.23968742187104e-05 wnfactor=-3.40460082719276e-06 pnfactor=1.95298119546119e-11
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-0.379651437465387 lpclm=8.01143053164889e-06 wpclm=4.29504058680203e-07 ppclm=-9.612275015519e-12
+  pdiblc1=0.39
+  pdiblc2=0.000405296608393313 lpdiblc2=-1.13509926428938e-08 wpdiblc2=-3.8706186055133e-10 ppdiblc2=1.88688568698144e-14
+  pdiblcb=0.613662666666666 wpdiblcb=-1.04446394349787e-6
+  drout=0.56
+  pscbe1=439287218.879787 lpscbe1=1452.9470110514 wpscbe1=449.192141507947 ppscbe1=-0.00180934097639713
+  pscbe2=4.45098752630226e-09 lpscbe2=2.04900503806104e-14 wpscbe2=9.46367816682035e-15 ppscbe2=-3.82952911317755e-20
+  pvag=0.0
+  delta=0.01
+  alpha0=8.84538062255031e-11 lalpha0=-1.1035629188035e-16 walpha0=-1.10159680333553e-16 palpha0=1.37436865128711e-22
+  alpha1=-3.73822490017055e-12 lalpha1=3.00125473664078e-17 walpha1=4.65555613251818e-18 palpha1=-3.73773923922548e-23
+  beta0=-27.0032871707239 lbeta0=-0.00022643806956225 wbeta0=7.09914492167796e-05 pbeta0=2.82004205615884e-10
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=7.47903123398794e-09 lagidl=-3.17826673537542e-14 wagidl=-9.2556323407431e-15 pagidl=4.02994655334521e-20
+  bgidl=3966969312.89599 lbgidl=-11950.9167887133 wbgidl=-3695.04043992003 pbgidl=0.0148835785515126
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=0.186398469974506 lkt1=-2.46675200882532e-06 wkt1=-1.01739641546399e-06 pkt1=3.921103900756e-12
+  kt2=0.02431255853778 lkt2=-6.22602151095355e-07 wkt2=-1.27925037027623e-07 pkt2=1.03455302123864e-12
+  at=675471.252361256 lat=-2.64928569868193 wat=-0.885544213947169 pat=3.75516072110389e-6
+  ute=7.0628460466625 lute=-3.01767055112135e-05 wute=-1.18563441880855e-05 pute=4.95576597126245e-11
+  ua1=1.63592766326956e-08 lua1=-5.37418505087121e-14 wua1=-2.34210943629082e-14 pua1=8.88340159808119e-20
+  ub1=-8.75036842041733e-18 lub1=3.27151204635645e-23 wub1=1.34067874769959e-23 pub1=-5.5944148868988e-29
+  uc1=1.1714002730292e-09 luc1=-5.8909274268119e-15 wuc1=-1.33804062695714e-15 puc1=6.44857124649433e-21
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.57 pmos
* DC IV MOS Parameters
+  lmin=2e-06 lmax=4e-06 wmin=1.26e-06 wmax=1.65e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.12867156978814+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0=9.0679159634416e-08 wvth0=1.27765709762442e-07 pvth0=-9.762185292737e-14
+  k1=0.265168445669288 lk1=8.39539998794508e-07 wk1=2.1539291851177e-07 pk1=-9.87174373456203e-13
+  k2=0.0856273628741691 lk2=-3.19808050342149e-07 wk2=-9.05294307711021e-08 pk2=3.80526908231913e-13
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=45318.1421598342 lvsat=-0.228649637546566 wvsat=-0.0167053450375289 pvsat=3.3914329288802e-7
+  ua=3.03286648306796e-09 lua=-6.31458268661959e-15 wua=-4.57121729763241e-15 pua=6.87506247322998e-21
+  ub=-5.22696945208319e-19 lub=2.58529754669449e-24 wub=1.67663855728637e-24 pub=-2.41377634374095e-30
+  uc=-2.40409777870372e-10 luc=2.30596924985318e-16 wuc=2.19397512427473e-16 puc=-2.38665996816509e-22
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0283131859947702 lu0=-3.17167556330772e-08 wu0=-2.39792761313862e-08 pu0=3.64142535401757e-14
+  a0=1.40658919479542 la0=-1.80378087665017e-06 wa0=-2.42873721691512e-07 pa0=1.86390554452218e-12
+  keta=-0.0255088303349823 lketa=-1.02364774729384e-07 wketa=4.59304424964556e-08 pketa=8.66050396127639e-14
+  a1=0.0
+  a2=0.8
+  ags=-0.359484025157291 lags=2.92839913565091e-06 wags=7.47591777005777e-07 pags=-3.13981346575076e-12
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.329461403567899+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff=1.79921175273331e-07 wvoff=1.14040913757977e-07 pvoff=-2.40679189709046e-13
+  nfactor={0.290510173684805+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor=2.07566383684219e-06 wnfactor=2.46799187544725e-06 pnfactor=-4.12492098050966e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=-0.17742104452954 leta0=1.03688887831245e-06 weta0=4.20984368339462e-07 peta0=-1.69571998385893e-12
+  etab=0.155041034103719 letab=-9.06462584877372e-07 wetab=-3.68030351853156e-07 petab=1.48242184090029e-12
+  dsub=-0.411400168036 ldsub=3.91278822004699e-06 wdsub=1.58862025788476e-06 pdsub=-6.39894333531674e-12
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=2.61390691618101 lpclm=-4.04658659413857e-06 wpclm=-3.60489378750164e-06 ppclm=6.63823109612733e-12
+  pdiblc1=0.39
+  pdiblc2=-0.0050772400939224 lpdiblc2=1.07325994035935e-08 wpdiblc2=8.65488817012797e-09 ppdiblc2=-1.75520093503615e-14
+  pdiblcb=0.513050544840932 lpdiblcb=4.05264419368596e-07 wpdiblcb=-9.19162391750647e-07 ppdiblcb=-5.04713146819179e-13
+  drout=0.56
+  pscbe1=800000128.626278 lpscbe1=-0.000260852548308321 wpscbe1=-0.000210354410228319 ppscbe1=4.26596220154396e-10
+  pscbe2=1.11468581127625e-08 lpscbe2=-6.48083599120423e-15 wpscbe2=-1.88228794583548e-15 ppscbe2=7.40612421840893e-21
+  pvag=0.0
+  delta=0.01
+  alpha0=-8.160051851811e-11 lalpha0=5.74620487535027e-16 walpha0=9.77743268490283e-17 palpha0=-7.00118820594641e-22
+  alpha1=-4.17731412310327e-10 lalpha1=1.69757213833627e-15 walpha1=5.2024313489642e-16 palpha1=-2.11415797260231e-21
+  beta0=-185.598762882832 lbeta0=0.000412382603460413 wbeta0=0.000302601163521992 pbeta0=-6.50916944288941e-10
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-7.16848772857567e-10 lagidl=1.23023896325937e-15 wagidl=1.26069838621703e-15 pagidl=-2.06018843877457e-21
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.364847550004784 lkt1=-2.46339655300978e-07 wkt1=-1.07859493134182e-07 pkt1=2.57500092054593e-13
+  kt2=-0.170792309756339 lkt2=1.63277917134937e-07 wkt2=2.03123735622088e-07 pkt2=-2.98907462409127e-13
+  at=-55858.7386285234 lat=0.296502729065006 wat=0.198771168019225 pat=-6.12448625672167e-7
+  ute=0.690267907861497 lute=-4.50803723906071e-06 wute=9.50580988685042e-08 pute=1.41755471760105e-12
+  ua1=6.32794014564931e-09 lua1=-1.33357475149277e-14 wua1=-2.87239977331795e-15 pua1=6.06412075827739e-21
+  ub1=-1.4615051626519e-18 lub1=3.35566672764443e-24 wub1=-1.66987781001835e-24 pub1=4.78447798712209e-30
+  uc1=-4.28906350315289e-10 luc1=5.55088448340219e-16 wuc1=2.55373994102955e-16 puc1=3.03162738397304e-23
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.58 pmos
* DC IV MOS Parameters
+  lmin=1e-06 lmax=2e-06 wmin=1.26e-06 wmax=1.65e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.1448185694017+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0=1.23425081086726e-07 wvth0=1.43613259850344e-07 pvth0=-1.29760494335035e-13
+  k1=0.79387414802023 lk1=-2.32668821104779e-07 wk1=-4.04502221379415e-07 pk1=2.69965531501442e-13
+  k2=-0.128470728595044 lk2=1.14380309980317e-07 wk2=1.65316886550679e-07 pk2=-1.38326353140851e-13
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=-381810.571122841 lvsat=0.637562267446141 wvsat=0.573583045656409 pvsat=-8.57954479978597e-7
+  ua=3.16896159175666e-09 lua=-6.59058193389897e-15 wua=-5.56434393969532e-15 pua=8.88911138581385e-21
+  ub=-1.20811943621247e-18 lub=3.97532613338102e-24 wub=3.15279460689899e-24 pub=-5.40740309848275e-30
+  uc=-2.87012869987101e-10 luc=3.25107436560938e-16 wuc=3.06030228213165e-16 puc=-4.14356104837304e-22
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0254502085362245 lu0=-2.5910671702876e-08 wu0=-2.29744054826539e-08 pu0=3.43763879229944e-14
+  a0=-1.67454845300352 la0=4.4447292994343e-06 wa0=4.05593439817176e-06 pa0=-6.85402573686312e-12
+  keta=-0.24421165376953 lketa=3.41161926761997e-07 wketa=3.40425824736073e-07 pketa=-5.10628061624594e-13
+  a1=0.0
+  a2=0.8
+  ags=3.49093756433381 lags=-4.88020964277798e-06 wags=-4.81377701565678e-06 pags=8.13857570934339e-12
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.199636694206759+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff=-8.33617774145498e-08 wvoff=-5.85521051712637e-08 pvoff=1.09337381563228e-13
+  nfactor={2.82345525672655+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor=-3.06111839622547e-06 wnfactor=-1.64755591761634e-06 pnfactor=4.22136055724979e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=-1.17253498357265 leta0=3.05496800532462e-06 weta0=1.35910888403547e-06 peta0=-3.59822524419625e-12
+  etab=97.5544912231146 letab=-0.000198431378774789 wetab=-0.000121485903530559 petab=2.47108015232837e-10
+  dsub=3.796003072144 ldsub=-4.61977506219917e-06 wdsub=-4.78778511629226e-06 pdsub=6.53233024664977e-12
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-0.22931844744514 lpclm=1.71944032459091e-06 wpclm=6.99888687835377e-07 ppclm=-2.09181610646645e-12
+  pdiblc1=0.424437536426877 lpdiblc1=-6.98389106232694e-08 wpdiblc1=-3.29526551686352e-08 ppdiblc1=6.68275892501298e-14
+  pdiblc2=-0.000711795294184933 lpdiblc2=1.87952973506352e-09 wpdiblc2=1.15422363037462e-09 ppdiblc2=-2.34075167171617e-15
+  pdiblcb=1.36700738435208 lpdiblcb=-1.32654980367794e-06 wpdiblcb=-2.23872322619321e-06 ppdiblcb=2.17134039070032e-12
+  drout=0.853457797042051 ldrout=-5.95128890907715e-07 wdrout=-8.15160829369292e-07 pdrout=1.65313638003097e-12
+  pscbe1=800000000.0
+  pscbe2=1.19731123413063e-08 lpscbe2=-8.15646965164032e-15 wpscbe2=-2.00728764009264e-15 ppscbe2=7.65962209836608e-21
+  pvag=0.0
+  delta=0.01
+  alpha0=3.06336815186522e-10 lalpha0=-2.12111769969963e-16 walpha0=-5.01833659036733e-16 palpha0=5.15878979485853e-22
+  alpha1=7.47619046947873e-10 lalpha1=-6.65744608833851e-16 walpha1=-1.05911113794999e-15 palpha1=1.08875354047893e-21
+  beta0=26.943601477197 lbeta0=-1.86507609533535e-05 wbeta0=-3.73739529080225e-05 pbeta0=3.85485121297318e-11
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-1.0542031428186e-09 lagidl=1.91438957728791e-15 wagidl=1.40656588175131e-15 pagidl=-2.35600596930814e-21
+  bgidl=144664071.537354 lbgidl=1734.6109988911 wbgidl=1065.22869368714 pbgidl=-0.00216027100805319
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.735007766417638 lkt1=5.04340821661694e-07 wkt1=3.83723432788211e-07 pkt1=-7.3942418272091e-13
+  kt2=-0.176395494710077 lkt2=1.74641108982899e-07 wkt2=1.86468070809098e-07 pkt2=-2.65129974036361e-13
+  at=-20741.8538763567 lat=0.225286108190229 wat=0.0152899827383116 pat=-2.40350983696698e-7
+  ute=-5.27204677078922 lute=7.5834653814668e-06 wute=5.83308002706275e-06 pute=-1.02190848965137e-11
+  ua1=-2.37914703018777e-09 lua1=4.32212079262382e-15 wua1=2.8836168207155e-15 pua1=-5.60901182222333e-21
+  ub1=-2.42128957956151e-19 lub1=8.82786417035899e-25 wub1=1.57299952126144e-24 pub1=-1.79203832618535e-30
+  uc1=-5.66195449366317e-10 luc1=8.33509093746516e-16 wuc1=8.00656074796896e-16 puc1=-1.07550924242261e-21
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=2.745e-6
+  sbref=2.74e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.59 pmos
* DC IV MOS Parameters
+  lmin=5e-07 lmax=1e-06 wmin=1.26e-06 wmax=1.65e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.937326459894059+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0=-8.9874317581819e-08 wvth0=-1.67072057757481e-07 pvth0=1.89620283942e-13
+  k1=0.887957685245111 lk1=-3.29385568369508e-07 wk1=-6.13925873613569e-07 pk1=4.85250532914325e-13
+  k2=-0.131553997279161 lk2=1.17549873188366e-07 wk2=1.91576700304927e-07 pk2=-1.65321126562453e-13
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=287749.806887545 lvsat=-0.0507377664240006 wvsat=-0.360614053116023 pvsat=1.02388927194277e-7
+  ua=-5.13726734439935e-09 lua=1.94812173772218e-15 wua=5.92939220381661e-15 pua=-2.92631144488269e-21
+  ub=3.89920672994557e-18 lub=-1.27494387751545e-24 wub=-3.98087261919051e-24 pub=1.92592120593054e-30
+  uc=1.83125086055043e-11 luc=1.12366112722829e-17 wuc=-1.18785271873642e-16 puc=2.2349131465933e-23
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=-0.00789810821079866 lu0=8.37099773326285e-09 wu0=2.30548257754481e-08 pu0=-1.29411094595593e-14
+  a0=4.82430819476674 la0=-2.23601734819375e-06 wa0=-6.08715437954725e-06 pa0=3.5729478095667e-12
+  keta=0.122642513329817 lketa=-3.59597547661261e-08 wketa=-2.05761544757069e-07 pketa=5.08459999659224e-14
+  a1=0.0
+  a2=0.617599761713941 la2=1.87505256155209e-07 wa2=2.27159834039599e-07 pa2=-2.33517583474699e-13
+  ags=-2.59619023946448 lags=1.37728469399302e-06 wags=4.67010866728703e-06 pags=-1.61074496609466e-12
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.263163280019567+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff=-1.80572095180129e-08 wvoff=2.66607336312529e-08 pvoff=2.17396058283072e-14
+  nfactor={-0.643670559204143+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor=5.03045337041487e-07 wnfactor=2.9651965357941e-06 pnfactor=-5.204936118267e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=3.18180398526346 leta0=-1.42124020257129e-06 weta0=-4.40215524142879e-06 peta0=2.3242851416115e-12
+  etab=-196.291022939917 letab=0.000103638283638638 wetab=0.000244441393643479 petab=-1.29060855134508e-10
+  dsub=-1.64585421998153 ldsub=9.74388931818378e-07 wdsub=3.06617363359588e-06 pdsub=-1.54144510073024e-12
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=2.32111193017591 lpclm=-9.02371498438997e-07 wpclm=-2.76334025153232e-06 ppclm=1.46834168445627e-12
+  pdiblc1=0.418673626660299 lpdiblc1=-6.39136805501449e-08 wpdiblc1=2.53268989619197e-07 ppdiblc1=-2.27404826932024e-13
+  pdiblc2=0.0014891195185207 lpdiblc2=-3.82984281420124e-10 wpdiblc2=-2.00391939382061e-09 ppdiblc2=9.05781459440242e-16
+  pdiblcb=1.06944181479077 lpdiblcb=-1.02065596895575e-06 wpdiblcb=-1.36300929949427e-06 ppdiblcb=1.27111698262093e-12
+  drout=-0.491545034084099 ldrout=7.87517879455995e-07 wdrout=1.63032165873858e-06 pdrout=-8.60790271954068e-13
+  pscbe1=800000000.0
+  pscbe2=-1.56219593460229e-09 lpscbe2=5.75766483229437e-15 wpscbe2=1.12259350786033e-14 ppscbe2=-5.94397205778075e-21
+  pvag=0.0
+  delta=0.01
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=6.98756819418803 lbeta0=1.86380178918031e-06 wbeta0=2.2109136288961e-06 pbeta0=-2.14425565182214e-12
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=1.83311053874086e-09 lagidl=-1.05373423959104e-15 wagidl=-2.17543304696496e-15 pagidl=1.32624594542504e-21
+  bgidl=2710671856.92529 lbgidl=-903.21421239427 wbgidl=-2130.45738737427 pbgidl=0.00112485593504497
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=0.0344448727151181 lkt1=-2.8664725793511e-07 wkt1=-6.89922196991645e-07 pkt1=3.64270640945225e-13
+  kt2=0.0448945178217516 lkt2=-5.2842368419671e-08 wkt2=-1.46886069722914e-07 pkt2=7.7554082180862e-14
+  at=299968.043039699 lat=-0.104399817320713 wat=-0.400296088583372 pat=1.86866510589137e-7
+  ute=4.92278758071041 lute=-2.89670199386261e-06 wute=-8.87012486132877e-06 pute=4.89563329029408e-12
+  ua1=3.1654279797503e-09 lua1=-1.3776357826924e-15 wua1=-5.28937666785927e-15 pua1=2.79272740810968e-21
+  ub1=1.27940151380933e-18 lub1=-6.81328649573358e-25 wub1=-1.08981691961199e-24 pub1=9.45305021235242e-31
+  uc1=4.77252595966668e-10 luc1=-2.39142975479249e-16 wuc1=-5.04888810808605e-16 puc1=2.66575233441214e-22
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.745e-6
+  sbref=1.74e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.60 pmos
* DC IV MOS Parameters
+  lmin=2.5e-07 lmax=5e-07 wmin=1.26e-06 wmax=1.65e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-2.07975597390621+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0=5.13314756662432e-07 wvth0=1.42614386876425e-06 pvth0=-6.51578606670354e-13
+  k1=-0.975762274849525 lk1=6.54636205920939e-07 wk1=1.75075021481023e-06 pk1=-7.63270065660382e-13
+  k2=0.536681092126767 lk2=-2.35270235196891e-07 wk2=-6.5561511956912e-07 pk2=2.81985988029205e-13
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=762754.910800918 lvsat=-0.301534761229014 wvsat=-1.04228218838741 pvsat=4.62301522599948e-7
+  ua=4.15988373254162e-10 lua=-9.83930642130266e-16 wua=-1.2963100020674e-15 pua=8.88772611397599e-22
+  ub=1.91353065663267e-19 lub=6.82758362981634e-25 wub=8.25945250227266e-25 pub=-6.12020947307607e-31
+  uc=1.13816472238423e-10 luc=-3.91883354783344e-17 wuc=-1.99153508177365e-16 puc=6.47825958154631e-23
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0188523964052498 lu0=-5.75294769795536e-09 wu0=-1.24899266387683e-08 pu0=5.82609327811797e-15
+  a0=1.79266250060043 la0=-6.35344801422266e-07 wa0=-3.71115335447697e-07 pa0=5.54947786750667e-13
+  keta=0.439202542680105 lketa=-2.03099651542726e-07 wketa=-6.20908404319153e-07 pketa=2.70038560052388e-13
+  a1=0.0
+  a2=0.183793948350163 la2=4.16549519941524e-07 wa2=1.15001075632407e-06 pa2=-7.20771796229831e-13
+  ags=-2.69407952106477 lags=1.42896906000659e-06 wags=6.22364733342076e-06 pags=-2.43099473934927e-12
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.264525644871572+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff=-1.73378972245326e-08 wvoff=8.57893838838389e-08 pvoff=-9.47961196125516e-15
+  nfactor={-1.19507566029197+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor=7.94180613554647e-07 wnfactor=3.88860367258087e-06 pnfactor=-1.00804149916447e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=1.40907929564448 leta0=-4.85262839148736e-07 weta0=-1.14461418597713e-06 peta0=6.04342554825691e-13
+  etab=-0.00407271239620571 letab=1.12936190922435e-09 wetab=5.14223646937897e-09 petab=-1.44762662349704e-15
+  dsub=0.311366999602107 ldsub=-5.90003854671497e-08 wdsub=-4.22562301261257e-07 pdsub=3.00565608043115e-13
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-0.404015103000011 lpclm=5.3646287355349e-07 wpclm=1.26792448281729e-06 ppclm=-6.60117720103511e-13
+  pdiblc1=0.463498165499105 lpdiblc1=-8.75804991625678e-08 wpdiblc1=-8.08872145081684e-07 ppdiblc1=3.33392946496425e-13
+  pdiblc2=0.00468698656823939 lpdiblc2=-2.07141970926699e-09 wpdiblc2=-1.9763723437588e-08 ppdiblc2=1.02827448769009e-14
+  pdiblcb=-2.04124148968242 lpdiblcb=6.21747487606441e-07 wpdiblcb=2.78797469408175e-06 ppdiblcb=-9.20552754179281e-13
+  drout=0.912796098788462 ldrout=4.60426133928776e-08 wdrout=8.95622452806606e-07 pdrout=-4.72877907612454e-13
+  pscbe1=799747395.294958 lpscbe1=0.133372253005973 wpscbe1=0.413107764308734 ppscbe1=-2.18115942262048e-7
+  pscbe2=9.41213875053695e-09 lpscbe2=-3.66521894429261e-17 wpscbe2=3.05418110883279e-17 ppscbe2=-3.29387572520408e-23
+  pvag=0.0
+  delta=0.01
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=13.6068399340374 lbeta0=-1.6310942581993e-06 wbeta0=-6.05943693852763e-06 pbeta0=2.22239020357078e-12
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-9.77542402835243e-09 lagidl=5.07543270941941e-15 wagidl=1.14743997043572e-14 pagidl=-5.88070194928006e-21
+  bgidl=1984841617.31006 lbgidl=-519.984555840304 wbgidl=-1610.60229918426 pbgidl=0.000850378686741698
+  cgidl=1415.43319898274 lcgidl=-0.000588935343864497 wcgidl=-0.00138915180563415 pcgidl=7.33455483553163e-10
+  egidl=-5.8025098039492 legidl=3.11645434636753e-06 wegidl=7.35093967026187e-06 pegidl=-3.88120793462222e-12
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.401305532454498 lkt1=-5.65762730104147e-08 wkt1=-1.28450151061577e-07 pkt1=6.78201383587002e-14
+  kt2=0.104727511900625 lkt2=-8.44334712973871e-08 wkt2=-2.51221086583453e-07 pkt2=1.32641719063024e-13
+  at=190157.372127418 lat=-0.04642110080708 wat=-0.15802478925681 pat=5.89501718003043e-8
+  ute=-0.449146735826713 lute=-6.03851379428055e-08 wute=1.8302168336633e-07 pute=1.15680552453606e-13
+  ua1=1.66248057888539e-09 lua1=-5.84097590404537e-16 wua1=-1.16493602190159e-15 pua1=6.15072240331775e-22
+  ub1=-2.95541006665669e-19 lub1=1.50222101927197e-25 wub1=1.21071640396917e-24 pub1=-2.69348967215724e-31
+  uc1=5.05951877602402e-11 luc1=-1.38729838351537e-17 wuc1=1.63233894500036e-19 puc1=-8.61855374892874e-26
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.245e-6
+  sbref=1.24e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.61 pmos
* DC IV MOS Parameters
+  lmin=1.8e-07 lmax=2.5e-07 wmin=1.26e-06 wmax=1.65e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={2.22484346353622+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0=-6.83312231753316e-07 wvth0=-3.89146029046782e-06 pvth0=8.2665153834625e-13
+  k1=3.25699492471341 lk1=-5.22019502471163e-07 wk1=-5.36291619643431e-06 pk1=1.21424383266867e-12
+  k2=-1.00997991442022 lk2=1.94682964691092e-07 wk2=1.98340106011207e-06 pk2=-4.51628841728009e-13
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=-1521119.01288601 lvsat=0.333354783068868 wvsat=2.39041391441115 pvsat=-4.9194680162482e-7
+  ua=-7.03564296571385e-09 lua=1.08753345052677e-15 wua=9.65449532203558e-15 pua=-2.15541985903914e-21
+  ub=5.69243973312517e-18 lub=-8.46477717532768e-25 wub=-7.5311195790003e-24 pub=1.7111427904397e-30
+  uc=-1.08808825423924e-10 luc=2.2698825768226e-17 wuc=1.34935914799101e-16 puc=-2.80902546989189e-23
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=-0.0234923292536868 lu0=6.01837789852111e-09 wu0=4.2834257346123e-08 pu0=-9.553365979474e-15
+  a0=-2.74344714060789 la0=6.25639245517952e-07 wa0=3.4108655421942e-06 pa0=-4.9639751346325e-13
+  keta=-1.19761119132802 lketa=2.51914924746724e-07 wketa=1.34182325995634e-06 pketa=-2.75577289836227e-13
+  a1=0.0
+  a2=4.82574774233174 la2=-8.73857931339827e-07 wa2=-5.96110409619524e-06 pa2=1.25603279939231e-12
+  ags=6.00088974435487 lags=-9.88128056148881e-07 wags=-1.00127923489471e-05 pags=2.08254065507281e-12
+  b0=0.0
+  b1=1.99947914368468e-23 lb1=-5.55831208194616e-30 wb1=-3.2699325956446e-29 pb1=9.09002022398052e-36
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.58750667077093+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff=7.24469522031785e-08 wvoff=5.2160924187731e-07 pvoff=-1.30632302645144e-13
+  nfactor={1.06256284363691+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor=1.66584201124464e-07 wnfactor=-8.15511184477273e-08 pnfactor=9.56138908839862e-14
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=-1.59877089367488 leta0=3.50883419279772e-07 weta0=3.63237795010199e-06 peta0=-7.23603935098672e-13
+  etab=0.676807644924325 letab=-1.88147206861595e-07 wetab=-7.26435440242819e-07 petab=2.01922188570373e-13
+  dsub=-0.434701030633388 ldsub=1.48397574121956e-07 wdsub=2.65011436504724e-06 pdsub=-5.53601633070653e-13
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=4.1009857964496 lpclm=-7.15873316482708e-07 wpclm=-4.25797538216956e-06 ppclm=8.76016131564455e-13
+  pdiblc1=-0.21865566962782 lpdiblc1=1.02050081156696e-07 wpdiblc1=1.99365829482302e-06 ppdiblc1=-4.45676885431805e-13
+  pdiblc2=-0.0391853663278757 lpdiblc2=1.01245679276182e-08 wpdiblc2=9.49722213694954e-08 ppdiblc2=-2.16124709481306e-14
+  pdiblcb=0.0666106693774444 lpdiblcb=3.57898816137075e-08 wpdiblcb=-9.18226723565734e-07 ppdiblcb=1.09726765509707e-13
+  drout=1.31144250432692 ldrout=-6.47763035899469e-08 wdrout=-3.19865161716644e-06 pdrout=6.65281152551214e-13
+  pscbe1=800902159.660864 lpscbe1=-0.187638383543799 wpscbe1=-1.47538487253405 ppscbe1=3.06862348868359e-7
+  pscbe2=7.85513692079348e-09 lpscbe2=3.96175635203805e-16 wpscbe2=1.02579438061818e-15 ppscbe2=-3.09607028550512e-22
+  pvag=0.0
+  delta=0.01
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=7.24841573438354 lbeta0=1.36471368214081e-07 wbeta0=4.39963162716508e-06 pbeta0=-6.85105348868998e-13
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=3.08768856488595e-08 lagidl=-6.22542155312938e-15 wagidl=-3.53144986809854e-14 pagidl=7.12605033506457e-21
+  bgidl=-2489269173.2653 lbgidl=723.764554610159 wbgidl=5706.32358965852 pbgidl=-0.00118363890724593
+  cgidl=-3683.68999636691 lcgidl=0.000828559714964361 wcgidl=0.00496125644869338 pcgidl=-1.03188180625084e-9
+  egidl=21.1803921569614 legidl=-4.38446860394209e-06 wegidl=-2.62533559652209e-05 pegidl=5.46038300049436e-12
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=1.8351044322773 lkt1=-6.78271406286277e-07 wkt1=-2.57392562276948e-06 pkt1=7.47632973787837e-13
+  kt2=-0.409321262373606 lkt2=5.84659193655578e-08 wkt2=8.66805131034239e-07 pkt2=-1.78156153120083e-13
+  at=-198016.981142164 lat=0.0614867113096245 wat=0.35692434708816 pat=-8.4199508713961e-8
+  ute=-0.959457948260193 lute=8.14752553791528e-08 wute=1.07847238481272e-06 pute=-1.33243997140075e-13
+  ua1=-1.99143215209431e-09 lua1=4.31646301855046e-16 wua1=3.91407813887122e-15 pua1=-7.96832748193137e-22
+  ub1=2.44849592666667e-19 wub1=2.41793402919755e-25
+  uc1=4.19143813318708e-12 luc1=-9.73298283828463e-19 wuc1=-5.8726739833067e-18 puc1=1.59172442164645e-24
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.1e-6
+  sbref=1.1e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.62 pmos
* DC IV MOS Parameters
+  lmin=1.5e-07 lmax=1.8e-07 wmin=1.26e-06 wmax=1.65e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.51385122841267+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0=9.42913998357504e-08 wvth0=9.03270579824166e-07 pvth0=-1.7059494590404e-13
+  k1=-2.8786037284572 lk1=7.54111390204487e-07 wk1=3.61189069226355e-06 pk1=-6.5240830249782e-13
+  k2=1.58581188824321 lk2=-3.45210580761269e-07 wk2=-1.71916981908741e-06 pk2=3.18461470294931e-13
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=635059.633148298 lvsat=-0.115104501162516 wvsat=-0.538184177625181 pvsat=1.17166458341633e-7
+  ua=2.91375518298587e-09 lua=-9.81821971624984e-16 wua=-6.02065696419456e-15 pua=1.10482371466929e-21
+  ub=-3.17865621549564e-18 lub=9.98603786628975e-25 wub=5.74348228133725e-24 pub=-1.04981510128818e-30
+  uc=3.04103421329749e-12 luc=-5.64602838000414e-19 wuc=-3.00093363989564e-18 puc=5.98954534211163e-25
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0180242998977479 lu0=-2.61658276542749e-09 wu0=-1.83537784891778e-08 pu0=3.17301121783853e-15
+  a0=-0.995446855747911 la0=2.62076162270492e-07 wa0=3.88022163842891e-06 pa0=-5.94017949206915e-13
+  keta=-0.98615600484481 lketa=2.07934783420454e-07 wketa=1.6135469769568e-06 pketa=-3.3209256228772e-13
+  a1=0.0
+  a2=-3.98600027042304 la2=9.58879914337014e-07 wa2=4.43863542678133e-06 pa2=-9.06988224512544e-13
+  ags=1.25
+  b0=0.0
+  b1=-4.66545133526427e-23 lb1=8.30394352261017e-30 wb1=7.62984272317077e-29 pb1=-1.35802044661172e-35
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-1.01373551645891+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff=1.6109743736013e-07 wvoff=8.91774107843087e-07 pvoff=-2.07622152787634e-13
+  nfactor={6.05631505776005+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor=-8.72056334386581e-07 wnfactor=-4.76736945544648e-06 pnfactor=1.07020787515968e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=-2.88612691530723 leta0=6.18638023507043e-07 weta0=3.86293641444409e-06 peta0=-7.71557328980257e-13
+  etab=-0.979181848994178 letab=1.56278735999526e-07 wetab=1.05584141566118e-06 petab=-1.68770010135388e-13
+  dsub=0.390269872085943 ldsub=-2.31864739928332e-08 wdsub=-8.03215504402415e-08 pdsub=1.42962721197574e-14
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=4.30419815299335 lpclm=-7.58139048095532e-07 wpclm=-4.54316717108289e-06 ppclm=9.3533260135696e-13
+  pdiblc1=4.09376441213614 lpdiblc1=-7.94881546809227e-07 wpdiblc1=-4.83417730151225e-06 ppdiblc1=9.74430984578775e-13
+  pdiblc2=0.105341514562286 lpdiblc2=-1.99352889749648e-08 wpdiblc2=-1.30791379941815e-07 ppdiblc2=2.53436489614062e-14
+  pdiblcb=-1.22221469936708 lpdiblcb=3.03850092408145e-07 wpdiblcb=1.99684215008237e-06 ppdiblcb=-4.96572579382616e-13
+  drout=1.0
+  pscbe1=800000000.0
+  pscbe2=9.62848312553808e-09 lpscbe2=2.73409047713684e-17 wpscbe2=1.2491479544417e-15 ppscbe2=-3.56061891662925e-22
+  pvag=0.0
+  delta=0.01
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=17.6681406545709 lbeta0=-2.03070637848585e-06 wbeta0=-4.74198220444115e-06 pbeta0=1.21624062873912e-12
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=7.12790547813983e-09 lagidl=-1.28591866538174e-15 wagidl=-1.0974981996375e-14 pagidl=2.06372293886582e-21
+  bgidl=934614593.368546 lbgidl=11.6378177555189 wbgidl=106.930783998905 pbgidl=-1.90323963823969e-5
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-7.5657952480431 lkt1=1.2770029164242e-06 wkt1=9.20714660814384e-06 pkt1=-1.70268867737536e-12
+  kt2=-0.176981045100124 lkt2=1.01419422552809e-08 wkt2=7.09637491155433e-08 pkt2=-1.26306957775774e-14
+  at=665986.148578232 lat=-0.118215571634661 wat=-0.695153303861862 pat=1.34620017751832e-7
+  ute=-2.67568311745295 lute=4.38429495869215e-07 wute=3.03551057441182e-06 pute=-5.40284456118411e-13
+  ua1=-4.88818078117511e-11 lua1=2.7619140848406e-17 wua1=7.94994426902696e-18 pua1=1.55950427457841e-23
+  ub1=-4.91192533348183e-19 lub1=1.53087929705576e-25 wub1=1.67633754288248e-24 pub1=-2.98367966582567e-31
+  uc1=-4.1642242286105e-11 luc1=8.55955723921926e-18 wuc1=1.2342623506882e-17 puc1=-2.19683887274292e-24
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.04e-6
+  sbref=1.04e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.63 pmos
* DC IV MOS Parameters
+  lmin=2.0e-05 lmax=1.0e-04 wmin=1e-06 wmax=1.26e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.019765+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+  k1=0.49177002
+  k2=-0.002690247
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=55237.817
+  ua=-1.4116341e-9
+  ub=1.370092e-18
+  uc=-3.8916596e-11
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0062318252
+  a0=1.212397
+  keta=0.0066402373
+  a1=0.0
+  a2=0.8
+  ags=0.28815017
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.25245591+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.5589128+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.0017402344
+  pdiblc1=0.39
+  pdiblc2=0.00056783834
+  pdiblcb=-0.225
+  drout=0.56
+  pscbe1=799985290.0
+  pscbe2=1.0771971e-8
+  pvag=0.0
+  delta=0.01
+  alpha0=0.0
+  alpha1=0.0
+  beta0=30.0
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=1.1890194e-10
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.54561
+  kt2=-0.052484
+  at=10000.0
+  ute=-1.2595
+  ua1=-2.5605e-10
+  ub1=4.9434e-19
+  uc1=8.1951e-12
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.64 pmos
* DC IV MOS Parameters
+  lmin=8e-06 lmax=2.0e-05 wmin=1e-06 wmax=1.26e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.019765+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+  k1=0.49177002
+  k2=-0.002690247
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=55237.817
+  ua=-1.4116341e-9
+  ub=1.370092e-18
+  uc=-3.8916596e-11
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0062318252
+  a0=1.212397
+  keta=0.0066402373
+  a1=0.0
+  a2=0.8
+  ags=0.28815017
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.25245591+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.5589128+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.0017402344
+  pdiblc1=0.39
+  pdiblc2=0.00056783834
+  pdiblcb=-0.225
+  drout=0.56
+  pscbe1=799985290.0
+  pscbe2=1.0771971e-8
+  pvag=0.0
+  delta=0.01
+  alpha0=0.0
+  alpha1=0.0
+  beta0=30.0
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=1.1890194e-10
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.54561
+  kt2=-0.052484
+  at=10000.0
+  ute=-1.2595
+  ua1=-2.5605e-10
+  ub1=4.9434e-19
+  uc1=8.1951e-12
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.65 pmos
* DC IV MOS Parameters
+  lmin=4e-06 lmax=8e-06 wmin=1e-06 wmax=1.26e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.016478161792+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0=-2.63866976917606e-8
+  k1=0.534075464395531 lk1=-3.39627599941981e-7
+  k2=-0.014860639538516 lk2=9.7703765254496e-08 pk2=-2.52435489670724e-29
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=67817.2708528591 lvsat=-0.100987704577306
+  ua=-1.99250034062952e-09 lua=4.6631872093789e-15
+  ub=1.75864839835032e-18 lub=-3.11932610327959e-24
+  uc=-2.3153039787075e-11 luc=-1.26549640114687e-16
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.00400447391202439 lu0=1.78811494116526e-8
+  a0=1.290013307769 la0=-6.23102787373838e-7
+  keta=0.010081996961465 lketa=-2.76304052611251e-8
+  a1=0.0
+  a2=0.8
+  ags=0.23401573324487 lags=4.34590608656943e-7
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.26378896640707+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff=9.09816408392809e-8
+  nfactor={1.1497465565696+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor=3.28478169226432e-6
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-0.0347769002070012 lpclm=2.9315911841939e-07 wpclm=-9.92616735063633e-24 ppclm=1.26217744835362e-29
+  pdiblc1=0.39
+  pdiblc2=9.45014544238799e-05 lpdiblc2=3.79994283736246e-9
+  pdiblcb=-0.225
+  drout=0.56
+  pscbe1=799970497.21407 lpscbe1=0.118756307932927
+  pscbe2=1.20499416283276e-08 lpscbe2=-1.02595328685664e-14
+  pvag=0.0
+  delta=0.01
+  alpha0=0.0
+  alpha1=0.0
+  beta0=30.0
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=4.71295882709498e-11 lagidl=5.76187578412592e-16
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.63053005701 lkt1=6.81737198635594e-7
+  kt2=-0.078406116774 lkt2=2.08102442396271e-7
+  at=-35585.2436945 lat=0.365957789356522 wat=1.38777878078145e-17 pat=-1.05879118406788e-22
+  ute=-2.4573229315 lute=9.61610812020682e-6
+  ua1=-2.44692302305e-09 lua1=1.75883023385691e-14 pua1=3.00926553810506e-36
+  ub1=2.01474435048e-18 lub1=-1.22057878808012e-23
+  uc1=9.70073011147e-11 luc1=-7.12983284802398e-16 wuc1=1.23259516440783e-32 puc1=9.4039548065783e-38
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.66 pmos
* DC IV MOS Parameters
+  lmin=2e-06 lmax=4e-06 wmin=1e-06 wmax=1.26e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.02608082788174+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0=1.22927260857104e-8
+  k1=0.43812032260554 lk1=4.68785597263962e-8
+  k2=0.01293585993148 lk2=-1.42602010526543e-8
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=31904.41993038 lvsat=0.0436688279842283
+  ua=-6.37637714430962e-10 lua=-7.94183190597387e-16
+  ub=8.2357658796972e-19 lub=6.47131928071745e-25
+  uc=-6.42423725923621e-11 luc=3.89576993530151e-17
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.00905878876040002 lu0=-2.47757014582607e-9
+  a0=1.211571334806 la0=-3.0713946158255e-7
+  keta=0.0113714733127004 lketa=-3.28244005301851e-8
+  a1=0.0
+  a2=0.8
+  ags=0.24080219552546 lags=4.07254820028274e-7
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.23789112252874+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff=-1.33345635285058e-8
+  nfactor={2.2722086903828+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.23648231318963e-6
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.160612523 leta0=-3.24706275293724e-7
+  etab=-0.140472581489149 letab=2.83862712567314e-7
+  dsub=0.864198200000001 ldsub=-1.2253066992216e-6
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-0.280678249441224 lpclm=1.28364680231865e-06 ppclm=4.03896783473158e-28
+  pdiblc1=0.39
+  pdiblc2=0.0018722880708822 lpdiblc2=-3.36096032029225e-9
+  pdiblcb=-0.225
+  drout=0.56
+  pscbe1=799999959.720119 lpscbe1=8.16871124698082e-5
+  pscbe2=9.635456366521e-09 lpscbe2=-5.34015207832602e-16
+  pvag=0.0
+  delta=0.01
+  alpha0=-3.091654524078e-12 lalpha0=1.24531473231319e-17
+  alpha1=2.964777003837e-15 lalpha1=-1.19420861941314e-20
+  beta0=57.377838 lbeta0=-0.000110277602929944
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=2.9544148094122e-10 lagidl=-4.24009745520543e-16
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.45145439814 lkt1=-3.9577406384857e-8
+  kt2=-0.00769209472199994 lkt2=-7.67327898609207e-8
+  at=103746.539146 lat=-0.195268959943618
+  ute=0.7665957497 lute=-3.3697976406426e-06 pute=1.61558713389263e-27
+  ua1=4.02151830254e-09 lua1=-8.46650169961149e-15
+  ub1=-2.80235008686e-18 lub1=7.19741070767103e-24 wub1=-1.46936793852786e-39 pub1=-2.80259692864963e-45
+  uc1=-2.23851272804e-10 luc1=5.79431200639238e-16
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.67 pmos
* DC IV MOS Parameters
+  lmin=1e-06 lmax=2e-06 wmin=1e-06 wmax=1.26e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.02950288021532+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0=1.92326071535865e-8
+  k1=0.469075083613521 lk1=-1.58973241406559e-8
+  k2=0.004272102579488 lk2=3.30979489209729e-9
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=78753.615529692 lvsat=-0.051340778500829
+  ua=-1.29898347783292e-09 lua=5.47018081432629e-16
+  ub=1.32344821524624e-18 lub=-3.66601733585513e-25
+  uc=-4.1282867652764e-11 luc=-7.60390115043052e-18
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.00700268214039999 lu0=1.69218940625448e-9
+  a0=1.582204237572 la0=-1.05877854079717e-6
+  keta=0.0291366334094596 lketa=-6.88519320244916e-08 pketa=6.31088724176809e-30
+  a1=0.0
+  a2=0.8
+  ags=-0.374332360800441 lags=1.65474031864252e-6
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.2466516868904+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff=4.43175587016839e-9
+  nfactor={1.5005339170744+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor=3.28464866982522e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=-0.0812250460000001 leta0=1.65737412587448e-07 weta0=-3.30872245021211e-24 peta0=3.07655753036195e-29
+  etab=0.00618191897829788 letab=-1.35508545266625e-08 wetab=-8.27180612553028e-25 petab=1.57772181044202e-30
+  dsub=-0.0483964000000001 ldsub=6.254241984432e-7
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.332664105388719 lpclm=3.97958668317801e-8
+  pdiblc1=0.39797787563196 lpdiblc1=-1.61790360471074e-8
+  pdiblc2=0.000215
+  pdiblcb=-0.4305976 lpdiblcb=4.169494656288e-07 wpdiblcb=4.2351647362715e-22
+  drout=0.1989163366336 ldrout=7.32273336303098e-7
+  pscbe1=800000000.0
+  pscbe2=1.03613408527e-08 lpscbe2=-2.00610023518976e-15
+  pvag=0.0
+  delta=0.01
+  alpha0=-9.66154909518441e-11 lalpha0=2.02118365312604e-16 walpha0=4.93038065763132e-32 palpha0=2.93873587705572e-38
+  alpha1=-1.02804729554008e-10 lalpha1=2.08480828324765e-16 walpha1=-1.93375403478631e-32 palpha1=5.68633912773262e-38
+  beta0=-3.06618412128561 lbeta0=1.23021486037577e-5
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=7.521286103248e-11 lagidl=2.26112529109428e-17
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.42689323608076 lkt1=-8.9387148307051e-8
+  kt2=-0.02666911067692 lkt2=-3.82476292285345e-8
+  at=-8464.61082126801 lat=0.0322939056562017
+  ute=-0.588317398578001 lute=-6.22050034892599e-7
+  ua1=-6.371834778916e-11 lua1=-1.81690795583757e-16
+  ub1=1.02092658491736e-18 lub1=-5.56148503373387e-25
+  uc1=7.6699274718912e-11 luc1=-3.00817031306568e-17
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=2.745e-6
+  sbref=2.74e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.68 pmos
* DC IV MOS Parameters
+  lmin=5e-07 lmax=1e-06 wmin=1e-06 wmax=1.26e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.0714786231704+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0=6.23831672024935e-8
+  k1=0.394999825372881 lk1=6.02511524276241e-8
+  k2=0.0222744113979824 lk2=-1.51963625456091e-8
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=-1808.81819138397 lvsat=0.0314764366152325
+  ua=-3.76203156092561e-10 lua=-4.01589015952602e-16
+  ub=7.0272563813328e-19 lub=2.71493627015686e-25
+  uc=-7.7067301765592e-11 luc=2.91820677043474e-17
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.01061399245552 lu0=-2.02019426196509e-9
+  a0=-0.0634326948480002 la0=6.32916478087406e-7
+  keta=-0.042575756671448 lketa=4.86754443000049e-9
+  a1=0.0
+  a2=0.8
+  ags=1.1537197626112 lags=8.39210724008375e-8
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.24175577993144+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff=-6.01177732758859e-10
+  nfactor={1.7372633632936+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor=8.5109837022539e-8
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=-0.35295016 leta0=4.4506756907808e-7
+  etab=-0.01438523215 letab=7.5919300274142e-9
+  dsub=0.81616026316352 ldsub=-2.63329676608941e-07 wdsub=-8.470329472543e-22
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.10226051009128 lpclm=2.76647997954405e-7
+  pdiblc1=0.62203846997568 lpdiblc1=-2.46510638305319e-7
+  pdiblc2=-0.000119947403386 lpdiblc2=3.44321911311968e-10
+  pdiblcb=-0.025
+  drout=0.817537886732799 ldrout=9.63378062597227e-8
+  pscbe1=800000000.0
+  pscbe2=7.45177980621521e-09 lpscbe2=9.84893605864053e-16
+  pvag=0.0
+  delta=0.01
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=8.7628431869944 lbeta0=1.42050479173602e-7
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=8.63250305572001e-11 lagidl=1.11880759855651e-17
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.51953498759848 lkt1=5.84746055214585e-9
+  kt2=-0.0730491064621599 lkt2=9.43044987874294e-9
+  at=-21453.665385464 lat=0.0456464978795404 pat=1.32348898008484e-23
+  ute=-2.199567016764 lute=1.03429523760719e-6
+  ua1=-1.08172939594168e-09 lua1=8.64812345784455e-16 pua1=3.76158192263132e-37
+  ub1=4.0432222584528e-19 lub1=7.77133785004025e-26
+  uc1=7.1847125458176e-11 luc1=-2.50937519164114e-17
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.745e-6
+  sbref=1.74e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.69 pmos
* DC IV MOS Parameters
+  lmin=2.5e-07 lmax=5e-07 wmin=1e-06 wmax=1.26e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.934619631504001+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0=-9.87673808946638e-9
+  k1=0.43001994765856 lk1=4.17609481022523e-8
+  k2=0.0102484393695712 lk2=-8.84679362627236e-9
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=-74155.8939940799 lvsat=0.0696748244741463
+  ua=-6.24896580150402e-10 lua=-2.70281872371151e-16
+  ub=8.54553983596802e-19 lub=1.91330082551093e-25
+  uc=-4.6095809352361e-11 luc=1.28294913680704e-17
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.008823486124 lu0=-1.07482840499851e-9
+  a0=1.49467176688 la0=-1.89743980451438e-7
+  keta=-0.0593620093695648 lketa=1.37304844195738e-8
+  a1=0.0
+  a2=1.10720647359648 la2=-1.62201331581259e-7
+  ags=2.30325973754048 lags=-5.23022239882123e-7
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.19564020951728+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff=-2.49496455245904e-8
+  nfactor={1.9273171671088+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor=-1.52362907462407e-8
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.49
+  etab=5.62972999999999e-05 letab=-3.30242238324e-11 wetab=-1.29246970711411e-26 petab=-6.16297582203915e-33
+  dsub=-0.0279335847931197 ldsub=1.8234174598599e-7
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.61407741662336 lpclm=6.41481310834537e-9
+  pdiblc1=-0.18599373358432 lpdiblc1=1.80120668787918e-07 ppdiblc1=5.04870979341448e-29
+  pdiblc2=-0.011182490884396 lpdiblc2=6.18521211876348e-09 wpdiblc2=8.27180612553028e-25 ppdiblc2=-1.18329135783152e-30
+  pdiblcb=0.1973904 lpdiblcb=-1.174194625152e-07 wpdiblcb=-5.29395592033938e-23
+  drout=1.63194501654032 ldrout=-3.3365938539309e-7
+  pscbe1=800079104.265282 lpscbe1=-0.0417661028168368
+  pscbe2=9.4366626002032e-09 lpscbe2=-6.31006907680859e-17
+  pvag=0.0
+  delta=0.01
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=8.7413550381728 lbeta0=1.53395963893621e-7
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-5.619411557624e-10 lagidl=3.53464843168078e-16 wagidl=1.97215226305253e-31 pagidl=-4.70197740328915e-38
+  bgidl=691592551.526402 lbgidl=162.835431904679
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.50444585328 lkt1=-2.11942129839932e-9
+  kt2=-0.096992947392 lkt2=2.20725105636073e-8
+  at=63269.802688 lat=0.000913523418368256
+  ute=-0.30218766272 lute=3.25017072242073e-8
+  ua1=7.2708366384e-10 lua1=-9.02192440235539e-17
+  ub1=6.7661571952e-19 lub1=-6.60543186379256e-26
+  uc1=5.072625803232e-11 luc1=-1.39421873659686e-17
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.245e-6
+  sbref=1.24e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.70 pmos
* DC IV MOS Parameters
+  lmin=1.8e-07 lmax=2.5e-07 wmin=1e-06 wmax=1.26e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.899843113485716+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0=-1.9544192780334e-8
+  k1=-1.04921174370343 lk1=4.52969607520589e-7
+  k2=0.582611608243943 lk2=-1.67956886215321e-07 wk2=-1.58818677610181e-22 pk2=5.04870979341448e-29
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=398287.511750286 lvsat=-0.0616587730019185
+  ua=7.16529660737141e-10 lua=-6.43182270222996e-16
+  ub=-3.54747312851425e-19 lub=5.27501331348142e-25
+  uc=-4.606963774268e-13 luc=1.43477582394365e-19 wuc=1.92592994438724e-34
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0109018618662857 lu0=-1.65259192084504e-9
+  a0=-0.00465887600000059 la0=2.27051946301488e-7
+  keta=-0.120180916787726 lketa=3.06374108549335e-08 wketa=5.29395592033938e-23 pketa=6.31088724176809e-30
+  a1=0.0
+  a2=0.0392201759994286 la2=1.34686043315151e-7
+  ags=-2.03898102803886 lags=6.84068586059746e-7
+  b0=0.0
+  b1=-6.26145615844572e-24 lb1=1.74060967457401e-30
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.168675364554856+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff=-3.24455488460044e-8
+  nfactor={0.997080565485717+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor=2.43358321665759e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=1.31788295248057 leta0=-2.30141526194169e-7
+  etab=0.0935091143547428 letab=-2.60117859312463e-08 wetab=-1.24077091882954e-23 petab=2.26797510251041e-30
+  dsub=1.693234542632 ldsub=-2.96122339420664e-7
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.682002296978858 lpclm=-1.24674885319186e-8
+  pdiblc1=1.382172001224 lpdiblc1=-2.55810587499977e-7
+  pdiblc2=0.03707351932236 lpdiblc2=-7.22937964659221e-9
+  pdiblcb=-0.670688571428571 lpdiblcb=1.23896074594286e-7
+  drout=-1.256946487644 ldrout=4.694177860721e-7
+  pscbe1=799717484.766857 lpscbe1=0.0587597783110141
+  pscbe2=8.67880867706288e-09 lpscbe2=1.47573605617857e-16
+  pvag=0.0
+  delta=0.01
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=10.7811435185828 lbeta0=-4.13640756198613e-7
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=2.52075921657143e-09 lagidl=-5.03488867936258e-16
+  bgidl=2092679862.27428 lbgidl=-226.650027435504
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.231654635885715 lkt1=-7.79521062394021e-8
+  kt2=0.286688501485714 lkt2=-8.45863280470107e-08 wkt2=5.29395592033938e-23
+  at=88578.9579428572 lat=-0.00612211803261897
+  ute=-0.0934878668571431 lute=-2.55143316281167e-8
+  ua1=1.15141565028571e-09 lua1=-2.08178444271625e-16
+  ub1=4.39e-19
+  uc1=-5.24083598285714e-13 luc1=3.0479260324025e-19
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.1e-6
+  sbref=1.1e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.71 pmos
* DC IV MOS Parameters
+  lmin=1.5e-07 lmax=1.8e-07 wmin=1e-06 wmax=1.26e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.788718570808747+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0=-4.26567641626294e-08 wvth0=1.96024078967603e-10 pvth0=-4.07706561370577e-17
+  k1=4.11830102617436 lk1=-6.21811038460751e-07 wk1=-5.10199991329752e-06 pk1=1.06115475796693e-12
+  k2=-1.38668350242437 lk2=2.41632865262361e-07 wk2=1.98275275498596e-06 pk2=-4.1238878000402e-13
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=-459891.739157119 lvsat=0.116832213035811 wvsat=0.825459720823284 pvsat=-1.71685716414593e-7
+  ua=-5.09677744853903e-09 lua=5.65915848821138e-16 wua=3.95559789295204e-15 pua=-8.22716894559309e-22
+  ub=3.63535079134925e-18 lub=-3.02391193148348e-25 wub=-2.74262889573271e-24 pub=5.70433898765656e-31
+  uc=2.22165827457476e-12 luc=-4.14419996966135e-19 wuc=-1.98048923694266e-18 puc=4.11917995413231e-25
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=-0.00492412921573533 lu0=1.63902431232236e-09 wu0=1.02260161310072e-08 pu0=-2.12688864305593e-15
+  a0=-2.08228480125189 la0=6.59173207242779e-07 wa0=5.23376113842361e-06 pa0=-1.08855951165845e-12
+  keta=0.761151985656444 lketa=-1.52669256858625e-07 wketa=-5.62536765411136e-07 pketa=1.17000896764331e-13
+  a1=0.0
+  a2=2.40751338627852 la2=-3.57890524904377e-07 wa2=-3.52379661186828e-06 pa2=7.32907409709259e-13
+  ags=1.25
+  b0=0.0
+  b1=1.46100643697067e-23 lb1=-2.60041613703535e-30
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={0.994569654925066+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff=-2.74386553957595e-07 wvoff=-1.60935348781818e-06 pvoff=3.34726213224328e-13
+  nfactor={-9.55756180582907+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor=2.43859727919078e-06 wnfactor=1.46780310022279e-05 pnfactor=-3.05285431209138e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=3.17607718361169 leta0=-6.16623627938668e-07 weta0=-3.68688528515757e-06 peta0=7.66827896689352e-13
+  etab=0.199797492392715 letab=-4.81184931026082e-08 wetab=-4.12450260063194e-07 petab=8.57847046900236e-14
+  dsub=0.467176730191369 ldsub=-4.11170271267622e-08 wdsub=-1.76100751651244e-07 pdsub=3.66268431344385e-14
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-2.99898054296121 lpclm=7.53132770381538e-07 wpclm=4.55215461206512e-06 ppclm=-9.46793533454201e-13
+  pdiblc1=-2.54577407474361 lpdiblc1=5.61155060948375e-07 wpdiblc1=3.43465214164761e-06 ppdiblc1=-7.14366429637004e-13
+  pdiblc2=-0.0496171610450667 lpdiblc2=1.08012415816681e-08 wpdiblc2=6.21929459819132e-08 ppdiblc2=-1.29353864488862e-14
+  pdiblcb=3.79591210725848 lpdiblcb=-8.05103267364477e-07 wpdiblcb=-4.25269383350002e-06 ppdiblcb=8.84509285042002e-13
+  drout=1.0
+  pscbe1=800000000.0
+  pscbe2=1.50686260347976e-08 lpscbe2=-1.18143172698268e-15 wpscbe2=-5.52596359163528e-15 ppscbe2=1.14933411549704e-21
+  pvag=0.0
+  delta=0.01
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=-1.5848823221769 lbeta0=2.15834422636934e-06 wbeta0=1.92355824372214e-05 pbeta0=-4.00077031995282e-12
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=9.98778569869926e-09 lagidl=-2.05654077190107e-15 wagidl=-1.4536654515994e-14 pagidl=3.02344969947256e-21
+  bgidl=1020475725.30667 lbgidl=-3.64443339588342
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=1.36130201414738 lkt1=-4.09267973966487e-07 wkt1=-1.91059069082956e-06 pkt1=3.97379936604259e-13
+  kt2=-0.12
+  at=-563008.159389326 lat=0.129400183327067 wat=0.835426621125335 pat=-1.73758712074616e-7
+  ute=-0.238289841333334 lute=4.60274143923742e-9
+  ua1=-1.73814038436491e-09 lua1=3.92814536263289e-16 wua1=2.11173939929144e-15 pua1=-4.39216454179828e-22
+  ub1=8.54839297333334e-19 lub1=-8.64895837737652e-26
+  uc1=2.28016756041765e-12 luc1=-2.7845798675616e-19 wuc1=-4.23580031211806e-17 puc1=8.80995635316812e-24
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.04e-6
+  sbref=1.04e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.72 pmos
* DC IV MOS Parameters
+  lmin=2.0e-05 lmax=1.0e-04 wmin=8.4e-07 wmax=1.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.019765+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+  k1=0.49177002
+  k2=-0.002690247
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=55237.817
+  ua=-1.4116341e-9
+  ub=1.370092e-18
+  uc=-3.8916596e-11
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0062318252
+  a0=1.212397
+  keta=0.0066402373
+  a1=0.0
+  a2=0.8
+  ags=0.28815017
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.25245591+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.5589128+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.0017402344
+  pdiblc1=0.39
+  pdiblc2=0.00056783834
+  pdiblcb=-0.225
+  drout=0.56
+  pscbe1=799985290.0
+  pscbe2=1.0771971e-8
+  pvag=0.0
+  delta=0.01
+  alpha0=0.0
+  alpha1=0.0
+  beta0=30.0
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=1.1890194e-10
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.54561
+  kt2=-0.052484
+  at=10000.0
+  ute=-1.2595
+  ua1=-2.5605e-10
+  ub1=4.9434e-19
+  uc1=8.1951e-12
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.73 pmos
* DC IV MOS Parameters
+  lmin=8e-06 lmax=2.0e-05 wmin=8.4e-07 wmax=1.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.019765+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+  k1=0.49177002
+  k2=-0.002690247
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=55237.817
+  ua=-1.4116341e-9
+  ub=1.370092e-18
+  uc=-3.8916596e-11
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0062318252
+  a0=1.212397
+  keta=0.0066402373
+  a1=0.0
+  a2=0.8
+  ags=0.28815017
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.25245591+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.5589128+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.0017402344
+  pdiblc1=0.39
+  pdiblc2=0.00056783834
+  pdiblcb=-0.225
+  drout=0.56
+  pscbe1=799985290.0
+  pscbe2=1.0771971e-8
+  pvag=0.0
+  delta=0.01
+  alpha0=0.0
+  alpha1=0.0
+  beta0=30.0
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=1.1890194e-10
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.54561
+  kt2=-0.052484
+  at=10000.0
+  ute=-1.2595
+  ua1=-2.5605e-10
+  ub1=4.9434e-19
+  uc1=8.1951e-12
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.74 pmos
* DC IV MOS Parameters
+  lmin=4e-06 lmax=8e-06 wmin=8.4e-07 wmax=1.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.016478161792+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0=-2.63866976917606e-8
+  k1=0.53407546439553 lk1=-3.39627599941978e-7
+  k2=-0.014860639538516 lk2=9.77037652544961e-08 wk2=-6.61744490042422e-24 pk2=5.04870979341448e-29
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=67817.2708528591 lvsat=-0.100987704577306
+  ua=-1.99250034062952e-09 lua=4.66318720937891e-15
+  ub=1.75864839835032e-18 lub=-3.11932610327959e-24
+  uc=-2.3153039787075e-11 luc=-1.26549640114687e-16
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.00400447391202441 lu0=1.78811494116526e-8
+  a0=1.290013307769 la0=-6.23102787373838e-7
+  keta=0.010081996961465 lketa=-2.7630405261125e-8
+  a1=0.0
+  a2=0.8
+  ags=0.23401573324487 lags=4.34590608656944e-7
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.26378896640707+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff=9.09816408392809e-8
+  nfactor={1.1497465565696+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor=3.28478169226435e-6
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-0.0347769002070012 lpclm=2.93159118419391e-07 wpclm=3.30872245021211e-24 ppclm=8.83524213847533e-29
+  pdiblc1=0.39
+  pdiblc2=9.45014544238799e-05 lpdiblc2=3.79994283736246e-9
+  pdiblcb=-0.225
+  drout=0.56
+  pscbe1=799970497.214071 lpscbe1=0.118756307929289
+  pscbe2=1.20499416283276e-08 lpscbe2=-1.02595328685664e-14
+  pvag=0.0
+  delta=0.01
+  alpha0=0.0
+  alpha1=0.0
+  beta0=30.0
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=4.712958827095e-11 lagidl=5.76187578412593e-16
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.63053005701 lkt1=6.81737198635594e-7
+  kt2=-0.078406116774 lkt2=2.08102442396271e-7
+  at=-35585.2436945 lat=0.365957789356522 wat=-1.38777878078145e-17 pat=-5.29395592033938e-23
+  ute=-2.4573229315 lute=9.61610812020682e-6
+  ua1=-2.44692302305e-09 lua1=1.75883023385691e-14
+  ub1=2.01474435048e-18 lub1=-1.22057878808012e-23 wub1=7.3468396926393e-40 pub1=5.60519385729927e-45
+  uc1=9.70073011147001e-11 luc1=-7.12983284802399e-16 wuc1=-1.23259516440783e-32 puc1=-3.29138418230241e-37
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.75 pmos
* DC IV MOS Parameters
+  lmin=2e-06 lmax=4e-06 wmin=8.4e-07 wmax=1.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.02608082788174+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0=1.22927260857138e-8
+  k1=0.43812032260554 lk1=4.68785597263962e-8
+  k2=0.01293585993148 lk2=-1.42602010526543e-8
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=31904.41993038 lvsat=0.0436688279842286
+  ua=-6.37637714430961e-10 lua=-7.94183190597387e-16
+  ub=8.23576587969721e-19 lub=6.47131928071748e-25
+  uc=-6.42423725923619e-11 luc=3.89576993530149e-17
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.00905878876040002 lu0=-2.47757014582607e-9
+  a0=1.211571334806 la0=-3.07139461582554e-7
+  keta=0.0113714733127004 lketa=-3.28244005301851e-8
+  a1=0.0
+  a2=0.8
+  ags=0.24080219552546 lags=4.07254820028274e-7
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.23789112252874+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff=-1.3334563528505e-8
+  nfactor={2.2722086903828+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.23648231318964e-6
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.160612523 leta0=-3.24706275293724e-7
+  etab=-0.140472581489149 letab=2.83862712567314e-7
+  dsub=0.8641982 ldsub=-1.2253066992216e-6
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-0.280678249441224 lpclm=1.28364680231865e-06 wpclm=-1.05879118406788e-22 ppclm=-3.02922587604869e-28
+  pdiblc1=0.39
+  pdiblc2=0.0018722880708822 lpdiblc2=-3.36096032029225e-9
+  pdiblcb=-0.225
+  drout=0.56
+  pscbe1=799999959.720119 lpscbe1=8.16871142887976e-5
+  pscbe2=9.635456366521e-09 lpscbe2=-5.34015207832627e-16
+  pvag=0.0
+  delta=0.01
+  alpha0=-3.091654524078e-12 lalpha0=1.24531473231319e-17
+  alpha1=2.964777003837e-15 lalpha1=-1.19420861941314e-20
+  beta0=57.377838 lbeta0=-0.000110277602929944
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=2.9544148094122e-10 lagidl=-4.24009745520542e-16
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.45145439814 lkt1=-3.9577406384857e-8
+  kt2=-0.007692094722 lkt2=-7.67327898609206e-8
+  at=103746.539146 lat=-0.195268959943618
+  ute=0.7665957497 lute=-3.3697976406426e-06 wute=-4.2351647362715e-22 pute=-1.41363874215605e-27
+  ua1=4.02151830254e-09 lua1=-8.46650169961149e-15
+  ub1=-2.80235008686e-18 lub1=7.19741070767104e-24 wub1=1.46936793852786e-39
+  uc1=-2.23851272804e-10 luc1=5.79431200639238e-16 wuc1=-9.86076131526265e-32 puc1=1.88079096131566e-37
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.76 pmos
* DC IV MOS Parameters
+  lmin=1e-06 lmax=2e-06 wmin=8.4e-07 wmax=1.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.02950288021532+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0=1.92326071535865e-8
+  k1=0.46907508361352 lk1=-1.58973241406542e-8
+  k2=0.004272102579488 lk2=3.30979489209729e-9
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=78753.615529692 lvsat=-0.0513407785008291
+  ua=-1.29898347783292e-09 lua=5.47018081432629e-16
+  ub=1.32344821524624e-18 lub=-3.66601733585511e-25
+  uc=-4.1282867652764e-11 luc=-7.60390115043042e-18
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.00700268214040001 lu0=1.69218940625449e-9
+  a0=1.582204237572 la0=-1.05877854079716e-6
+  keta=0.0291366334094596 lketa=-6.88519320244915e-08 wketa=6.61744490042422e-24 pketa=-6.31088724176809e-30
+  a1=0.0
+  a2=0.8
+  ags=-0.374332360800441 lags=1.65474031864252e-6
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.2466516868904+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff=4.43175587016839e-9
+  nfactor={1.5005339170744+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor=3.28464866982522e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=-0.081225046 leta0=1.65737412587448e-07 weta0=-1.73707928636136e-23 peta0=-1.65660790096412e-29
+  etab=0.00618191897829788 letab=-1.35508545266625e-08 wetab=-2.48154183765908e-24 petab=6.31088724176809e-30
+  dsub=-0.0483964000000001 ldsub=6.25424198443201e-7
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.332664105388719 lpclm=3.97958668317805e-8
+  pdiblc1=0.39797787563196 lpdiblc1=-1.61790360471074e-8
+  pdiblc2=0.000215
+  pdiblcb=-0.4305976 lpdiblcb=4.169494656288e-7
+  drout=0.1989163366336 ldrout=7.322733363031e-7
+  pscbe1=800000000.0
+  pscbe2=1.03613408527e-08 lpscbe2=-2.00610023518978e-15
+  pvag=0.0
+  delta=0.01
+  alpha0=-9.6615490951844e-11 lalpha0=2.02118365312604e-16 walpha0=1.23259516440783e-32 palpha0=6.46521892952258e-38
+  alpha1=-1.02804729554008e-10 lalpha1=2.08480828324765e-16 walpha1=2.60301469046087e-32 palpha1=-2.28957371358892e-38
+  beta0=-3.0661841212856 lbeta0=1.23021486037577e-05 pbeta0=-6.46234853557053e-27
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=7.52128610324799e-11 lagidl=2.26112529109428e-17
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.426893236080759 lkt1=-8.9387148307051e-8
+  kt2=-0.02666911067692 lkt2=-3.82476292285343e-8
+  at=-8464.61082126801 lat=0.0322939056562017 pat=1.32348898008484e-23
+  ute=-0.588317398578001 lute=-6.22050034892598e-7
+  ua1=-6.371834778916e-11 lua1=-1.81690795583757e-16
+  ub1=1.02092658491736e-18 lub1=-5.56148503373388e-25
+  uc1=7.66992747189121e-11 luc1=-3.00817031306569e-17
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=2.745e-6
+  sbref=2.74e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.77 pmos
* DC IV MOS Parameters
+  lmin=5e-07 lmax=1e-06 wmin=8.4e-07 wmax=1.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.0714786231704+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0=6.23831672024926e-8
+  k1=0.39499982537288 lk1=6.02511524276237e-8
+  k2=0.0222744113979824 lk2=-1.51963625456091e-08 pk2=6.31088724176809e-30
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=-1808.81819138397 lvsat=0.0314764366152325
+  ua=-3.7620315609256e-10 lua=-4.015890159526e-16
+  ub=7.0272563813328e-19 lub=2.71493627015684e-25
+  uc=-7.7067301765592e-11 luc=2.91820677043474e-17
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.01061399245552 lu0=-2.02019426196509e-9
+  a0=-0.0634326948479993 la0=6.32916478087406e-7
+  keta=-0.042575756671448 lketa=4.86754443000046e-9
+  a1=0.0
+  a2=0.8
+  ags=1.1537197626112 lags=8.39210724008375e-8
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.24175577993144+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff=-6.01177732758859e-10
+  nfactor={1.7372633632936+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor=8.5109837022539e-8
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=-0.35295016 leta0=4.4506756907808e-07 peta0=1.0097419586829e-28
+  etab=-0.01438523215 letab=7.59193002741421e-9
+  dsub=0.81616026316352 ldsub=-2.63329676608941e-7
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.10226051009128 lpclm=2.76647997954406e-7
+  pdiblc1=0.62203846997568 lpdiblc1=-2.46510638305319e-7
+  pdiblc2=-0.000119947403386 lpdiblc2=3.44321911311968e-10
+  pdiblcb=-0.025
+  drout=0.817537886732801 ldrout=9.63378062597227e-8
+  pscbe1=800000000.0
+  pscbe2=7.4517798062152e-09 lpscbe2=9.84893605864059e-16
+  pvag=0.0
+  delta=0.01
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=8.76284318699442 lbeta0=1.42050479173596e-7
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=8.63250305572001e-11 lagidl=1.11880759855651e-17
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.51953498759848 lkt1=5.84746055214585e-9
+  kt2=-0.07304910646216 lkt2=9.43044987874294e-9
+  at=-21453.665385464 lat=0.0456464978795403
+  ute=-2.199567016764 lute=1.03429523760719e-6
+  ua1=-1.08172939594168e-09 lua1=8.64812345784456e-16 pua1=-1.88079096131566e-37
+  ub1=4.04322225845279e-19 lub1=7.77133785004025e-26
+  uc1=7.1847125458176e-11 luc1=-2.50937519164114e-17
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.745e-6
+  sbref=1.74e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.78 pmos
* DC IV MOS Parameters
+  lmin=2.5e-07 lmax=5e-07 wmin=8.4e-07 wmax=1.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.934619631503999+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0=-9.87673808946595e-9
+  k1=0.430019947658559 lk1=4.17609481022523e-8
+  k2=0.0102484393695712 lk2=-8.84679362627236e-09 pk2=-3.15544362088405e-30
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=-74155.8939940801 lvsat=0.0696748244741463 pvsat=2.64697796016969e-23
+  ua=-6.24896580150399e-10 lua=-2.70281872371151e-16
+  ub=8.54553983596799e-19 lub=1.91330082551092e-25
+  uc=-4.60958093523609e-11 luc=1.28294913680704e-17
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.008823486124 lu0=-1.07482840499851e-9
+  a0=1.49467176688 la0=-1.89743980451438e-7
+  keta=-0.0593620093695648 lketa=1.37304844195738e-08 pketa=1.26217744835362e-29
+  a1=0.0
+  a2=1.10720647359648 la2=-1.62201331581258e-7
+  ags=2.30325973754048 lags=-5.23022239882123e-7
+  b0=0.0
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.19564020951728+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff=-2.49496455245903e-8
+  nfactor={1.9273171671088+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor=-1.52362907462415e-8
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.49
+  etab=5.62973e-05 letab=-3.30242238324e-11 wetab=1.29246970711411e-26 petab=-3.08148791101958e-33
+  dsub=-0.0279335847931206 ldsub=1.8234174598599e-7
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.614077416623358 lpclm=6.41481310834558e-9
+  pdiblc1=-0.18599373358432 lpdiblc1=1.80120668787918e-7
+  pdiblc2=-0.011182490884396 lpdiblc2=6.18521211876347e-09 wpdiblc2=-8.27180612553028e-25 ppdiblc2=9.86076131526265e-31
+  pdiblcb=0.1973904 lpdiblcb=-1.174194625152e-07 wpdiblcb=1.05879118406788e-22 ppdiblcb=-3.78653234506086e-29
+  drout=1.63194501654032 ldrout=-3.3365938539309e-7
+  pscbe1=800079104.265278 lpscbe1=-0.0417661028168368
+  pscbe2=9.43666260020318e-09 lpscbe2=-6.31006907680828e-17
+  pvag=0.0
+  delta=0.01
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=8.74135503817278 lbeta0=1.53395963893621e-7
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-5.619411557624e-10 lagidl=3.53464843168078e-16 pagidl=9.4039548065783e-38
+  bgidl=691592551.526398 lbgidl=162.835431904679
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.504445853279999 lkt1=-2.11942129839953e-9
+  kt2=-0.0969929473919998 lkt2=2.20725105636073e-8
+  at=63269.8026879999 lat=0.000913523418368284
+  ute=-0.30218766272 lute=3.25017072242073e-8
+  ua1=7.27083663839999e-10 lua1=-9.02192440235541e-17
+  ub1=6.7661571952e-19 lub1=-6.60543186379258e-26 wub1=-7.3468396926393e-40
+  uc1=5.072625803232e-11 luc1=-1.39421873659686e-17
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.245e-6
+  sbref=1.24e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.79 pmos
* DC IV MOS Parameters
+  lmin=1.8e-07 lmax=2.5e-07 wmin=8.4e-07 wmax=1.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.899843113485709+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0=-1.95441927803331e-8
+  k1=-1.04921174370343 lk1=4.52969607520589e-7
+  k2=0.582611608243943 lk2=-1.67956886215321e-7
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=398287.511750286 lvsat=-0.0616587730019185
+  ua=7.16529660737154e-10 lua=-6.43182270222999e-16
+  ub=-3.54747312851432e-19 lub=5.27501331348143e-25
+  uc=-4.606963774268e-13 luc=1.43477582394365e-19 puc=4.59177480789956e-41
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0109018618662857 lu0=-1.65259192084503e-9
+  a0=-0.00465887600000059 la0=2.27051946301489e-7
+  keta=-0.120180916787726 lketa=3.06374108549335e-08 wketa=2.64697796016969e-23 pketa=6.31088724176809e-30
+  a1=0.0
+  a2=0.0392201759994251 la2=1.34686043315151e-7
+  ags=-2.03898102803886 lags=6.84068586059746e-7
+  b0=0.0
+  b1=-6.26145615844572e-24 lb1=1.74060967457401e-30
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.168675364554855+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff=-3.24455488460046e-8
+  nfactor={0.99708056548571+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor=2.43358321665758e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=1.31788295248057 leta0=-2.30141526194169e-7
+  etab=0.0935091143547429 letab=-2.60117859312463e-08 wetab=4.54949336904165e-24 petab=1.17343059651626e-29
+  dsub=1.693234542632 ldsub=-2.96122339420665e-07 wdsub=1.6940658945086e-21
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.682002296978856 lpclm=-1.24674885319186e-8
+  pdiblc1=1.382172001224 lpdiblc1=-2.55810587499977e-7
+  pdiblc2=0.03707351932236 lpdiblc2=-7.22937964659221e-9
+  pdiblcb=-0.67068857142857 lpdiblcb=1.23896074594286e-7
+  drout=-1.256946487644 ldrout=4.694177860721e-7
+  pscbe1=799717484.766857 lpscbe1=0.0587597783110141
+  pscbe2=8.67880867706283e-09 lpscbe2=1.47573605617844e-16
+  pvag=0.0
+  delta=0.01
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=10.7811435185828 lbeta0=-4.13640756198613e-7
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=2.52075921657142e-09 lagidl=-5.03488867936258e-16
+  bgidl=2092679862.27428 lbgidl=-226.650027435504
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.231654635885713 lkt1=-7.79521062394021e-8
+  kt2=0.286688501485715 lkt2=-8.45863280470108e-08 wkt2=5.29395592033938e-23
+  at=88578.9579428567 lat=-0.00612211803261897
+  ute=-0.0934878668571422 lute=-2.55143316281165e-8
+  ua1=1.15141565028571e-09 lua1=-2.08178444271625e-16
+  ub1=4.39e-19
+  uc1=-5.24083598285719e-13 luc1=3.0479260324025e-19
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.1e-6
+  sbref=1.1e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.80 pmos
* DC IV MOS Parameters
+  lmin=1.5e-07 lmax=1.8e-07 wmin=8.4e-07 wmax=1.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.749710940395602+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0=-5.07698831969992e-08 wvth0=-3.8241790670624e-08 pvth0=7.9538335580017e-15
+  k1=-5.85428844906348 lk1=1.45236790131502e-06 wk1=4.72491196940394e-06 pk1=-9.82724990692385e-13
+  k2=2.23290028267025 lk2=-5.111971270319e-07 wk2=-1.58395687409276e-06 pk2=3.29444022328805e-13
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=343925.411286352 lvsat=-0.0503521084506259 wvsat=0.0333845705500604 pvsat=-6.94359005956604e-9
+  ua=-1.61065089243855e-09 lua=-1.59156641329088e-16 wua=5.20395976357762e-16 pua=-1.08236118330697e-22
+  ub=2.52206562900939e-18 lub=-7.08412388036046e-26 wub=-1.64560638038729e-24 pub=3.4226637984399e-31
+  uc=-2.16467088758533e-12 luc=4.97883832813219e-19 wuc=2.34176530608242e-18 puc=-4.87059082481471e-25
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0056713973312255 lu0=-5.64718063126932e-10 wu0=-2.1473308326092e-10 pu0=4.46619045212702e-17
+  a0=13.0631229413606 la0=-2.4908898583277e-06 wa0=-9.69040551696633e-06 pa0=2.01548806266279e-12
+  keta=3.15941242683372 lketa=-6.51478649498204e-07 wketa=-2.92576389771578e-06 pketa=6.08523781558111e-13
+  a1=0.0
+  a2=-1.16852122396933 la2=3.85881761611854e-7
+  ags=-19.2893357426319 lags=4.27193536243852e-06 wags=2.02393012339707e-05 pags=-4.20953178505109e-12
+  b0=0.0
+  b1=1.46100643697067e-23 lb1=-2.60041613703535e-30
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={0.75275727111028+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff=-2.24092479872725e-07 wvoff=-1.37107345094369e-06 pvoff=2.85166824914875e-13
+  nfactor={-5.41969190609261+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor=1.57796999448439e-06 wnfactor=1.06006062784128e-05 pnfactor=-2.20479889863452e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=1.24878542050382 leta0=-2.15770068713389e-07 weta0=-1.78774701466683e-06 peta0=3.71829926086525e-13
+  etab=-1.48931911887505 letab=3.03197492641753e-07 wetab=1.2519920735705e-06 petab=-2.60399327397781e-13
+  dsub=0.0959968937635232 ldsub=3.6083924692192e-08 wdsub=1.89656963962031e-07 pdsub=-3.94463726205349e-14
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-3.53376297321431 lpclm=8.64361098485018e-07 wpclm=5.07912504753356e-06 ppclm=-1.05639706038641e-12
+  pdiblc1=0.939794556353335 lpdiblc1=-1.63801387496217e-7
+  pdiblc2=0.01349775500756 lpdiblc2=-2.32590357828559e-9
+  pdiblcb=-0.519825152991825 lpdiblcb=9.25182939204638e-8
+  drout=1.0
+  pscbe1=-147376080.210926 lpscbe1=197.042856170909 wpscbe1=933.536999906417 ppscbe1=-0.000194164493536536
+  pscbe2=-8.12769301278432e-09 lpscbe2=3.64312427908578e-15 wpscbe2=1.73315082665633e-14 ppscbe2=-3.60474574134596e-21
+  pvag=0.0
+  delta=0.01
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=18.2284323446247 lbeta0=-1.9625874645494e-06 wbeta0=-2.88303291590499e-07 pbeta0=5.9963625011327e-14
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-2.614334899479e-08 lagidl=5.45830167072838e-15 wagidl=2.10666837881197e-14 pagidl=-4.38161742772344e-21
+  bgidl=1020475725.30666 lbgidl=-3.64443339588342
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.426233527438381 lkt1=-3.74820317431458e-08 wkt1=-1.49167110928165e-07 pkt1=3.10249690677273e-14
+  kt2=-0.12
+  at=284803.119333333 lat=-0.0469343889119013 pat=5.29395592033938e-23
+  ute=-0.238289841333334 lute=4.60274143923742e-9
+  ua1=4.04904181333334e-10 lua1=-5.29130168671572e-17
+  ub1=8.54839297333336e-19 lub1=-8.64895837737656e-26
+  uc1=-4.07057654733333e-11 luc1=8.66210025306766e-18
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.04e-6
+  sbref=1.04e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.81 pmos
* DC IV MOS Parameters
+  lmin=2.0e-05 lmax=1.0e-04 wmin=6.4e-07 wmax=8.4e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.950462476053101+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} wvth0=-5.72017627060836e-8
+  k1=0.53274593583127 wk1=-3.38212013149867e-8
+  k2=-0.0043856305323825 wk2=1.39935634363696e-9
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=151381.852093917 wvsat=-0.0793565366430454
+  ua=-2.96695920428551e-09 wua=1.28375320954145e-15
+  ub=2.46710918726135e-18 wub=-9.05469429631458e-25
+  uc=5.20559427867161e-11 wuc=-7.50880239287529e-17
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=-0.000746420104814099 wu0=5.75978924428018e-9
+  a0=1.0919001832572 wa0=9.94571326643377e-8
+  keta=0.0042407059278715 wketa=1.98055447821016e-9
+  a1=0.0
+  a2=0.8
+  ags=0.45446425121193 wags=-1.37274345382494e-7
+  b0=3.5784941684e-07 wb0=-2.95366117434285e-13
+  b1=-8.7307878081e-07 wb1=7.20632415666084e-13
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.14070598491445+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} wvoff=-9.22375165161974e-8
+  nfactor={1.2571207257031+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} wnfactor=2.49096824146482e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.0017402344
+  pdiblc1=0.39
+  pdiblc2=-0.00027655585819909 wpdiblc2=6.96956384918783e-10
+  pdiblcb=-0.225
+  drout=0.56
+  pscbe1=830904617.828781 wpscbe1=-25.5205720191179
+  pscbe2=1.46936572682486e-08 wpscbe2=-3.2369292566595e-15
+  pvag=0.0
+  delta=0.01
+  alpha0=-3.126961e-10 walpha0=2.5809692191042e-16
+  alpha1=-3.126961e-10 walpha1=2.5809692191042e-16
+  beta0=114.427947 wbeta0=-6.96861689158134e-5
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-9.33726204948599e-11 wagidl=1.75209766490886e-16
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.60814922 wkt1=5.16193843820841e-8
+  kt2=-0.052484
+  at=10000.0
+  ute=-1.2595
+  ua1=-2.5605e-10
+  ub1=4.9434e-19
+  uc1=8.1951e-12
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.82 pmos
* DC IV MOS Parameters
+  lmin=8e-06 lmax=2.0e-05 wmin=6.4e-07 wmax=8.4e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.9504624760531+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} wvth0=-5.72017627060844e-8
+  k1=0.53274593583127 wk1=-3.38212013149867e-8
+  k2=-0.0043856305323825 wk2=1.39935634363696e-9
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=151381.852093917 wvsat=-0.0793565366430454
+  ua=-2.96695920428551e-09 wua=1.28375320954145e-15
+  ub=2.46710918726135e-18 wub=-9.05469429631458e-25
+  uc=5.2055942786716e-11 wuc=-7.50880239287529e-17
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=-0.000746420104814099 wu0=5.75978924428018e-9
+  a0=1.0919001832572 wa0=9.94571326643368e-8
+  keta=0.0042407059278715 wketa=1.98055447821017e-9
+  a1=0.0
+  a2=0.8
+  ags=0.45446425121193 wags=-1.37274345382494e-7
+  b0=3.5784941684e-07 wb0=-2.95366117434285e-13
+  b1=-8.7307878081e-07 wb1=7.20632415666084e-13
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.14070598491445+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} wvoff=-9.22375165161972e-8
+  nfactor={1.2571207257031+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} wnfactor=2.49096824146482e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.0017402344
+  pdiblc1=0.39
+  pdiblc2=-0.000276555858199089 wpdiblc2=6.96956384918783e-10
+  pdiblcb=-0.225
+  drout=0.56
+  pscbe1=830904617.82878 wpscbe1=-25.5205720191175
+  pscbe2=1.46936572682486e-08 wpscbe2=-3.2369292566595e-15
+  pvag=0.0
+  delta=0.01
+  alpha0=-3.126961e-10 walpha0=2.5809692191042e-16
+  alpha1=-3.126961e-10 walpha1=2.5809692191042e-16
+  beta0=114.427947 wbeta0=-6.96861689158134e-5
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-9.337262049486e-11 wagidl=1.75209766490886e-16
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.60814922 wkt1=5.16193843820844e-8
+  kt2=-0.052484
+  at=10000.0
+  ute=-1.2595
+  ua1=-2.5605e-10
+  ub1=4.9434e-19
+  uc1=8.1951e-12
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.83 pmos
* DC IV MOS Parameters
+  lmin=4e-06 lmax=8e-06 wmin=6.4e-07 wmax=8.4e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.80032033666693+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0=-1.2053392932865e-06 wvth0=-1.78414982827196e-07 pvth0=9.73098276573647e-13
+  k1=0.656080299923008 lk1=-9.90126794916101e-07 wk1=-1.00701839606663e-07 pk1=5.36916961637919e-13
+  k2=-0.00169830334201462 lk2=-2.15738304363471e-08 wk2=-1.08640896303699e-08 pk2=9.84507971179755e-14
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=302434.794026307 lvsat=-1.21265120519792 wvsat=-0.193651473610683 pvsat=9.1755838243695e-7
+  ua=-5.15378635516125e-09 lua=1.75558221253047e-14 wua=2.60930081836358e-15 pua=-1.06414802970528e-20
+  ub=2.75485325774249e-18 lub=-2.31000594489376e-24 wub=-8.22259720544395e-25 pub=-6.68006546034432e-31
+  uc=1.0239789727854e-10 luc=-4.04144606556908e-16 wuc=-1.03628764156649e-16 puc=2.2912472006067e-22
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=-0.0149702268071506 lu0=1.14188549520677e-07 wu0=1.56615699709415e-08 pu0=-7.9491376852268e-14
+  a0=1.40286571325168 la0=-2.49642754320936e-06 wa0=-9.31474952366449e-08 pa0=1.54622764153354e-12
+  keta=0.0286207430774165 lketa=-1.95722645676101e-07 wketa=-1.53017364418867e-08 pketa=1.38742024119046e-13
+  a1=0.0
+  a2=0.8
+  ags=0.228150153725404 lags=1.81684685885266e-06 wags=4.84140358384657e-09 pags=-1.14090352731279e-12
+  b0=7.91876123627729e-07 lb0=-3.48436119377141e-12 wb0=-6.53608375808563e-13 pb0=2.87596455132161e-18
+  b1=-1.71341295281859e-06 lb1=6.74619264887489e-12 wb1=1.41423768663543e-12 pb1=-5.56825479207868e-18
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={0.00226276346076126+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff=-1.14775139633121e-06 wvoff=-2.19597022629415e-07 pvoff=1.02244058676284e-12
+  nfactor={0.431089270255342+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor=6.63137061195712e-06 wnfactor=5.93174118596954e-07 pnfactor=-2.76224839092085e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=1.10455555171378 lpclm=-8.85338813361125e-06 wpclm=-9.40396119022292e-07 ppclm=7.54948875875753e-12
+  pdiblc1=0.39
+  pdiblc2=-0.00351433207547088 lpdiblc2=2.59928286189433e-08 wpdiblc2=2.9787030466736e-09 ppdiblc2=-1.83178348196078e-14
+  pdiblcb=-0.225
+  drout=0.56
+  pscbe1=862025558.385254 lpscbe1=-249.838537336094 wpscbe1=-51.2197634612185 ppscbe1=0.00020631280050689
+  pscbe2=2.01615025709145e-08 lpscbe2=-4.38957964756584e-14 wpscbe2=-6.69521913183589e-15 ppscbe2=2.77631096184376e-20
+  pvag=0.0
+  delta=0.01
+  alpha0=-5.60565689369467e-10 lalpha0=1.98989408902301e-15 walpha0=4.62686547593181e-16 palpha0=-1.6424430599057e-21
+  alpha1=-6.27580028736629e-10 lalpha1=2.52788440129051e-15 walpha1=5.17999660594989e-16 palpha1=-2.08649606732686e-21
+  beta0=179.501412415642 lbeta0=-0.000522408999475192 wbeta0=-0.000123397299696854 pbeta0=4.31192313376628e-10
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=4.08150439564903e-09 lagidl=-3.35158625870789e-14 wagidl=-3.32994149788637e-15 pagidl=2.81393122886054e-20
+  bgidl=2012767503.31827 lbgidl=-8130.48536342901 wbgidl=-835.930397652373 pbgidl=0.00671083920118848
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.540885823082166 lkt1=-5.39989743295614e-07 wkt1=-7.39916514590096e-08 pkt1=1.00840388839987e-12
+  kt2=-0.178494104302999 lkt2=1.01160760522323e-06 wkt2=8.26118442201334e-08 pkt2=-6.632068940571e-13
+  at=-11866.5628524492 lat=0.175544504180708 wat=-0.0195772141613182 pat=1.57165640360492e-7
+  ute=-3.38260966720648 lute=1.70442989310176e-05 wute=7.63724454415591e-07 pute=-6.13117075535491e-12
+  ua1=-7.31153498536269e-09 lua1=5.66413487966719e-14 wua1=4.01521276971959e-15 pua1=-3.22340799327556e-20
+  ub1=6.54537531720348e-18 lub1=-4.85776389140857e-23 wub1=-3.73954746101202e-24 pub1=3.00210421424349e-29
+  uc1=2.09108936411466e-10 luc1=-1.61293386774521e-15 wuc1=-9.25278153811954e-17 puc1=7.42812191546452e-22
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.84 pmos
* DC IV MOS Parameters
+  lmin=2e-06 lmax=4e-06 wmin=6.4e-07 wmax=8.4e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.25753459422649+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0=6.36314249592316e-07 wvth0=1.91040133401579e-07 pvth0=-5.15062498134467e-13
+  k1=0.321160683423464 lk1=3.5892540130866e-07 wk1=9.65375738956997e-08 pk1=-2.57561029076637e-13
+  k2=-0.0115142773622294 lk2=1.796479512539e-08 wk2=2.01809526111569e-08 pk2=-2.65982604903875e-14
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=-118454.570645007 lvsat=0.482686105025755 wvsat=0.124105138020798 pvsat=-3.62361436135315e-7
+  ua=7.02274779863739e-10 lua=-6.0323218538424e-15 wua=-1.10595332147339e-15 pua=4.32351879516086e-21
+  ub=2.49796314127376e-18 lub=-1.27525563843909e-24 wub=-1.38202560088203e-24 pub=1.58672370277502e-30
+  uc=-1.79935970959967e-11 luc=8.07908880857929e-17 wuc=-3.81733785542511e-17 puc=-3.45287876811628e-23
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0259886752641049 lu0=-5.0793416515515e-08 wu0=-1.39737962670433e-08 pu0=3.98795227299395e-14
+  a0=0.824588632002593 la0=-1.67134399262993e-07 wa0=3.19412504428851e-07 pa0=-1.15559086399074e-13
+  keta=-0.0368938819187056 lketa=6.81694776327784e-08 wketa=3.98378477382317e-08 pketa=-8.33595592834604e-14
+  a1=0.0
+  a2=0.8
+  ags=1.32952570042773 lags=-2.61948062675775e-06 wags=-8.98623888902996e-07 pags=2.4982438292407e-12
+  b0=-3.95062481831673e-07 lb0=1.2966132657558e-12 wb0=3.26081491016504e-13 pb0=-1.07021447597136e-18
+  b1=1.3294477068416e-09 lb1=-1.60769163532736e-13 wb1=-1.09731576753494e-15 pb1=1.32697613580445e-19
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.371907071953499+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff=3.594002106794e-07 wvoff=1.10615719330791e-07 pvoff=-3.07652375299967e-13
+  nfactor={3.57053313598733+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor=-6.01427160588491e-06 wnfactor=-1.0716268704713e-06 pnfactor=3.9435500154342e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.160612523 leta0=-3.24706275293724e-7
+  etab=-0.140472576764777 letab=2.83862693537599e-07 wetab=-3.89946006240709e-15 petab=1.57069784342903e-20
+  dsub=0.864198200000001 ldsub=-1.2253066992216e-6
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-2.72301199405387 lpclm=6.56400800993033e-06 wpclm=2.01588322260007e-06 ppclm=-4.35836895394526e-12
+  pdiblc1=0.39
+  pdiblc2=0.00593487442439421 lpdiblc2=-1.20684617720353e-08 wpdiblc2=-3.35322708801526e-09 ppdiblc2=7.18710377975736e-15
+  pdiblcb=0.4091439384468 lpdiblcb=-2.55432417433645e-06 wpdiblcb=-5.23417460471269e-07 ppdiblcb=2.10831924976875e-12
+  drout=0.56
+  pscbe1=799999833.766506 lpscbe1=0.000337119528921903 wpscbe1=0.000103961129752861 ppscbe1=-2.10831924835064e-10
+  pscbe2=9.64880370804336e-09 lpscbe2=-1.55077160839974e-15 wpscbe2=-1.10167915833004e-17 ppscbe2=8.39222802328199e-22
+  pvag=0.0
+  delta=0.01
+  alpha0=-1.35008944937042e-10 lalpha0=2.75756629130135e-16 walpha0=1.08883502551995e-16 palpha0=-2.17328640116342e-22
+  alpha1=1.04123206521175e-14 lalpha1=-4.23642029235366e-20 walpha1=-6.14714443645029e-21 palpha1=2.51101778559406e-26
+  beta0=97.2682858590333 lbeta0=-0.000191174952502689 wbeta0=-3.29252645173528e-05 pbeta0=6.67720413380173e-11
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-8.33822410973684e-09 lagidl=1.65106547958733e-14 wagidl=7.12616023595406e-15 pagidl=-1.3977740022083e-20
+  bgidl=-1025535006.63654 lbgidl=4107.76068703882 wbgidl=1671.86079530475 pbgidl=-0.00339051363054848
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.944475077367157 lkt1=1.08566292989328e-06 wkt1=4.06935423072798e-07 pkt1=-9.28764596689352e-13
+  kt2=0.15452570783273 lkt2=-3.29792201821745e-07 wkt2=-1.33893308929814e-07 pkt2=2.08873264769051e-13
+  at=159274.741919703 lat=-0.513810617745863 wat=-0.0458325454494327 pat=2.62921799725042e-7
+  ute=2.39403337397805 lute=-6.22394991915717e-06 wute=-1.34327432106563e-06 pute=2.35579502829815e-12
+  ua1=1.42087134312964e-08 lua1=-3.00419535826498e-14 wua1=-8.4084313991535e-15 pua1=1.78082096957352e-20
+  ub1=-1.25943146465141e-17 lub1=2.85168025834891e-23 wub1=8.08221117021491e-24 pub1=-1.75968597630436e-29
+  uc1=-4.9793710461712e-10 luc1=1.23503910096544e-15 wuc1=2.26228307709061e-16 puc1=-5.41133647187624e-22
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.85 pmos
* DC IV MOS Parameters
+  lmin=1e-06 lmax=2e-06 wmin=6.4e-07 wmax=8.4e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.884632724190526+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0=-1.19926268018177e-07 wvth0=-1.19574696795648e-07 pvth0=1.14860650127547e-13
+  k1=0.644716835770763 lk1=-2.97242592977832e-07 wk1=-1.44973332224921e-07 pk1=2.32220190405108e-13
+  k2=-0.0340285625151805 lk2=6.36234952441529e-08 wk2=3.16130702239516e-08 pk2=-4.9782457823724e-14
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=398654.417530706 lvsat=-0.566004717686734 wvsat=-0.264043626745382 pvsat=4.2479960102532e-7
+  ua=-6.73437798725114e-09 lua=9.04912071803336e-15 wua=4.48633223199662e-15 pua=-7.01756919984968e-21
+  ub=4.57710644369682e-18 lub=-5.49173330603344e-24 wub=-2.68554412322893e-24 pub=4.23024362387225e-30
+  uc=1.70316151541443e-10 luc=-3.01099022433951e-16 wuc=-1.74652179970549e-16 puc=2.42248583845472e-22
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=-0.0172205642434901 lu0=3.68344026950135e-08 wu0=1.99936786239411e-08 pu0=-2.90061087392781e-14
+  a0=3.08837480440868 la0=-4.75806559146846e-06 wa0=-1.24318143773657e-06 pa0=3.05336267718509e-12
+  keta=0.155795943219055 lketa=-3.22603175468699e-07 wketa=-1.04543606374224e-07 pketa=2.0944429707915e-13
+  a1=0.0
+  a2=-0.485791353787201 la2=2.6075694359842e-06 wa2=1.0612821542434e-06 pa2=-2.15226747341976e-12
+  ags=-3.71204363597739 lags=7.60476148863979e-06 wags=2.75492085238311e-06 pags=-4.91110106355062e-12
+  b0=3.6813473484763e-07 lb0=-2.51141531303228e-13 wb0=-3.03855538692302e-13 pb0=2.0729026103374e-19
+  b1=-1.35319374292177e-07 lb1=1.1635300769541e-13 wb1=1.11691556049644e-13 pb1=-9.60368649983313e-20
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.225170202535416+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff=6.18196003419603e-08 wvoff=-1.7730649631026e-08 pvoff=-4.73674792018301e-14
+  nfactor={-1.39723128963658+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor=4.06029503610725e-06 wnfactor=2.39179279905063e-06 pnfactor=-3.08022351332024e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=1.23671109163188 leta0=-2.50702125929636e-06 weta0=-1.08781420809948e-06 peta0=2.20607416025525e-12
+  etab=-0.501705675216391 letab=1.01643908240029e-06 wetab=4.19206458725062e-07 petab=-8.50145660018e-13
+  dsub=-1.0127399153404 ldsub=2.58110127543135e-06 wdsub=7.95961615682547e-07 pdsub=-1.61420060506482e-12
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=1.64596131932591 lpclm=-2.29621744192411e-06 wpclm=-1.08398527666548e-06 ppclm=1.9281271641433e-12
+  pdiblc1=0.424558783130533 lpdiblc1=-7.00847974833219e-08 wpdiblc1=-2.19396737182433e-08 ppdiblc1=4.44933950245121e-14
+  pdiblc2=0.000437487774803728 lpdiblc2=-9.19827615305554e-10 wpdiblc2=-1.83639673918353e-10 ppdiblc2=7.59218539017805e-16
+  pdiblcb=-2.3417811537872 lpdiblcb=3.024518901613e-06 wpdiblcb=1.57747599806424e-06 ppdiblcb=-2.15226747341976e-12
+  drout=0.12536052068447 ldrout=8.81443648378144e-07 wdrout=6.07123967490479e-08 pdrout=-1.23124012058308e-13
+  pscbe1=796130700.223832 lpscbe1=7.84689351447105 wpscbe1=3.19368985471101 ppscbe1=-6.47676470107508e-6
+  pscbe2=1.12929380733249e-08 lpscbe2=-4.88505637157819e-15 wpscbe2=-7.6893307944542e-16 ppscbe2=2.37626793911713e-21
+  pvag=0.0
+  delta=0.01
+  alpha0=-1.00838691094847e-10 lalpha0=2.0645976438121e-16 walpha0=3.4857964570735e-18 palpha0=-3.58335692831407e-24
+  alpha1=-1.02820048141589e-10 lalpha1=2.08496575648976e-16 walpha1=1.26438427045347e-20 palpha1=-1.2997718574203e-26
+  beta0=-6.20504158031115 lbeta0=1.86677138643721e-05 wbeta0=2.59078846359151e-06 pbeta0=-5.25408791470202e-12
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-3.06255224564405e-10 lagidl=2.21918280370195e-16 wagidl=3.14860782400601e-16 pagidl=-1.64506465870053e-22
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.316910684426488 lkt1=-1.8703012821768e-07 wkt1=-9.07787402715334e-08 pkt1=8.05937540029894e-14
+  kt2=0.0626045910175198 lkt2=-1.433772799739e-07 wkt2=-7.36858170437173e-08 pkt2=8.67731937139491e-14
+  at=-54145.3067505522 lat=-0.08099732008317 wat=0.037704490110603 pat=9.35096940537166e-8
+  ute=3.11446327404258 lute=-7.68497311132924e-06 wute=-3.05624628549178e-06 pute=5.82968161649081e-12
+  ua1=3.01809803043835e-09 lua1=-7.34751983709457e-15 wua1=-2.54370720042124e-15 pua1=5.9146193973965e-21
+  ub1=-6.24425004782261e-19 lub1=4.24201002873262e-24 wub1=1.35806036839567e-24 pub1=-3.96036262676375e-30
+  uc1=1.56350819388653e-11 luc1=1.9352086949614e-16 wuc1=5.04019084199468e-17 puc1=-1.84559819346092e-22
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=2.745e-6
+  sbref=2.74e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.86 pmos
* DC IV MOS Parameters
+  lmin=5e-07 lmax=1e-06 wmin=6.4e-07 wmax=8.4e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.17819267424358+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0=1.81849837916961e-07 wvth0=8.80809453862028e-08 pvth0=-9.86068581676895e-14
+  k1=0.284432272997548 lk1=7.31256141382783e-08 wk1=9.12615953036901e-08 pk1=-1.0626480275173e-14
+  k2=0.0381590533819347 lk2=-1.05845076466908e-08 wk2=-1.31110595933467e-08 pk2=-3.806589061099e-15
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=-267328.597220904 lvsat=0.118617829681745 wvsat=0.219157954556689 pvsat=-7.19258261342333e-8
+  ua=3.23754187697586e-09 lua=-1.20189323935362e-15 wua=-2.98275696308342e-15 pua=6.60564863622258e-22
+  ub=-1.36265473387054e-18 lub=6.14269907371677e-25 wub=1.70474884908505e-24 pub=-2.82924868150848e-31
+  uc=-2.0025731090297e-10 luc=7.98460500773559e-17 wuc=1.0168007265992e-16 puc=-4.18176558716188e-23
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0250705899864342 lu0=-6.64039635949789e-09 wu0=-1.19323628405558e-08 pu0=3.81347877372721e-15
+  a0=-4.4680483272819 la0=3.00984671083187e-06 wa0=3.63553538700901e-06 pa0=-1.96189967405146e-12
+  keta=-0.209895172663364 lketa=5.33229033650372e-08 wketa=1.38104140868282e-07 pketa=-3.99946753131797e-14
+  a1=0.0
+  a2=3.3715827075744 la2=-1.35776481060679e-06 wa2=-2.12256430848679e-06 pa2=1.12068848410932e-12
+  ags=4.60932970800124 lags=-9.49510452490119e-07 wags=-2.85223349516737e-06 pags=8.52986319879101e-13
+  b0=2.93276636540517e-08 lb0=9.7148072198916e-14 wb0=-2.42068248242778e-14 pb0=-8.01852610380221e-20
+  b1=-4.44131221110458e-08 lb1=2.2902471328233e-14 wb1=3.66582445681047e-14 pb1=-1.89035211950472e-20
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.116278783849872+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff=-5.01194713697536e-08 wvoff=-1.03567733845156e-07 pvoff=4.08720133252851e-14
+  nfactor={3.46968243908804+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor=-9.42833874056907e-07 wnfactor=-1.42992519229194e-06 pnfactor=8.48456721164027e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=-2.98882243526376 leta0=1.83677649995004e-06 weta0=2.17562841619896e-06 peta0=-1.14870569621206e-12
+  etab=1.00138993734189 letab=-5.28725170162269e-07 wetab=-8.38412901852283e-07 petab=4.42671951223183e-13
+  dsub=2.67956436099563 ldsub=-1.21454321299077e-06 wdsub=-1.53803920779866e-06 pdsub=7.85124233463982e-13
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-1.85485478310782 lpclm=1.30257950158453e-06 wpclm=1.61538769750725e-06 ppclm=-8.46795860830579e-13
+  pdiblc1=0.704329441393986 lpdiblc1=-3.57685676930253e-07 wpdiblc1=-6.79223259390925e-08 ppdiblc1=9.17630097157193e-14
+  pdiblc2=-0.00016724460365879 lpdiblc2=-2.98169987034628e-10 wpdiblc2=3.90387401869989e-11 ppdiblc2=5.30307801458473e-16
+  pdiblcb=0.6003922 wpdiblcb=-5.1619384382084e-7
+  drout=0.42109693342068 ldrout=5.77430164922273e-07 wdrout=3.27219270624388e-07 pdrout=-3.97089880319671e-13
+  pscbe1=807738599.552336 lpscbe1=-4.08588770043889 wpscbe1=-6.38737970942202 ppscbe1=3.37245983801811e-6
+  pscbe2=-2.38539883508921e-08 lpscbe2=3.12455622293997e-14 wpscbe2=2.58395368518847e-14 ppscbe2=-2.49769198486511e-20
+  pvag=0.0
+  delta=0.01
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=15.129968555878 lbeta0=-3.26442053550879e-06 wbeta0=-5.25537561589866e-06 pbeta0=2.81167460504493e-12
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-1.35460173060417e-10 lagidl=4.63430169647138e-17 wagidl=1.83059777141393e-16 pagidl=-2.90166140756497e-23
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.491803336822593 lkt1=-7.24258026631223e-09 wkt1=-2.28894882435408e-08 pkt1=1.08044175892376e-14
+  kt2=-0.167164157473485 lkt2=9.28222362498715e-08 wkt2=7.76818290073502e-08 pkt2=-6.88309300147958e-14
+  at=-338982.735166071 lat=0.211812138278842 wat=0.262086017470169 pat=-1.37151823493589e-7
+  ute=-8.22187538224392 lute=3.96864699126942e-06 wute=4.97076635086188e-06 pute=-2.42199104952912e-12
+  ua1=-9.88220749747184e-09 lua1=5.91383944193077e-15 wua1=7.2638459812738e-15 pua1=-4.16742758274782e-21
+  ub1=6.37173816541423e-18 lub1=-2.94996175627133e-24 wub1=-4.92545857067588e-24 pub1=2.49901944037454e-30
+  uc1=3.9350575589662e-10 luc1=-1.94925648884345e-16 wuc1=-2.65494524626574e-16 puc1=1.40177923068536e-22
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.745e-6
+  sbref=1.74e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.87 pmos
* DC IV MOS Parameters
+  lmin=2.5e-07 lmax=5e-07 wmin=6.4e-07 wmax=8.4e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.682127902238233+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0=-8.00664089245983e-08 wvth0=-2.08404703900477e-07 pvth0=5.79340068278854e-14
+  k1=0.248004431126993 lk1=9.23590775118292e-08 wk1=1.50234187624126e-07 pk1=-4.17633013492557e-14
+  k2=0.0622434603725366 lk2=-2.33007855248447e-08 wk2=-4.29162847746838e-08 pk2=1.19302121719448e-14
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=-286355.350088983 lvsat=0.128663726875056 wvsat=0.175147775904975 pvsat=-4.86889799282723e-8
+  ua=3.80594257632444e-09 lua=-1.50200198780128e-15 wua=-3.65718007920891e-15 pua=1.01665217585913e-21
+  ub=-2.13632510239344e-18 lub=1.02275857790735e-24 wub=2.46864826871947e-24 pub=-6.86254594924788e-31
+  uc=-1.0361126603803e-10 luc=2.8818098141206e-17 wuc=4.74728093277888e-17 puc=-1.31968713194133e-23
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0208743178024781 lu0=-4.42481500163527e-09 wu0=-9.94666247092871e-09 pu0=2.76505280696853e-15
+  a0=1.70005590370782 la0=-2.46838305879929e-07 wa0=-1.69522464541414e-07 pa0=4.71252108729386e-14
+  keta=-0.218911148872376 lketa=5.80832306116812e-08 wketa=1.31690615262332e-07 pketa=-3.66084107555452e-14
+  a1=0.0
+  a2=1.10720647359648 la2=-1.62201331581258e-7
+  ags=5.46761597336305 lags=-1.40267530116597e-06 wags=-2.61183495506931e-06 pags=7.26058775489808e-13
+  b0=4.50530906705166e-07 lb0=-1.25242185693156e-13 wb0=-3.71864696253371e-13 pb0=1.03373923182082e-19
+  b1=-2.1884967557354e-09 lb1=6.08375836133373e-16 wb1=1.80636815190931e-15 pb1=-5.02148669812964e-22
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.128711991236801+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff=-4.35548870679443e-08 wvoff=-5.5242029328605e-08 pvoff=1.53566212490002e-14
+  nfactor={1.47432825475324+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor=1.10689191021657e-07 wnfactor=3.73893514944764e-07 pnfactor=-1.03937910432465e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.49
+  etab=5.62973e-05 letab=-3.30242238324e-11 wetab=6.46234853557053e-27 petab=-1.54074395550979e-33
+  dsub=0.102632280904263 ldsub=1.46046002112506e-07 wdsub=-1.07768047132867e-07 pdsub=2.99582238863715e-14
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.584469873441449 lpclm=1.46453548223983e-08 wpclm=2.44378352035122e-08 ppclm=-6.79342493255385e-15
+  pdiblc1=-0.456899306415221 lpdiblc1=2.55429167168034e-07 wpdiblc1=2.23603346751158e-07 ppdiblc1=-6.21590471566608e-14
+  pdiblc2=-0.0138523478944929 lpdiblc2=6.92740032928629e-09 wpdiblc2=2.2036791512493e-09 ppdiblc2=-6.12596359897492e-16
+  pdiblcb=1.5181887075744 lpdiblcb=-4.84585542441192e-07 wpdiblcb=-1.09017662084511e-06 ppdiblcb=3.03056018475491e-13
+  drout=2.71905018696108 ldrout=-6.35861577508017e-07 wdrout=-8.97288128244968e-07 pdrout=2.49435332194562e-13
+  pscbe1=800079104.265281 lpscbe1=-0.0417661028166094
+  pscbe2=6.43630574234068e-08 lpscbe2=-1.53319793348808e-14 wpscbe2=-4.53358178611927e-14 ppscbe2=1.26028133355972e-20
+  pvag=0.0
+  delta=0.01
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=8.56253413650776 lbeta0=2.0310602870568e-07 wbeta0=1.47597377431285e-07 pbeta0=-4.10302997573688e-14
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-8.89721096196439e-10 lagidl=4.44583733249456e-16 wagidl=2.70547006150721e-16 pagidl=-7.52088211458265e-23
+  bgidl=691592551.5264 lbgidl=162.835431904679
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.498238101234401 lkt1=-3.84510187405127e-09 wkt1=-5.12383011797179e-09 pkt1=1.42436328683466e-15
+  kt2=0.0378077278790432 lkt2=-1.54004595536395e-08 wkt2=-1.11263425923452e-07 pkt2=3.09298972456086e-14
+  at=57326.2103039152 lat=0.00256577077803524 wat=0.00490579479380299 pat=-1.36375208313971e-9
+  ute=-1.28360684516316 lute=3.05324462913216e-07 wute=8.10055738118959e-07 pute=-2.25185774528213e-13
+  ua1=2.33700472094244e-09 lua1=-5.37757978845346e-16 wua1=-1.32881628314811e-15 pua1=3.69394980919776e-22
+  ub1=1.1688112088376e-18 lub1=-2.02878758322347e-25 wub1=-4.06254317757931e-25 pub1=1.12933825284892e-31
+  uc1=5.072625803232e-11 luc1=-1.39421873659686e-17
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.245e-6
+  sbref=1.24e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.88 pmos
* DC IV MOS Parameters
+  lmin=1.8e-07 lmax=2.5e-07 wmin=6.4e-07 wmax=8.4e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.92394398099186+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0=-1.28444408240355e-08 wvth0=1.98926680528029e-08 pvth0=-5.52992300666298e-15
+  k1=-2.40846499358988 lk1=8.30825699950024e-07 wk1=1.12191703028093e-06 pk1=-3.11879471413736e-13
+  k2=0.856328152214882 lk2=-2.44046800840715e-07 wk2=-2.25923500404571e-07 pk2=6.28040220304658e-14
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=543459.46810475 lvsat=-0.102014834804983 wvsat=-0.119823800433715 pvsat=3.33095786349676e-8
+  ua=-5.60434370133591e-11 lua=-4.28416219925532e-16 wua=6.37675808813097e-16 pua=-1.77266222740336e-22
+  ub=6.68390258815575e-19 lub=2.43081364075577e-25 wub=-8.44489771180884e-25 pub=2.34758022511031e-31
+  uc=-1.88949989961328e-12 luc=5.4066781591994e-19 wuc=1.17932328254525e-18 puc=-3.27837720668188e-25
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0098341395479334 lu0=-1.35577792901091e-09 wu0=8.81289673333922e-10 pu0=-2.44987953710752e-16
+  a0=1.98082893666874 la0=-3.24889839766669e-07 wa0=-1.63880615377184e-06 pa0=4.55568445074725e-13
+  keta=0.188768187392565 lketa=-5.52467327179371e-08 wketa=-2.55004180787399e-07 pketa=7.08881022087276e-14
+  a1=0.0
+  a2=-0.129692156859157 la2=1.81641644901844e-07 wa2=1.39418922025282e-07 pa2=-3.87567872959642e-14
+  ags=-2.03898102803885 lags=6.84068586059746e-7
+  b0=-7.05986321635221e-07 lb0=1.96255725578732e-13 wb0=5.82715603184402e-13 pb0=-1.61987945098026e-19
+  b1=6.71488819302796e-08 lb1=-1.86665833900346e-14 wb1=-5.54241633839737e-14 pb1=1.54072523307841e-20
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-1.30744990194489+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff=2.84120107253977e-07 wvoff=9.39935620720343e-07 pvoff=-2.61290823332807e-13
+  nfactor={-11.4875599540154+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor=3.71393857040084e-06 wnfactor=1.03047249046002e-05 pnfactor=-2.86458986678e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.503041913103093 leta0=-3.62549533970225e-09 weta0=6.72563438142064e-07 peta0=-1.86964565042236e-13
+  etab=-0.532087212115869 letab=1.47896485671666e-07 wetab=5.16362328217497e-07 petab=-1.43542530896525e-13
+  dsub=1.61531859349785 ldsub=-2.7446264055276e-07 wdsub=6.4311216670925e-08 pdsub=-1.78777464999171e-14
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.718485472944057 lpclm=-2.2609373652132e-08 wpclm=-3.01129288729016e-08 ppclm=8.37103287152006e-15
+  pdiblc1=1.53929200445416 lpdiblc1=-2.99488062957922e-07 wpdiblc1=-1.29685625130147e-07 ppdiblc1=3.60510475586792e-14
+  pdiblc2=0.046985619865208 lpdiblc2=-9.98482465229743e-09 wpdiblc2=-8.18137047368248e-09 ppdiblc2=2.27432281523804e-15
+  pdiblcb=0.0260830744133318 lpdiblcb=-6.97980816900133e-08 wpdiblcb=-5.7510988165907e-07 ppdiblcb=1.59873645782641e-13
+  drout=-1.256946487644 ldrout=4.694177860721e-7
+  pscbe1=799717484.766857 lpscbe1=0.0587597783105593
+  pscbe2=-6.92572842854773e-08 lpscbe2=2.18128722160884e-14 wpscbe2=6.43278432297555e-14 ppscbe2=-1.78823684837533e-20
+  pvag=0.0
+  delta=0.01
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=6.91463038118624 lbeta0=6.61203497839997e-07 wbeta0=3.1913897848047e-06 pbeta0=-8.87168063498287e-13
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=3.69441107258675e-09 lagidl=-8.29750000086244e-16 wagidl=-9.68723087470566e-16 pagidl=2.69293393639768e-22
+  bgidl=2065239807.49686 lbgidl=-219.022021488037 wbgidl=22.6488071808599 pbgidl=-6.29609661059304e-6
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-3.77565282594474 lkt1=9.07236862618726e-07 wkt1=2.92518846288884e-06 pkt1=-8.13167290421542e-13
+  kt2=0.286688501485714 lkt2=-8.45863280470107e-08 wkt2=-2.64697796016969e-23
+  at=423445.367602224 lat=-0.0992109615210069 wat=-0.276396122574846 pat=7.68348053223362e-8
+  ute=0.687421120764791 lute=-2.42597659279163e-07 wute=-6.44556187293041e-07 pute=1.79178885393218e-13
+  ua1=1.2910594585422e-09 lua1=-2.46997747241229e-16 wua1=-1.15260910113199e-16 pua1=3.20411498805481e-23
+  ub1=-1.77551105515664e-19 lub1=1.71393808720088e-25 wub1=5.08896473394005e-25 pub1=-1.41467112845853e-31
+  uc1=2.16687075276997e-10 luc1=-6.00773030301819e-17 wuc1=-1.79284396288619e-16 puc1=4.98389107554807e-23
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.1e-6
+  sbref=1.1e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.89 pmos
* DC IV MOS Parameters
+  lmin=1.5e-07 lmax=1.8e-07 wmin=6.4e-07 wmax=8.4e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.469244128796294+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0=-1.07416553682487e-07 wvth0=-2.69736909323571e-07 pvth0=5.47095535326941e-14
+  k1=2.87063228078955 lk1=-2.67163183953605e-07 wk1=-2.47656954663507e-06 pk1=4.36562554745868e-13
+  k2=-0.219073747550769 lk2=-2.03761105122567e-08 wk2=4.39883365054233e-07 pk2=-7.56758163025798e-14
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=593220.662634369 lvsat=-0.112364566132809 wvsat=-0.172381785409631 pvsat=4.42410088141384e-8
+  ua=-3.57520475541252e-11 lua=-4.32636585436376e-16 wua=-7.79513245998855e-16 pua=1.17492094391894e-22
+  ub=-1.65455691486622e-18 lub=7.26226500835309e-25 wub=1.80174528967182e-24 pub=-3.15627115325602e-31
+  uc=3.80520059730702e-12 luc=-6.43761551033518e-19 wuc=-2.58572005255014e-18 puc=4.55246112511631e-25
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.00357970291373789 lu0=-5.49301623378517e-11 wu0=1.51173517371691e-09 pu0=-3.76113052444409e-16
+  a0=-3.11032092071965 la0=7.34008236771827e-07 wa0=3.65902889393257e-06 pa0=-6.46317670827218e-13
+  keta=-2.90179189141525 lketa=5.87552676953143e-07 wketa=2.07710686917323e-06 pketa=-4.14163010850485e-13
+  a1=0.0
+  a2=-0.774392447299292 la2=3.15731568909907e-07 wa2=-3.2531081805899e-07 pa2=5.79014218846835e-14
+  ags=17.6814685941055 lags=-3.41754828995082e-06 wags=-1.02761122932986e-05 pags=2.13730804365858e-12
+  b0=4.18392337074251e-06 lb0=-8.20786811519528e-13 wb0=-3.45337771560858e-12 pb0=6.77471032091088e-19
+  b1=-1.44630239680196e-07 lb1=2.53809325554851e-14 wb1=1.19376671716165e-13 pb1=-2.09492237600235e-20
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={0.309599767841256+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff=-5.22068194655049e-08 wvoff=-1.00529470437396e-06 pvoff=1.43293741522907e-13
+  nfactor={28.070582695607+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor=-4.51368040300882e-06 wnfactor=-1.70420051536881e-05 pnfactor=2.82320182458327e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=-0.00637465344417176 leta0=1.0232703750333e-07 weta0=-7.51747679878731e-07 peta0=1.09275055772673e-13
+  etab=2.25739932157671 letab=-4.32283239497985e-07 wetab=-1.84052010277455e-06 petab=3.46660732160648e-13
+  dsub=0.596558858858248 ldsub=-6.25728408645384e-08 wdsub=-2.23502977643825e-07 pdsub=4.19841521472192e-14
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=1.37267020192843 lpclm=-1.58671947064135e-07 wpclm=1.02939337494951e-06 ppclm=-2.11993564247895e-13
+  pdiblc1=0.392298716780865 lpdiblc1=-6.09272230413295e-08 wpdiblc1=4.51898795515568e-07 ppdiblc1=-8.49115329225817e-14
+  pdiblc2=-0.0136191705894393 lpdiblc2=2.62024450478374e-09 wpdiblc2=2.23820988757436e-08 ppdiblc2=-4.08251204781038e-15
+  pdiblcb=-2.25935770971245 lpdiblcb=4.05546176118739e-07 wpdiblcb=1.43579660396326e-06 ppdiblcb=-2.58370772348975e-13
+  drout=1.0
+  pscbe1=1557294026.57566 lpscbe1=-157.508069999418 wpscbe1=-473.484409808392 ppscbe1=9.84790754272277e-5
+  pscbe2=1.9905375425348e-07 lpscbe2=-3.39926040675522e-14 wpscbe2=-1.53674442291722e-13 ppscbe2=2.74594908772879e-20
+  pvag=0.0
+  delta=0.01
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=35.2315556743004 lbeta0=-5.22837716002422e-06 wbeta0=-1.43225486635428e-05 pbeta0=2.75552096649661e-12
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=2.45100569382934e-08 lagidl=-5.15915455240284e-15 wagidl=-2.07422423724811e-14 pagidl=4.38194812269053e-21
+  bgidl=1084502519.78733 lbgidl=-15.040434491907 wbgidl=-52.8472167553409 pbgidl=9.4061704158494e-6
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=5.18207495156557 lkt1=-9.55863022370089e-07 wkt1=-4.7782211846919e-06 pkt1=7.8904947535948e-13
+  kt2=-0.12
+  at=-112598.585960197 lat=0.012279748292534 wat=0.32801226781598 pat=-4.88748869782707e-8
+  ute=-1.48770899348361 lute=2.09803302923133e-07 wute=1.03126082271545e-06 pute=-1.69370942884428e-13
+  ua1=1.32279813775936e-09 lua1=-2.53599011654247e-16 wua1=-7.5762251206118e-16 pua1=1.65644654746505e-22
+  ub1=2.29345854353655e-18 lub1=-3.42546546166984e-25 wub1=-1.18742510458602e-24 pub1=2.11347419515056e-31
+  uc1=-5.47531802848994e-10 luc1=9.88710529934868e-17 wuc1=4.18330258006779e-16 puc1=-7.44577659621106e-23
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.04e-6
+  sbref=1.04e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.90 pmos
* DC IV MOS Parameters
+  lmin=2.0e-05 lmax=1.0e-04 wmin=5.5e-07 wmax=6.4e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.0419279+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+  k1=0.47866595
+  k2=-0.0021480645
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=24491.02
+  ua=-9.1424219e-10
+  ub=1.01926665e-18
+  uc=-6.8009552e-11
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0084634633
+  a0=1.2509318
+  keta=0.0074076058
+  a1=0.0
+  a2=0.8
+  ags=0.23496304
+  b0=-1.1444e-7
+  b1=2.7921e-7
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.28819346+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.6554257+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.0017402344
+  pdiblc1=0.39
+  pdiblc2=0.00083787503
+  pdiblcb=-0.225
+  drout=0.56
+  pscbe1=790097310.0
+  pscbe2=9.5178184e-9
+  pvag=0.0
+  delta=0.01
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=3.0
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=1.867872e-10
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.52561
+  kt2=-0.052484
+  at=10000.0
+  ute=-1.2595
+  ua1=-2.5605e-10
+  ub1=4.9434e-19
+  uc1=8.1951e-12
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.91 pmos
* DC IV MOS Parameters
+  lmin=8e-06 lmax=2.0e-05 wmin=5.5e-07 wmax=6.4e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.0419279+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+  k1=0.47866595
+  k2=-0.0021480645
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=24491.02
+  ua=-9.1424219e-10
+  ub=1.01926665e-18
+  uc=-6.8009552e-11
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0084634633
+  a0=1.2509318
+  keta=0.0074076058
+  a1=0.0
+  a2=0.8
+  ags=0.23496304
+  b0=-1.1444e-7
+  b1=2.7921e-7
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.28819346+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.6554257+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.0017402344
+  pdiblc1=0.39
+  pdiblc2=0.00083787503
+  pdiblcb=-0.225
+  drout=0.56
+  pscbe1=790097310.0
+  pscbe2=9.5178184e-9
+  pvag=0.0
+  delta=0.01
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=3.0
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=1.867872e-10
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.52561
+  kt2=-0.052484
+  at=10000.0
+  ute=-1.2595
+  ua1=-2.5605e-10
+  ub1=4.9434e-19
+  uc1=8.1951e-12
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.92 pmos
* DC IV MOS Parameters
+  lmin=4e-06 lmax=8e-06 wmin=5.5e-07 wmax=6.4e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.0856052871783+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0=3.50641540138743e-7
+  k1=0.49505840101435 lk1=-1.31598400033788e-7
+  k2=-0.0190699456975955 lk2=1.35848659191723e-07 wk2=3.30872245021211e-24
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=-7213.25340806 lvsat=0.254521526468625
+  ua=-9.8152322433938e-10 lua=5.40131336304132e-16
+  ub=1.44006276220322e-18 lub=-3.37814613921411e-24
+  uc=-6.3304144027139e-11 luc=-3.77749587412317e-17
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0100725702903211 lu0=-1.29178916090139e-8
+  a0=1.2539231852882 la0=-2.40148051970651e-8
+  keta=0.00415331856862559 lketa=2.61253788420269e-8
+  a1=0.0
+  a2=0.8
+  ags=0.23589154158385 lags=-7.45399957312793e-9
+  b0=-2.53241445489e-07 lb0=1.11429633876835e-12 wb0=1.0097419586829e-28
+  b1=5.47948296387e-07 lb1=-2.15742781853528e-12
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.34887212857885+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff=4.87127623206986e-7
+  nfactor={1.3795726677089+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor=2.21454483299657e-6
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-0.399134643050864 lpclm=3.218218705677e-06 wpclm=-9.42985898310452e-23 ppclm=-2.39813715187188e-28
+  pdiblc1=0.39
+  pdiblc2=0.00124860396158491 lpdiblc2=-3.29732693401648e-9
+  pdiblcb=-0.225
+  drout=0.56
+  pscbe1=780125330.878071 lpscbe1=80.0549287271133
+  pscbe2=9.45586995855402e-09 lpscbe2=4.97321344547225e-16
+  pvag=0.0
+  delta=0.01
+  alpha0=1.79268526012786e-10 lalpha0=-6.36366775608334e-16
+  alpha1=2.00699666141224e-10 lalpha1=-8.08415711385755e-16
+  beta0=-17.810449959447 lbeta0=0.000167066042549041 wbeta0=6.7762635780344e-21 pbeta0=-2.58493941422821e-26
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-1.2430607298616e-09 lagidl=1.14788020227538e-14 pagidl=2.25694915357879e-36
+  bgidl=676117641.595701 lbgidl=2600.12368668142
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.659198222020001 lkt1=1.0724446433179e-6
+  kt2=-0.0463980464689979 lkt2=-4.88579619154418e-8
+  at=-43170.461687961 lat=0.426851828385411 wat=1.38777878078145e-17 pat=-5.29395592033938e-23
+  ute=-2.16141686305 lute=7.24057775356305e-6
+  ua1=-8.9122342772e-10 lua1=5.09916465565503e-15 wua1=-3.94430452610506e-31
+  ub1=5.65851650275721e-19 lub1=-5.74094670273675e-25
+  uc1=6.1157274428481e-11 luc1=-4.25179700765752e-16 wuc1=1.23259516440783e-32 puc1=-9.4039548065783e-38
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.93 pmos
* DC IV MOS Parameters
+  lmin=2e-06 lmax=4e-06 wmin=5.5e-07 wmax=6.4e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.9520620709018+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0=-1.87268932504399e-7
+  k1=0.47552393562856 lk1=-5.2913807873411e-8
+  k2=0.020754997200448 lk2=-2.45657329022821e-8
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=79989.122801758 lvsat=-0.0967285984760076
+  ua=-1.0661408183375e-09 lua=8.80969989517428e-16 wua=7.88860905221012e-31
+  ub=2.88108907591218e-19 lub=1.26191016371678e-24
+  uc=-7.90326995252419e-11 luc=2.55794740624601e-17
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.003644622576778 lu0=1.29738046457651e-8
+  a0=1.3353281398328 la0=-3.51912985243237e-7
+  keta=0.0268067010726264 lketa=-6.51221740434983e-8
+  a1=0.0
+  a2=0.8
+  ags=-0.1073708404997 lags=1.37520275631082e-6
+  b0=1.26340712862e-07 lb0=-4.14656040083582e-13 wb0=-5.04870979341448e-29
+  b1=-4.25156471999993e-10 lb1=5.14138690993382e-14
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.1950329130964+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff=-1.32534890685738e-7
+  nfactor={1.857005416148+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor=2.9145145147685e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.160612523 leta0=-3.24706275293724e-7
+  etab=-0.140472583 letab=2.83862718653004e-7
+  dsub=0.864198200000001 ldsub=-1.2253066992216e-6
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.50037842015352 lpclm=-4.05009118753497e-7
+  pdiblc1=0.39
+  pdiblc2=0.0005730757194931 lpdiblc2=-5.76307281209572e-10
+  pdiblcb=-0.4277988 lpdiblcb=8.16871132814399e-7
+  drout=0.56
+  pscbe1=800000000.0
+  pscbe2=9.63118789578462e-09 lpscbe2=-2.0885720280246e-16
+  pvag=0.0
+  delta=0.01
+  alpha0=3.90954051843623e-11 lalpha0=-7.17511269888927e-17
+  alpha1=5.83057612939408e-16 lalpha1=-2.21311396537472e-21 walpha1=1.41059322098675e-37 palpha1=8.96831017167883e-44
+  beta0=44.620899918894 lbeta0=-8.44066855847181e-5
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=3.05648186189834e-09 lagidl=-5.83970394234418e-15
+  bgidl=1647764716.8086 lbgidl=-1313.65907251125
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.293786720408439 lkt1=-3.99428500235448e-7
+  kt2=-0.059569237594818 lkt2=4.19543788506765e-9
+  at=85988.65768419 lat=-0.093399554536181 wat=5.55111512312578e-17
+  ute=0.24614230487672 lute=-2.45704168413577e-06 pute=8.07793566946316e-28
+  ua1=7.63660232434117e-10 lua1=-1.56668686884183e-15
+  ub1=3.2911351618912e-19 lub1=3.79483692969539e-25
+  uc1=-1.36198810297074e-10 luc1=3.69768240235766e-16 wuc1=-4.93038065763132e-32
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.94 pmos
* DC IV MOS Parameters
+  lmin=1e-06 lmax=2e-06 wmin=5.5e-07 wmax=6.4e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.0758322575324+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0=6.37355207402162e-8
+  k1=0.4129049707924 lk1=7.40767013867425e-8
+  k2=0.016520629214348 lk2=-1.59784854388872e-8
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=-23550.443267656 lvsat=0.113248399037971
+  ua=4.39251987661599e-10 lua=-2.17194855633507e-15
+  ub=2.82930527801281e-19 lub=1.27241185579021e-24
+  uc=-1.089520900045e-10 luc=8.62556389217099e-17
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0147492598508 lu0=-9.54626649030418e-9
+  a0=1.1005319152 la0=1.24250940757385e-7
+  keta=-0.0113689276799161 lketa=1.22975429591129e-8
+  a1=0.0
+  a2=1.2111952 la2=-8.33898931257601e-7
+  ags=0.693065433792119 lags=-2.48072402717693e-7
+  b0=-1.177292377e-07 lb0=8.03148908167476e-14
+  b1=4.3275043818e-08 lb1=-3.72096126863782e-14
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.25352145096964+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff=-1.39208377412623e-8
+  nfactor={2.4272372583412+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor=-8.64971881708853e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=-0.502700126000001 leta0=1.02048381712649e-06 weta0=4.30133918527574e-23 peta0=-3.06078031225753e-28
+  etab=0.168604026 letab=-3.42940935479688e-07 wetab=-4.30133918527574e-23 petab=-9.78187522474055e-29
+  dsub=0.26
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-0.0873274499703598 lpclm=7.86851333387291e-7
+  pdiblc1=0.389477319501401 lpdiblc1=1.05998977899449e-9
+  pdiblc2=0.0001438485610138 lpdiblc2=2.94160245460547e-10
+  pdiblcb=0.1805976 lpdiblcb=-4.169494656288e-07 wpdiblcb=-2.64697796016969e-23 ppdiblcb=-5.04870979341448e-29
+  drout=0.22243943652168 ldrout=6.84568772007271e-7
+  pscbe1=801237399.43548 lpscbe1=-2.50943120636111
+  pscbe2=1.00634166954672e-08 lpscbe2=-1.08541202181314e-15
+  pvag=0.0
+  delta=0.01
+  alpha0=-9.52649144198684e-11 lalpha0=2.00729988844652e-16 walpha0=-2.46519032881566e-32 palpha0=2.93873587705572e-38
+  alpha1=-1.02799830680123e-10 lalpha1=2.08475792341198e-16 walpha1=-4.34161785510107e-33 palpha1=3.93163543278263e-38
+  beta0=-2.0623796417844 lbeta0=1.0266445164983e-5
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=1.9720609522916e-10 lagidl=-4.11269988482738e-17
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.462065581260081 lkt1=-5.81609897746535e-8
+  kt2=-0.055218779730816 lkt2=-4.62723845763395e-9
+  at=6144.04465261986 lat=0.0685243625564864
+  ute=-1.77246413805463 lute=1.63666795885169e-6
+  ua1=-1.04928112846583e-09 lua1=2.10993645576693e-15 wua1=-1.35585468084861e-31 pua1=2.11588983148012e-37
+  ub1=1.54710890369256e-18 lub1=-2.09059633694279e-24 pub1=-7.00649232162409e-46
+  uc1=9.62275620176813e-11 luc1=-1.01589653702089e-16
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=2.745e-6
+  sbref=2.74e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.95 pmos
* DC IV MOS Parameters
+  lmin=5e-07 lmax=1e-06 wmin=5.5e-07 wmax=6.4e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.0373515422528+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0=2.41778072013713e-8
+  k1=0.430359253384721 lk1=5.61339083332286e-8
+  k2=0.0171945137005208 lk2=-1.6671230604059e-08 wk2=-4.96308367531817e-24 pk2=-5.52202633654708e-30
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=83104.2264642799 lvsat=0.00360867840957768
+  ua=-1.5318763586264e-09 lua=-1.45652269891164e-16
+  ub=1.3632328756728e-18 lub=1.6187400580647e-25
+  uc=-3.767122067044e-11 luc=1.29797606167283e-17
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.00599078240239999 lu0=-5.42656775078368e-10
+  a0=1.3451603872 la0=-1.27224192916953e-7
+  keta=0.0109328787070922 lketa=-1.0628446385055e-08 wketa=2.48154183765908e-24 pketa=3.15544362088405e-30
+  a1=0.0
+  a2=-0.0223903999999999 la2=4.342122625152e-7
+  ags=0.0486180535108804 lags=4.14411770842858e-7
+  b0=-9.37896688e-09 lb0=-3.10678873829625e-14
+  b1=1.420328622936e-08 lb1=-7.32419474634733e-15
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.28188323789512+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff=1.52347388766883e-8
+  nfactor={1.183236921712+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor=4.13845536341924e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.49
+  etab=-0.33922944015 letab=1.79105773720918e-7
+  dsub=0.22024490066552 ldsub=4.08677650546537e-8
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.728144649100079 lpclm=-5.14441987919331e-8
+  pdiblc1=0.59572187331256 lpdiblc1=-2.10956936604232e-7
+  pdiblc2=-0.000104821790923039 lpdiblc2=5.49790383207395e-10 ppdiblc2=1.97215226305253e-31
+  pdiblcb=-0.225
+  drout=0.944319433836238 ldrout=-5.75152026721289e-8
+  pscbe1=797525201.12904 lpscbe1=1.30666410627964
+  pscbe2=1.74633431602536e-08 lpscbe2=-8.69244762849598e-15
+  pvag=0.0
+  delta=0.01
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=6.7266408266568 lbeta0=1.23143759167113e-6
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=1.5725178775616e-10 lagidl=-5.44502177193565e-20
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.528403550646081 lkt1=1.00336466985229e-8
+  kt2=-0.0429511771911121 lkt2=-1.72381866572192e-8
+  at=80091.9150616879 lat=-0.00749316084959051
+  ute=-0.273636899477624 lute=9.58915435213917e-8
+  ua1=1.7326575124752e-09 lua1=-7.49863083856756e-16
+  ub1=-1.50405333098736e-18 lub1=1.04596182636135e-24 pub1=3.50324616081204e-46
+  uc1=-3.10190856773144e-11 luc1=2.92183731685939e-17 wuc1=-9.24446373305873e-33 puc1=5.87747175411144e-39
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.745e-6
+  sbref=1.74e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.96 pmos
* DC IV MOS Parameters
+  lmin=2.5e-07 lmax=5e-07 wmin=5.5e-07 wmax=6.4e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.0153663147104+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0=1.25698708817146e-8
+  k1=0.48822838598944 lk1=2.55797007475276e-8
+  k2=-0.00637953296617763 lk2=-4.22441685260222e-9
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=-6294.65233007981 lvsat=0.0508102136264543
+  ua=-2.0418759273424e-09 lua=1.23621382396059e-16
+  ub=1.811035080096e-18 lub=-7.45601845025277e-26
+  uc=-2.77024054417689e-11 luc=7.71634580177271e-18
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.00496963835344 lu0=-3.5049709560796e-12
+  a0=1.42899005968 la0=-1.71485254030323e-7
+  keta=-0.00833830312480799 lketa=-4.53493631993675e-10
+  a1=0.0
+  a2=1.10720647359648 la2=-1.62201331581258e-7
+  ags=1.29130076657072 lags=-2.41709789460181e-7
+  b0=-1.44079477392e-07 lb0=4.00523657612473e-14
+  b1=6.9987977328e-10 lb1=-1.94558178414561e-16
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.2170438081808+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff=-1.89997019393162e-8
+  nfactor={2.0721827130352+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor=-5.550717412723e-8
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.49
+  etab=5.62972999999999e-05 letab=-3.30242238324e-11 petab=4.62223186652937e-33
+  dsub=-0.0696884597971197 ldsub=1.93949100178602e-7
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.62354588878592 lpclm=3.78269146881947e-9
+  pdiblc1=-0.0993583157358398 lpdiblc1=1.56037062251055e-07 ppdiblc1=-5.04870979341448e-29
+  pdiblc2=-0.0103286724293219 lpdiblc2=5.94786083407434e-09 wpdiblc2=1.65436122510606e-24 ppdiblc2=-1.18329135783152e-30
+  pdiblcb=-0.225
+  drout=1.28428952278112 ldrout=-2.37015329993958e-7
+  pscbe1=800079104.265282 lpscbe1=-0.0417661028168368
+  pscbe2=-8.12876108854878e-09 lpscbe2=4.8198763096207e-15 wpscbe2=1.57772181044202e-30 ppscbe2=-3.76158192263132e-37
+  pvag=0.0
+  delta=0.01
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=8.7985418408432 lbeta0=1.37498718992877e-7
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-4.5711735385568e-10 lagidl=3.24325084123633e-16 pagidl=9.4039548065783e-38
+  bgidl=691592551.5264 lbgidl=162.835431904679
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.50643108816 lkt1=-1.56754982457856e-9
+  kt2=-0.140102111616 lkt2=3.40563409079086e-8
+  at=65170.5594880001 lat=0.00038513583704991
+  ute=0.011669524 lute=-5.4746824397712e-8
+  ua1=2.12232005280001e-10 lua1=5.29033388362234e-17
+  ub1=5.19211936959999e-19 lub1=-2.22979559316367e-26
+  uc1=5.072625803232e-11 luc1=-1.39421873659686e-17
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.245e-6
+  sbref=1.24e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.97 pmos
* DC IV MOS Parameters
+  lmin=1.8e-07 lmax=2.5e-07 wmin=5.5e-07 wmax=6.4e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.892135672457144+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0=-2.16867688969838e-8
+  k1=-0.614523479319423 lk1=3.3213148628101e-7
+  k2=0.495077243737657 lk2=-1.43623383294948e-07 wk2=1.05879118406788e-22 pk2=-2.52435489670724e-29
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=351861.618893142 lvsat=-0.0487529318983468
+  ua=9.63598011685718e-10 lua=-7.11864306966487e-16
+  ub=-6.81946012057137e-19 lub=6.18458643342941e-25
+  uc=-3.76598328805711e-15 luc=1.64564159885244e-20
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0112433187371428 lu0=-1.74751283346087e-9
+  a0=-0.639616527428572 la0=4.03562553906815e-7
+  keta=-0.218982630074297 lketa=5.81031015280409e-08 wketa=-2.64697796016969e-23 pketa=6.31088724176809e-30
+  a1=0.0
+  a2=0.0932382251080011 la2=1.19669673879558e-7
+  ags=-2.03898102803885 lags=6.84068586059746e-7
+  b0=2.25773945257143e-07 lb0=-6.27624474941426e-14
+  b1=-2.14741667485714e-08 lb1=5.96956066610188e-15
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={0.195503957601716+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff=-1.33683030253665e-7
+  nfactor={4.98966010821142+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor=-8.66530880257481e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=1.57846856239943 leta0=-3.02581198724292e-7
+  etab=0.293574393861143 letab=-8.16275328506714e-08 wetab=5.91434137975415e-23 petab=1.97215226305253e-31
+  dsub=1.71815201014571 ldsub=-3.03049096379867e-7
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.670335002130859 lpclm=-9.22412057171261e-9
+  pdiblc1=1.33192513110629 lpdiblc1=-2.41842560569694e-7
+  pdiblc2=0.0339036363136342 lpdiblc2=-6.34819020876257e-9
+  pdiblcb=-0.893515669637313 lpdiblcb=1.85839333971137e-7
+  drout=-1.256946487644 ldrout=4.69417786072101e-7
+  pscbe1=799717484.766857 lpscbe1=0.0587597783114688
+  pscbe2=3.36027181733885e-08 lpscbe2=-6.78097414744674e-15
+  pvag=0.0
+  delta=0.01
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=12.01765178888 lbeta0=-7.57375217241974e-7
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=2.14542615165142e-09 lagidl=-3.99150779885276e-16
+  bgidl=2101455173.12 lbgidl=-229.089458546882
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=0.901713573714288 lkt1=-3.93014868089686e-7
+  kt2=0.286688501485714 lkt2=-8.45863280470106e-08 pkt2=1.89326617253043e-29
+  at=-18511.0919999997 lat=0.023647630770896
+  ute=-0.343222029714286 lute=4.39087688362148e-8
+  ua1=1.10675765542857e-09 lua1=-1.95764057597278e-16
+  ub1=6.36172624000001e-19 lub1=-5.48116234005122e-26
+  uc1=-6.99880644011428e-11 luc1=1.96149456986649e-17 wuc1=2.31111593326468e-32 puc1=-3.30607786168768e-39
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.1e-6
+  sbref=1.1e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.98 pmos
* DC IV MOS Parameters
+  lmin=1.5e-07 lmax=1.8e-07 wmin=5.5e-07 wmax=6.4e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.01282225636613+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0=3.41459231707771e-09 wvth0=7.02126117492048e-08 pvth0=-1.46033806924937e-14
+  k1=-4.88851898234773 lk1=1.22107126296486e-06 wk1=2.37594313195114e-06 pk1=-4.94167660128254e-13
+  k2=1.50150398554703 lk2=-3.52948068470396e-07 wk2=-6.36152528718813e-07 pk2=1.32312092143168e-13
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=654850.776176014 lvsat=-0.111771040743297 wvsat=-0.210924777703691 pvsat=4.38698226650353e-8
+  ua=3.14196323311354e-09 lua=-1.16493813264082e-15 wua=-2.76683159634921e-15 pua=5.7546777006148e-22
+  ub=-1.28134486079427e-18 lub=7.4312641109408e-25 wub=1.56834138210924e-24 pub=-3.26196187382136e-31
+  uc=1.7810784520001e-13 luc=-2.13711578510518e-20 wuc=-3.17364536705885e-19 puc=6.60080152603835e-26
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0164927877086097 lu0=-2.83933938589832e-09 wu0=-6.56400733493454e-09 pu0=1.36523475757837e-15
+  a0=-11.8177787646799 la0=2.72848616130825e-06 wa0=9.10460511137415e-06 pa0=-1.89364860790449e-12
+  keta=-0.457162210384712 lketa=1.07641596077644e-07 wketa=5.48254534768247e-07 pketa=-1.14030364177378e-13
+  a1=0.0
+  a2=-8.33568581458309 la2=1.87278472704683e-06 wa2=4.40346307575203e-06 pa2=-9.15867478199513e-13
+  ags=23.3086543735184 lags=-4.58793540583935e-06 wags=-1.37953103876943e-05 pags=2.86925901691577e-12
+  b0=-5.21268025187409e-06 lb0=1.06837076405879e-12 wb0=2.42318489646759e-12 pb0=-5.03993380246502e-19
+  b1=1.12349204198144e-07 lb1=-2.18640946103636e-14 wb1=-4.13362680456873e-14 pb1=8.5974477182864e-21
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-2.98901113441656+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff=5.28657894705032e-07 wvoff=1.05763082473304e-06 pvoff=-2.19974519974576e-13
+  nfactor={54.7127670491404+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor=-1.12083404466874e-05 wnfactor=-3.370381943935e-05 pnfactor=7.00998999755152e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=-7.15720513546989 leta0=1.51433410234815e-06 weta0=3.72032592710239e-06 peta0=-7.73783148926172e-13
+  etab=-1.47286370581888 letab=2.85770394625578e-07 wetab=4.92357298507041e-07 petab=-1.02404409801882e-13
+  dsub=0.0699005973160887 ldsub=3.97674184717412e-08 wdsub=1.058649911902e-07 pdsub=-2.20186477876675e-14
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=16.953341025109 lpclm=-3.3958939772789e-06 wpclm=-8.71463662863521e-06 ppclm=1.81253984311658e-12
+  pdiblc1=7.04922961070779 lpdiblc1=-1.43097328467305e-06 wpdiblc1=-3.71129386148536e-06 ppdiblc1=7.71904587662617e-13
+  pdiblc2=0.142856403880401 lpdiblc2=-2.90090584294393e-08 wpdiblc2=-7.5476504888214e-08 ppdiblc2=1.56982072986899e-14
+  pdiblcb=-2.39333422744247 lpdiblcb=4.97783596171917e-07 wpdiblcb=1.51958447313478e-06 ppdiblcb=-3.16055335398356e-13
+  drout=1.0
+  pscbe1=801348527.984619 lpscbe1=-0.280477638466436 wpscbe1=-0.721991364451242 ppscbe1=1.50165539909448e-7
+  pscbe2=-3.3724744808313e-08 lpscbe2=7.22233022319138e-15 wpscbe2=-8.09658465076991e-15 ppscbe2=1.68399244834433e-21
+  pvag=0.0
+  delta=0.01
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=14.1084083939135 lbeta0=-1.19222750200969e-06 wbeta0=-1.11229711493766e-06 pbeta0=2.31344452341652e-13
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-1.60692094359455e-08 lagidl=3.38927484670784e-15 wagidl=4.63571429969026e-15 pagidl=-9.64172945763979e-22
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-1.82151287806877 lkt1=1.73383555163768e-07 wkt1=-3.98231984023647e-07 pkt1=8.28274738931105e-14
+  kt2=-0.12
+  at=1006593.23617672 lat=-0.189561768237925 wat=-0.371921568052239 pat=7.73552230960491e-8
+  ute=6.56922441422295 lute=-1.3937971421454e-06 wute=-4.00748248638365e-06 pute=8.33508267377963e-13
+  ua1=-7.16984270367696e-10 lua1=1.83552378065237e-16 wua1=5.18041495678697e-16 pua1=-1.07746414603221e-22
+  ub1=5.26415890634492e-19 lub1=-3.19835399412866e-26 wub1=-8.23304123937596e-26 pub1=1.71237378129534e-32
+  uc1=7.09478228921501e-10 luc1=-1.42504689716925e-16 wuc1=-3.67794011184241e-16 puc1=7.64967407981879e-23
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.04e-6
+  sbref=1.04e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.99 pmos
* DC IV MOS Parameters
+  lmin=2.0e-05 lmax=1.0e-04 wmin=4.2e-07 wmax=5.5e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.12634583620754+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} wvth0=4.51967045856135e-8
+  k1=0.5433973549272 wk1=-3.46566892930645e-8
+  k2=-0.0852793716207807 wk2=4.45078534082705e-8
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=-211476.0232462 wvsat=0.126334914411078
+  ua=-1.38898106038814e-09 wua=2.5417148824262e-16
+  ub=2.4656318328274e-18 wub=-7.74372637237363e-25
+  uc=-1.35202780985493e-11 wuc=-2.91731322305003e-17
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0121208655760572 wu0=-1.95814465086329e-9
+  a0=0.178394076144155 wa0=5.74228331558174e-7
+  keta=-0.0465029744780326 wketa=2.88633041783325e-8
+  a1=0.0
+  a2=0.177878893076924 wa2=3.33078788101981e-7
+  ags=0.543504299226646 wags=-1.65190583568124e-7
+  b0=-2.48443950910769e-07 wb0=7.17446700868087e-14
+  b1=1.14984639526395e-06 wb1=-4.66131935060433e-13
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.415461382931554+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} wvoff=6.8138253247755e-8
+  nfactor={3.05861128106077+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} wnfactor=-7.51254615252403e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.00672845800311313 wpclm=-2.67065600896267e-9
+  pdiblc1=0.39
+  pdiblc2=-0.00408148750021257 wpdiblc2=2.63378832764807e-9
+  pdiblcb=-0.225
+  drout=0.56
+  pscbe1=1242087877.74128 wpscbe1=-241.992224442251
+  pscbe2=8.32815351435955e-09 wpscbe2=6.36937300385794e-16
+  pvag=0.0
+  delta=0.01
+  alpha0=4.11840153846154e-10 walpha0=-1.66956786016031e-16
+  alpha1=4.11840153846154e-10 walpha1=-1.66956786016031e-16
+  beta0=-81.1968415384615 wbeta0=4.50783322243283e-5
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-2.26198494850246e-10 wagidl=2.21109319734402e-16
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-1.10903174383077 wkt1=3.12359450957392e-7
+  kt2=-0.0323186599922416 wkt2=-1.07963657505018e-8
+  at=-223997.4452425 wat=0.125280407002762
+  ute=-4.24929865901538 wute=1.6007148816073e-6
+  ua1=-2.98627144930512e-09 wua1=1.46173926823066e-15
+  ub1=1.27170642412126e-18 wub1=-4.16195920016415e-25
+  uc1=-1.81977917287344e-10 wuc1=1.01817150106109e-16
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.100 pmos
* DC IV MOS Parameters
+  lmin=8e-06 lmax=2.0e-05 wmin=4.2e-07 wmax=5.5e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.15044424502738+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0=4.8264264266288e-07 wvth0=5.80988047001683e-08 pvth0=-2.58403106269095e-13
+  k1=0.564852267623844 lk1=-4.29698734029446e-07 wk1=-4.6143482202529e-08 pk1=2.30057350549239e-13
+  k2=-0.107540793365244 lk2=4.45851487561056e-07 wk2=5.64264449711666e-08 pk2=-2.38705408798586e-13
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=-292319.756188324 lvsat=1.61913731324007 wvsat=0.169618018447174 pvsat=-8.66873488237688e-7
+  ua=-1.43985562967835e-09 lua=1.01891526324946e-15 wua=2.81409335818957e-16 pua=-5.45519284404705e-22
+  ub=2.55171561834692e-18 lub=-1.72408502337961e-24 wub=-8.2046122455099e-25 pub=9.2306167365426e-31
+  uc=-3.94116632973286e-12 luc=-1.91850335556514e-16 wuc=-3.43017139544528e-17 puc=1.0271517322434e-22
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0126258656919944 lu0=-1.01141362619876e-08 wu0=-2.22851777393513e-09 pu0=5.41502966440533e-15
+  a0=-0.504927130230127 la0=1.36855489214096e-05 wa0=9.40073175545553e-07 pa0=-7.32713614524112e-12
+  keta=-0.0770795812570842 lketa=6.12387913651565e-07 wketa=4.52337809503038e-08 pketa=-3.27867712343321e-13
+  a1=0.0
+  a2=-0.238319505333507 la2=8.33561652898333e-06 wa2=5.55908164263418e-07 pa2=-4.46282407180875e-12
+  ags=0.729584329189762 lags=-3.72680860714094e-06 wags=-2.64816380186143e-07 pags=1.99530425915613e-12
+  b0=5.09372579307787e-08 lb0=-5.99600325810402e-12 wb0=-8.85416939535271e-14 pb0=3.21021337556348e-18
+  b1=1.89873890827308e-06 lb1=-1.49988102638369e-11 wb1=-8.67083145163925e-13 pb1=8.03024602453821e-18
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.398443040851588+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff=-3.40843150957435e-07 wvoff=5.90267656412101e-08 pvoff=1.82484764446033e-13
+  nfactor={4.40818246636896+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor=-2.70291955044983e-05 wnfactor=-1.47380450121116e-06 pnfactor=1.44712204453835e-11
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-4.31037554146123e-07 lcit=2.08912694961988e-10 wcit=5.58469614439691e-12 pcit=-1.11850227363628e-16
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=1.28515221638871 lpclm=-2.56042556918617e-05 wpclm=-6.87128764543298e-07 ppclm=1.37083187842284e-11
+  pdiblc1=0.39
+  pdiblc2=-0.00808025555849981 lpdiblc2=8.00872786861604e-08 wpdiblc2=4.77469755566421e-09 ppdiblc2=-4.28781043277965e-14
+  pdiblcb=-0.225
+  drout=0.56
+  pscbe1=1539133660.72275 lpscbe1=-5949.22937700359 wpscbe1=-401.028219693426 ppscbe1=0.00318517100445858
+  pscbe2=7.46574891732366e-09 lpscbe2=1.72722289205794e-14 wpscbe2=1.09866199488295e-15 ppscbe2=-9.24741664069265e-21
+  pvag=0.0
+  delta=0.01
+  alpha0=6.20460904929076e-10 lalpha0=-4.17825389923976e-15 walpha0=-2.78650708903969e-16 palpha0=2.23700454727256e-21
+  alpha1=6.20460904929076e-10 lalpha1=-4.17825389923976e-15 walpha1=-2.78650708903969e-16 palpha1=2.23700454727256e-21
+  beta0=-133.715720785245 lbeta0=0.00105184748332804 wbeta0=7.31965305257983e-05 pbeta0=-5.63150938163463e-10
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-3.41550686918799e-10 lagidl=2.31027231852267e-15 wagidl=2.82867983620807e-16 pagidl=-1.23690177921296e-21
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-1.21334211937223 lkt1=2.08912694961988e-06 wkt1=3.68206412401361e-07 pkt1=-1.11850227363628e-12
+  kt2=-0.0323186599922415 wkt2=-1.07963657505018e-8
+  at=-223997.4452425 wat=0.125280407002762
+  ute=-4.24929865901538 wute=1.6007148816073e-6
+  ua1=-2.98627144930512e-09 wua1=1.46173926823066e-15
+  ub1=1.27170642412126e-18 wub1=-4.16195920016415e-25
+  uc1=-1.96164128360983e-10 luc1=2.84121265148304e-16 wuc1=1.09412336862489e-16 puc1=-1.52116309214534e-22
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.101 pmos
* DC IV MOS Parameters
+  lmin=4e-06 lmax=8e-06 wmin=4.2e-07 wmax=5.5e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.28339293515391+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0=1.54995313161439e-06 wvth0=1.05893963982487e-07 pvth0=-6.42102071445644e-13
+  k1=0.578837878854054 lk1=-5.41975053158237e-07 wk1=-4.48548789554506e-08 pk1=2.19712459144934e-13
+  k2=-0.132263169415061 lk2=6.44322425820473e-07 wk2=6.06027690711861e-08 pk2=-2.72232888557653e-13
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=-284068.204935431 lvsat=1.55289395880046 wvsat=0.148225981579132 pvsat=-6.9513847296549e-7
+  ua=-1.58292081804459e-09 lua=2.16744087867137e-15 wua=3.21983580768536e-16 pua=-8.7124883596899e-22
+  ub=4.07000450455871e-18 lub=-1.39128899824212e-23 wub=-1.40805029531154e-24 pub=5.64021968265111e-30
+  uc=-8.4600927856893e-12 luc=-1.55572448195213e-16 wuc=-2.93630772510725e-17 puc=6.30678570332432e-23
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0184496687232666 lu0=-5.68675571114051e-08 wu0=-4.48503315963127e-09 pu0=2.35303081025893e-14
+  a0=1.21212221414844 la0=-9.89026106693711e-08 wa0=2.2379913900653e-08 pa0=4.00943469249966e-14
+  keta=-0.0142004248313807 lketa=1.07594800415894e-07 wketa=9.82645105716485e-09 pketa=-4.36180928491603e-14
+  a1=0.0
+  a2=0.8
+  ags=0.269181293730407 lags=-3.06985633096655e-08 wags=-1.78230736392001e-08 pags=1.24449581169448e-14
+  b0=-1.60618771923214e-06 lb0=7.30737617306016e-12 wb0=7.24356881981142e-13 pb0=-3.31572663725713e-18
+  b1=1.28943405233568e-06 lb1=-1.01073181920297e-11 wb1=-3.96985690146027e-13 pb1=4.25630929682399e-18
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.711656369270886+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff=2.17362969103274e-06 wvoff=1.94231852749439e-07 pvoff=-9.02940052397784e-13
+  nfactor={0.0109069084194164+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor=8.27207990741392e-06 wnfactor=7.32772971930666e-07 pnfactor=-3.24315703006947e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=2.55920076923077e-05 wcit=-8.34783930080153e-12
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.08
+  etab=-0.07
+  dsub=0.56
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-3.55518543240045 lpclm=1.32539168685659e-05 wpclm=1.68972497542161e-06 ppclm=-5.37303451796503e-12
+  pdiblc1=0.39
+  pdiblc2=0.00358729987432153 lpdiblc2=-1.35797163178641e-08 wpdiblc2=-1.25211954985107e-09 ppdiblc2=5.50511107347484e-15
+  pdiblcb=-0.225
+  drout=0.56
+  pscbe1=757003976.593337 lpscbe1=329.698341631138 wpscbe1=12.3789927374828 ppscbe1=-0.000133657136050199
+  pscbe2=9.36212194753825e-09 lpscbe2=2.0481689904929e-15 wpscbe2=5.0191953863338e-17 ppscbe2=-8.30311733027708e-22
+  pvag=0.0
+  delta=0.01
+  alpha0=4.26459619482637e-10 lalpha0=-2.62081390769117e-15 walpha0=-1.32344183353229e-16 palpha0=1.06245751582952e-21
+  alpha1=5.14721659958582e-10 lalpha1=-3.32938050948757e-15 walpha1=-1.68124926118261e-16 palpha1=1.34970488937829e-21
+  beta0=-88.3989569000244 lbeta0=0.000688045046658652 wbeta0=3.7792536025631e-05 pbeta0=-2.78928095164053e-10
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-6.12462556978797e-09 lagidl=4.87367280812978e-14 wagidl=2.61355173909082e-15 pagidl=-1.99476029999212e-20
+  bgidl=-333877603.132822 lbgidl=10708.3533914191 wbgidl=540.743576064741 pbgidl=-0.00434108293972483
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-1.55751699082723 lkt1=4.85215868756214e-06 wkt1=4.80952861932993e-07 pkt1=-2.02362941751882e-12
+  kt2=0.00424056330456918 lkt2=-2.93497005916117e-07 wkt2=-2.71115166916116e-08 pkt2=1.30977835973418e-13
+  at=-509706.415220086 lat=2.29366818247242 wat=0.249779710540662 pat=-9.99478914810623e-7
+  ute=-9.06389947841203 lute=3.86515576029065e-05 wute=3.69553535290043e-06 pute=-1.68171936056956e-11
+  ua1=-7.63719412710378e-09 lua1=3.73375514462955e-14 wua1=3.61174009387862e-15 pua1=-1.72601808282919e-20
+  ub1=3.05734698815079e-18 lub1=-1.43351010203423e-23 wub1=-1.33392717023468e-24 pub1=7.36753546397722e-30
+  uc1=-9.2654929824246e-13 luc1=-1.28324367671643e-15 wuc1=3.32391949694627e-17 puc1=4.5940075982498e-22
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.102 pmos
* DC IV MOS Parameters
+  lmin=2e-06 lmax=4e-06 wmin=4.2e-07 wmax=5.5e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.700823006190248+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0=-7.96631551412099e-07 wvth0=-1.34511435581861e-07 pvth0=3.26247993134753e-13
+  k1=0.427985192937786 lk1=6.56577554802654e-08 wk1=2.54518720344479e-08 pk1=-6.34822901613645e-14
+  k2=0.0801979339213927 lk2=-2.11468348885523e-07 wk2=-3.18252846654874e-08 pk2=1.00066202757023e-13
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=225623.524728826 lvsat=-0.500138211986417 wvsat=-0.0779715228434174 pvsat=2.15982360478488e-7
+  ua=-1.78008953695845e-09 lua=2.9616341124318e-15 wua=3.82242575149653e-16 pua=-1.11397134222819e-21
+  ub=-9.59433986835266e-19 lub=6.34562790765184e-24 wub=6.67924734841365e-25 pub=-2.72178282710443e-30
+  uc=-5.74447059131038e-11 luc=4.17369856666548e-17 wuc=-1.15580433935887e-17 puc=-8.65060568429516e-24
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=-0.00893928652546171 lu0=5.34548259630098e-08 wu0=6.73732677884816e-09 pu0=-2.16732230612866e-14
+  a0=1.52326109204192 la0=-1.35216627715779e-06 wa0=-1.00617836735738e-07 pa0=5.35527810515373e-13
+  keta=0.0545380124998506 lketa=-1.69282800293058e-07 wketa=-1.48471278339067e-08 pketa=5.57667868411293e-14
+  a1=0.0
+  a2=0.8
+  ags=-0.694088580084904 lags=3.84934092917993e-06 wags=3.1412410137555e-07 pags=-1.32463427947637e-12
+  b0=7.56537846142931e-07 lb0=-2.20965405156384e-12 wb0=-3.37402629620971e-13 pb0=9.61027934362043e-19
+  b1=-2.56075921569258e-06 lb1=5.40121408926893e-12 wb1=1.37078288470104e-12 pb1=-2.86424130943708e-18
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.00572646503784502+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff=-6.69847492059097e-07 wvoff=-1.01353195700256e-07 pvoff=2.87672975737006e-13
+  nfactor={1.87556588426301+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor=7.61255928623639e-07 wnfactor=-9.93712985712451e-09 pnfactor=-2.51529652589471e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=2.55920076923077e-05 wcit=-8.34783930080154e-12
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.160612523 leta0=-3.24706275293724e-7
+  etab=-0.140472583 letab=2.83862718653004e-7
+  dsub=0.8641982 ldsub=-1.2253066992216e-6
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.0961805721275844 lpclm=-1.453741581281e-06 wpclm=2.16404375089872e-07 ppclm=5.61483180324017e-13
+  pdiblc1=0.39
+  pdiblc2=0.00325723443517498 lpdiblc2=-1.22502166897671e-08 wpdiblc2=-1.43707763993809e-09 ppdiblc2=6.25012004084831e-15
+  pdiblcb=-1.06020688991815 lpdiblcb=3.36420333010764e-06 wpdiblcb=3.38586358559078e-07 ppdiblcb=-1.36382178923966e-12
+  drout=0.56
+  pscbe1=878255437.650689 lpscbe1=-158.701088490347 wpscbe1=-41.8973509257657 ppscbe1=8.49673249092419e-5
+  pscbe2=9.97523101600994e-09 lpscbe2=-4.21426980002176e-16 wpscbe2=-1.84198003032306e-16 ppscbe2=1.13808200668466e-22
+  pvag=0.0
+  delta=0.01
+  alpha0=-4.67033621947176e-10 lalpha0=9.78166146869217e-16 walpha0=2.70977533319814e-16 palpha0=-5.62117519068896e-22
+  alpha1=-6.2804179753986e-10 lalpha1=1.27365698415466e-15 walpha1=3.36248991841319e-16 palpha1=-6.81907199675885e-22
+  beta0=248.320664665369 lbeta0=-0.000668257548371293 wbeta0=-0.000109059265187098 pbeta0=3.12589197899203e-10
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=1.25986671978585e-08 lagidl=-2.66804705072689e-14 wagidl=-5.10881159982743e-15 pagidl=1.11579838608815e-20
+  bgidl=3667755206.26564 lbgidl=-5410.17554524424 wbgidl=-1081.48715212948 pbgidl=0.00219324296667276
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.102613801415074 lkt1=-1.00817390055175e-06 wkt1=-1.0235248968028e-07 pkt1=3.25917539115222e-13
+  kt2=-0.0729134658922656 lkt2=1.7278497840383e-08 wkt2=7.14439574547267e-09 pkt2=-7.0045682522081e-15
+  at=188057.184210266 lat=-0.516915222869843 wat=-0.054646692967554 pat=2.2674698540363e-7
+  ute=2.52936313191256 lute=-8.04596507232968e-06 wute=-1.22241862167254e-06 pute=2.99226598843659e-12
+  ua1=3.2341880759269e-09 lua1=-6.45224561092569e-15 wua1=-1.32270133728886e-15 pua1=2.61569004315351e-21
+  ub1=-8.89528535135056e-19 lub1=1.56286622494682e-24 wub1=6.52451448870964e-25 pub1=-6.33573777236884e-31
+  uc1=-6.97576530921233e-10 luc1=1.5228540894612e-15 wuc1=3.00557252875954e-16 puc1=-6.17353169605671e-22
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.103 pmos
* DC IV MOS Parameters
+  lmin=1e-06 lmax=2e-06 wmin=4.2e-07 wmax=5.5e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.29322771319337+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0=4.04758085533743e-07 wvth0=1.16391831276327e-07 pvth0=-1.82580821214449e-13
+  k1=0.307608382905939 lk1=3.09780481703131e-07 wk1=5.63749718410262e-08 pk1=-1.26193965491908e-13
+  k2=-0.0135669873388701 lk2=-2.13142137487654e-08 wk2=1.61086752191839e-08 pk2=2.85670731842799e-15
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=-251934.189863779 lvsat=0.468343102514813 wvsat=0.122274876534341 pvsat=-1.90114934502814e-7
+  ua=2.56729247533979e-09 lua=-5.85480443992489e-15 wua=-1.1393362783871e-15 pua=1.9717723137981e-21
+  ub=1.9374185703351e-18 lub=4.70845683941016e-25 wub=-8.85799992965876e-25 pub=4.29152276191922e-31
+  uc=-1.11385513785976e-10 luc=1.51128296743145e-16 wuc=1.30283611189661e-18 puc=-3.47323149908651e-23
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0370647341049756 lu0=-3.98407758272694e-08 wu0=-1.19475308549864e-08 pu0=1.62194440018384e-14
+  a0=-0.460648598564658 la0=2.67117876847607e-06 wa0=8.3584386986159e-07 pa0=-1.36360529292353e-12
+  keta=-0.0865780177215923 lketa=1.16898815603666e-07 wketa=4.02663601774111e-08 pketa=-5.60027054839671e-14
+  a1=0.0
+  a2=2.493466944288 la2=-3.43433064141273e-06 wa2=-6.86518290172189e-07 pa2=1.39225085424972e-12
+  ags=2.56634612704128 lags=-2.76278153165549e-06 wags=-1.00293987157619e-06 pags=1.34635565290209e-12
+  b0=-5.20682153676703e-07 lb0=3.80532781430375e-13 wb0=2.15737848181182e-13 pb0=-1.60734316934989e-19
+  b1=-9.88778115966359e-07 lb1=2.21325528279735e-12 wb1=5.52553211733899e-13 pb1=-1.20488135141581e-18
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.505117774979488+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff=3.42912091806837e-07 wvoff=1.34702709423545e-07 pvoff=-1.91045567183201e-13
+  nfactor={3.16233025622179+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.84828677653629e-06 wnfactor=-3.93563057339881e-07 pnfactor=5.2645912483443e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=2.55920076923077e-05 wcit=-8.34783930080154e-12
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=-0.502700126 leta0=1.02048381712649e-06 weta0=2.85377311330795e-23 peta0=-9.86076131526265e-31
+  etab=-0.0958645212593997 letab=1.93398104739807e-07 wetab=1.41594397348014e-07 petab=-2.87151738689004e-13
+  dsub=0.26
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-2.10406536529312 lpclm=3.00833077685695e-06 wpclm=1.07974574930807e-06 ppclm=-1.189362766494e-12
+  pdiblc1=0.377007194731406 lpdiblc1=2.63492531710464e-08 wpdiblc1=6.67640753488177e-09 ppdiblc1=-1.35396743638498e-14
+  pdiblc2=-0.00608661918204546 lpdiblc2=6.69900631971255e-09 wpdiblc2=3.33574383198553e-09 ppdiblc2=-3.42910463035514e-15
+  pdiblcb=1.44541377983631 lpdiblcb=-1.71716532070636e-06 wpdiblcb=-6.77172717118156e-07 ppdiblcb=6.96125427124859e-13
+  drout=-0.248320924845185 ldrout=1.63926513573494e-06 wdrout=2.52041425545001e-07 pdrout=-5.11136986508156e-13
+  pscbe1=729431656.367858 lpscbe1=143.111754065861 wpscbe1=38.4442347536087 ppscbe1=-7.79644467495018e-5
+  pscbe2=1.06741197222242e-08 lpscbe2=-1.83876488954022e-15 wpscbe2=-3.26965637042088e-16 ppscbe2=4.03339249228711e-22
+  pvag=0.0
+  delta=0.01
+  alpha0=-7.17712340361928e-11 lalpha0=1.76578767334398e-16 walpha0=-1.25783332267129e-17 palpha0=1.29303756170621e-23
+  alpha1=-1.02803044754604e-10 lalpha1=2.08479096371196e-16 walpha1=1.72079040750854e-21 palpha1=-1.76895188943389e-27
+  beta0=-177.846304375612 lbeta0=0.000196003950840187 wbeta0=9.41133421878783e-05 pbeta0=-9.94424117859599e-11
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-1.05304425311941e-09 lagidl=1.00503649477684e-15 wagidl=6.69374284553109e-16 pagidl=-5.60107774411636e-22
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.592176172339096 lkt1=-1.53472870662801e-08 wkt1=6.96601956010945e-08 pkt1=-2.29221224831813e-14
+  kt2=-0.0790969944556881 lkt2=2.98186195646609e-08 wkt2=1.27842099136216e-08 pkt2=-1.84420437074441e-14
+  at=-251839.851460247 lat=0.375190686705529 wat=0.138122565704439 pat=-1.64186757952069e-7
+  ute=-4.48789203866116 lute=6.18494420653178e-06 wute=1.45381891764711e-06 pute=-2.43511162645319e-12
+  ua1=-4.54665601797395e-09 lua1=9.32721284137611e-15 wua1=1.87246723631851e-15 pua1=-3.86407348209934e-21
+  ub1=4.45772694948955e-18 lub1=-9.28130373080606e-24 wub1=-1.55832219889895e-24 pub1=3.84984865115673e-30
+  uc1=2.0787211949509e-10 luc1=-3.13384908199301e-16 wuc1=-5.97736252458561e-17 puc1=1.13393527254822e-22
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=2.745e-6
+  sbref=2.74e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.104 pmos
* DC IV MOS Parameters
+  lmin=5e-07 lmax=1e-06 wmin=4.2e-07 wmax=5.5e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.889525665814068+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0=-1.02427747476064e-08 wvth0=-7.91448212034604e-08 pvth0=1.84285110949436e-14
+  k1=0.603238458959026 lk1=5.8763110814697e-09 wk1=-9.25581782066799e-08 pk1=2.69075255593331e-14
+  k2=-0.0288760627544941 lk2=-5.57666793040898e-09 wk2=2.46658272835186e-08 pk2=-5.93994231788334e-15
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=285283.684686246 lvsat=-0.0839104259081192 wvsat=-0.108245304932267 pvsat=4.68570458026813e-8
+  ua=-3.97443494142799e-09 lua=8.70012843783389e-16 wua=1.30772681327503e-15 pua=-5.43779179673469e-22
+  ub=2.77119159498454e-18 lub=-3.86262980122309e-25 wub=-7.53810116241494e-25 pub=2.93468266797778e-31
+  uc=5.71460387077809e-11 luc=-2.21201168418071e-17 wuc=-5.07644210964763e-17 puc=1.87922006122556e-23
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=-0.00602715216639765 lu0=4.45716615706696e-09 wu0=6.43430842824463e-09 pu0=-2.67686619925174e-15
+  a0=3.6315066925976 la0=-1.53550776497524e-06 wa0=-1.22409197840869e-06 pa0=7.53984039868143e-13
+  keta=-0.0129908778027087 lketa=4.12521188127327e-08 wketa=1.28085926300466e-08 pketa=-2.7776449938487e-14
+  a1=0.0
+  a2=-2.586933888576 la2=1.78826044996147e-06 wa2=1.37303658034438e-06 pa2=-7.24946837982868e-13
+  ags=0.209281556720716 lags=-3.39747438140794e-07 wags=-8.60179864432211e-08 pags=4.03770958048017e-13
+  b0=-1.56272830956639e-07 lb0=5.92437058602257e-15 wb0=7.8645829054493e-14 pb0=-1.98053663769824e-20
+  b1=2.40684925154549e-06 lb1=-1.27740890347641e-12 wb1=-1.28100398719173e-12 pb1=6.7999344639335e-19
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.178390273289819+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff=7.0401407998778e-09 wvoff=-5.54093260045541e-08 pvoff=4.3873238924596e-15
+  nfactor={0.856087110130421+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor=5.22503502727878e-07 wnfactor=1.75153457352247e-07 pnfactor=-5.81746276709018e-14
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=4.20567936072e-05 lcit=-1.69256023430783e-11 wcit=-1.71629572543047e-11 pcit=9.06183547478585e-18
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.49
+  etab=0.189717944859997 letab=-1.00177243441338e-07 wetab=-2.83194304144749e-07 petab=1.49525948981138e-13
+  dsub=0.349430903910948 ldsub=-9.19338960496078e-08 wdsub=-6.91651784867769e-08 pdsub=7.11009735022648e-14
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=1.10799899993606 lpclm=-2.93632845826269e-07 wpclm=-2.03371056573647e-07 ppclm=1.29665912550737e-13
+  pdiblc1=1.13078485510816 lpdiblc1=-7.48525136364332e-07 wpdiblc1=-2.86468546962106e-07 ppdiblc1=2.87809821119599e-13
+  pdiblc2=0.00284137468502792 lpdiblc2=-2.47886423971249e-09 wpdiblc2=-1.57737061289163e-09 ppdiblc2=1.62151806160524e-15
+  pdiblcb=0.433591436595692 lpdiblcb=-6.77024093723132e-07 wpdiblcb=-3.52604718140128e-07 ppdiblcb=3.62473418991434e-13
+  drout=1.96188892814783 ldrout=-6.3280407062365e-07 wdrout=-5.44798770212372e-07 pdrout=3.08005172648075e-13
+  pscbe1=941136687.264283 lpscbe1=-74.518477235295 wpscbe1=-76.8884695072179 ppscbe1=4.05961892381769e-5
+  pscbe2=4.45126514006198e-08 lpscbe2=-3.66243693925508e-14 wpscbe2=-1.44819886472878e-14 ppscbe2=1.49545330434852e-20
+  pvag=0.0
+  delta=0.01
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=17.5977248012758 lbeta0=-4.91016582530341e-06 wbeta0=-5.82029356555601e-06 pbeta0=3.28816656494152e-12
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-2.03246599267786e-10 lagidl=1.31454704189215e-16 wagidl=1.93008024525202e-16 pagidl=-7.04089754980682e-23
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.710280397833605 lkt1=1.06062439491369e-07 wkt1=9.73754453447931e-08 pkt1=-5.14130666367064e-14
+  kt2=-0.0953472908233255 lkt2=4.65237292270359e-08 wkt2=2.80524705490008e-08 pkt2=-3.41376324214863e-14
+  at=120078.995856369 lat=-0.00713742530978467 wat=-0.0214087711582422 pat=-1.90458033274866e-10
+  ute=3.07093472158738 lute=-1.58543899708259e-06 wute=-1.79065755825956e-06 pute=9.00171257061154e-13
+  ua1=9.24417835983556e-09 lua1=-4.84959940899953e-15 wua1=-4.02160967181413e-15 pua1=2.1949668505381e-21
+  ub1=-9.94912100968526e-18 lub1=5.52876308905013e-24 wub1=4.52142336364696e-24 pub1=-2.40005683019372e-30
+  uc1=-2.25071063967566e-10 luc1=1.31675489082107e-16 wuc1=1.0389391557117e-16 puc1=-5.48547406945908e-23
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.745e-6
+  sbref=1.74e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.105 pmos
* DC IV MOS Parameters
+  lmin=2.5e-07 lmax=5e-07 wmin=4.2e-07 wmax=5.5e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.84084748710978+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0=-3.59442689653262e-08 wvth0=-9.34360190505159e-08 pvth0=2.5974092063815e-14
+  k1=0.652310580953471 lk1=-2.00331804661336e-08 wk1=-8.78483273426215e-08 pk1=2.44207808213207e-14
+  k2=-0.0593001283568993 lk2=1.04868736188737e-08 wk2=2.83332739915483e-08 pk2=-7.87631017036254e-15
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=70622.2415499309 lvsat=0.0294282401305378 wvsat=-0.0411807050315856 pvsat=1.14477418303204e-8
+  ua=-3.13778195670918e-09 lua=4.28270107687672e-16 wua=5.86739540055946e-16 pua=-1.63106551261072e-22
+  ub=2.59202836954875e-18 lub=-2.91666947050918e-25 wub=-4.18137715425344e-25 pub=1.1623726723566e-31
+  uc=3.2147585302442e-11 luc=-8.92123342522901e-18 wuc=-3.20432182145228e-17 puc=8.90763014501876e-24
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=-0.000412370866419993 lu0=1.49262900805436e-09 wu0=2.88148575664113e-09 pu0=-8.01018462517153e-16
+  a0=0.624509423823941 la0=5.21507089700311e-08 wa0=4.30712657488374e-07 pa0=-1.19732950229878e-13
+  keta=0.148658132257956 lketa=-4.40966187111775e-08 wketa=-8.40546669317359e-08 pketa=2.33661887510194e-14
+  a1=0.0
+  a2=1.10720647359648 la2=-1.62201331581259e-7
+  ags=-1.38602246243287 lags=5.02553940324069e-07 wags=1.43341797368734e-06 pags=-3.98472995669395e-13
+  b0=-3.06343235540447e-07 lb0=8.51597433614177e-14 wb0=8.68747504553648e-14 pb0=-2.4150138129586e-20
+  b1=-2.64855234056606e-08 lb1=7.36265768049279e-15 wb1=1.455485281586e-14 pb1=-4.0460744245753e-21
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.0312500269039497+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff=-7.06481436089048e-08 wvoff=-9.94725413041316e-08 pvoff=2.7652172812053e-14
+  nfactor={1.81588987970968+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor=1.57391580232668e-08 wnfactor=1.37217183878385e-07 pnfactor=-3.81447305119846e-14
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=0.49
+  etab=3.57163176063846e-05 letab=-2.73029576987636e-11 wetab=1.1018897441879e-11 petab=-3.06312126207307e-18
+  dsub=-0.328060466287976 ldsub=2.65773417518982e-07 wdsub=1.38330356973554e-07 pdsub=-3.84541792743643e-14
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.457025456605324 lpclm=5.00733733698394e-08 wpclm=8.91537405301201e-08 ppclm=-2.4783670022487e-14
+  pdiblc1=-1.11960378024706 lpdiblc1=4.396530584396e-07 wpdiblc1=5.46231463784684e-07 ppdiblc1=-1.51845792154577e-13
+  pdiblc2=-0.0162210653812238 lpdiblc2=7.58587536598766e-09 wpdiblc2=3.15474122578327e-09 ppdiblc2=-8.7698020387304e-16
+  pdiblcb=-1.54218287319138 lpdiblcb=3.66161032552727e-07 wpdiblcb=7.05209436280256e-07 ppdiblcb=-1.96039760772676e-13
+  drout=1.1321919796254 ldrout=-1.94734038167184e-07 wdrout=8.14318382447382e-08 pdrout=-2.26370738499783e-14
+  pscbe1=800079104.265281 lpscbe1=-0.0417661028166094
+  pscbe2=-6.272960750791e-08 lpscbe2=1.99982564040461e-14 wpscbe2=2.92328672863239e-14 ppscbe2=-8.12638631119062e-21
+  pvag=0.0
+  delta=0.01
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=7.19133571530959 lbeta0=5.84282735417716e-07 wbeta0=8.60485623402909e-07 pbeta0=-2.39204677478528e-13
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-6.9243602569994e-10 lagidl=3.89740851072275e-16 wagidl=1.25987781419777e-16 pagidl=-3.50230913813209e-23
+  bgidl=691592551.5264 lbgidl=162.83543190468
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.506431088159999 lkt1=-1.56754982457793e-9
+  kt2=0.00428747494323944 lkt2=-6.08223148052129e-09 wkt2=-7.73050584050417e-08 pkt2=2.14898785759007e-14
+  at=151044.296905712 lat=-0.0234867326802252 wat=-0.0459761291982913 pat=1.27808122035746e-8
+  ute=0.349922085835547 lute=-1.48776977557252e-07 wute=-1.8109778323677e-07 pute=5.03430105664232e-14
+  ua1=-3.22741818666681e-10 lua1=2.01619642207514e-16 wua1=2.86420812545226e-16 pua1=-7.96215488378224e-23
+  ub1=6.14839413553695e-19 lub1=-4.88812468949642e-26 wub1=-5.11982050739465e-26 pub1=1.42324866320963e-32
+  uc1=5.072625803232e-11 luc1=-1.39421873659686e-17
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.245e-6
+  sbref=1.24e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.106 pmos
* DC IV MOS Parameters
+  lmin=1.8e-07 lmax=2.5e-07 wmin=4.2e-07 wmax=5.5e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.892135672457146+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0=-2.16867688969838e-8
+  k1=-0.614523479319425 lk1=3.32131486281009e-7
+  k2=0.495077243737657 lk2=-1.43623383294948e-07 wk2=2.64697796016969e-23 pk2=6.31088724176809e-30
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=351861.618893142 lvsat=-0.048752931898347
+  ua=9.63598011685708e-10 lua=-7.11864306966488e-16
+  ub=-6.81946012057137e-19 lub=6.18458643342942e-25
+  uc=-3.76598328805701e-15 luc=1.64564159885245e-20
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.0112433187371429 lu0=-1.74751283346087e-9
+  a0=-0.639616527428569 la0=4.03562553906814e-7
+  keta=-0.218982630074297 lketa=5.81031015280409e-08 wketa=-2.64697796016969e-23 pketa=-6.31088724176809e-30
+  a1=0.0
+  a2=0.0932382251080011 la2=1.19669673879557e-7
+  ags=-2.03898102803886 lags=6.84068586059746e-7
+  b0=2.25773945257143e-07 lb0=-6.27624474941426e-14
+  b1=-2.14741667485714e-08 lb1=5.96956066610187e-15
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={0.195503957601713+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff=-1.33683030253665e-7
+  nfactor={4.98966010821143+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor=-8.66530880257478e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=1.57846856239943 leta0=-3.02581198724292e-7
+  etab=0.293574393861143 letab=-8.16275328506713e-08 wetab=-3.05022850878929e-23 petab=3.8087190580202e-30
+  dsub=1.71815201014572 ldsub=-3.03049096379867e-7
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.670335002130859 lpclm=-9.22412057171261e-9
+  pdiblc1=1.33192513110629 lpdiblc1=-2.41842560569694e-7
+  pdiblc2=0.0339036363136343 lpdiblc2=-6.34819020876257e-9
+  pdiblcb=-0.893515669637313 lpdiblcb=1.85839333971137e-7
+  drout=-1.256946487644 ldrout=4.694177860721e-7
+  pscbe1=799717484.766859 lpscbe1=0.0587597783114688
+  pscbe2=3.36027181733886e-08 lpscbe2=-6.78097414744674e-15
+  pvag=0.0
+  delta=0.01
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=12.01765178888 lbeta0=-7.57375217241974e-7
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=2.14542615165143e-09 lagidl=-3.99150779885277e-16 wagidl=-7.88860905221012e-31
+  bgidl=2101455173.12 lbgidl=-229.089458546882
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=0.901713573714284 lkt1=-3.93014868089687e-7
+  kt2=0.286688501485714 lkt2=-8.45863280470108e-08 wkt2=-1.32348898008484e-23 pkt2=6.31088724176809e-30
+  at=-18511.0919999995 lat=0.023647630770896
+  ute=-0.343222029714286 lute=4.39087688362147e-8
+  ua1=1.10675765542857e-09 lua1=-1.95764057597278e-16 wua1=-3.94430452610506e-31
+  ub1=6.36172624000001e-19 lub1=-5.48116234005122e-26
+  uc1=-6.99880644011428e-11 luc1=1.96149456986649e-17 wuc1=-2.31111593326468e-33 puc1=9.18354961579912e-40
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.1e-6
+  sbref=1.1e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8__model.107 pmos
* DC IV MOS Parameters
+  lmin=1.5e-07 lmax=1.8e-07 wmin=4.2e-07 wmax=5.5e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.3994e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=7.3039e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=-2.0e-7
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.76784156345736+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0=-4.75384520396319e-08 wvth0=-6.0948140384743e-08 pvth0=1.26764818223416e-14
+  k1=-4.07900378532117 lk1=1.0527018161657e-06 wk1=1.94253500968166e-06 pk1=-4.04023971593668e-13
+  k2=1.29649356002937 lk2=-3.1030836008783e-07 wk2=-5.26391545977979e-07 pk2=1.09483124864868e-13
+  k3=-15.845
+  dvt0=4.4955
+  dvt1=0.294
+  dvt2=0.015
+  dvt0w=-4.9772
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  w0=0.0
+  k3b=2.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=830171.693055405 lvsat=-0.148235687603207 wvsat=-0.304790229097765 pvsat=6.33927101695859e-8
+  ua=-1.13013872242038e-09 lua=-2.76392191113232e-16 wua=-4.79581531751624e-16 pua=9.97472036259565e-23
+  ub=1.1406395781353e-18 lub=2.39382711609998e-25 wub=2.71629804984974e-25 pub=-5.64957398792145e-32
+  uc=8.38613022801412e-13 luc=-1.58748308730012e-19 wuc=-6.7099385685329e-19 puc=1.39558670299202e-25
+  rdsw=547.88
+  prwb=-0.32348
+  prwg=0.1376
+  wr=1.0
+  u0=0.00851953177556823 lu0=-1.18099783089689e-09 wu0=-2.2951882997804e-09 pu0=4.77371624094727e-16
+  a0=9.35601258824698 la0=-1.67540835460431e-06 wa0=-2.23167762341037e-06 pa0=4.64162165537875e-13
+  keta=1.25740201008753 lketa=-2.48967187009938e-07 wketa=-3.69709775271674e-07 pketa=7.68951967392049e-14
+  a1=0.0
+  a2=-4.87718884908827 la2=1.15345886018749e-06 wa2=2.55181077670244e-06 pa2=-5.30746019824786e-13
+  ags=-14.0213761047436 lags=3.17626297327342e-06 wags=6.19089675612945e-06 pags=-1.28763223451385e-12
+  b0=-2.12154650021876e-06 lb0=4.25452037319499e-13 wb0=7.68215996674591e-13 pb0=-1.59779708716355e-19
+  b1=3.73452524038533e-08 lb1=-6.26417268457264e-15 wb1=-1.17973728584803e-15 pb1=2.45371198608958e-22
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-2.41507012617082+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff=4.09285052282016e-07 wvoff=7.50347285658135e-07 pvoff=-1.56063231249464e-13
+  nfactor={-7.07292750829983+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor=1.64234259292547e-06 wnfactor=-6.24240501714043e-07 pnfactor=1.298345334705e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=1.0e-5
+  cdsc=0.00013
+  cdscb=0.00078
+  cdscd=0.0
+  eta0=-2.10768448899337 leta0=4.64094402128792e-07 weta0=1.01685195923991e-06 peta0=-2.1149300529839e-13
+  etab=-1.00242774536384 letab=1.87925360082455e-07 wetab=2.40489554679903e-07 petab=-5.00189414987637e-14
+  dsub=0.267634130210667 ldsub=-1.35878356793621e-9
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=3.82107240499831 lpclm=-6.64539691519309e-07 wpclm=-1.68372244112318e-06 ppclm=3.50194063084328e-13
+  pdiblc1=2.71046970141515 lpdiblc1=-5.28563288659095e-07 wpdiblc1=-1.38835564837737e-06 ppdiblc1=2.88761314594713e-13
+  pdiblc2=0.06202563151509 lpdiblc2=-1.21972277467229e-08 wpdiblc2=-3.22003398438507e-08 ppdiblc2=6.69728428344282e-15
+  pdiblcb=1.82981488155382 lpdiblcb=-3.80580740710005e-07 wpdiblcb=-7.41456619258789e-07 ppdiblcb=1.54214079326397e-13
+  drout=-0.670911346534268 ldrout=3.4752950914297e-07 wdrout=8.94592901825945e-07 pdrout=-1.86064588464975e-13
+  pscbe1=745143924.105118 lpscbe1=11.4094055132259 wpscbe1=29.3695151567299 ppscbe1=-6.10850671841799e-6
+  pscbe2=-7.30189637019774e-08 lpscbe2=1.53950562224469e-14 wpscbe2=1.29412336499907e-14 ppscbe2=-2.69162130439426e-21
+  pvag=0.0
+  delta=0.01
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=29.926269521579 lbeta0=-4.48215280223057e-06 wbeta0=-9.58105658337296e-06 pbeta0=1.99274479666258e-12
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=-7.82692672324005e-10 lagidl=2.09862798075726e-16 wagidl=-3.54856754072194e-15 pagidl=7.38059465659676e-22
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-5.60745301490793 lkt1=9.60813672344669e-07 wkt1=1.62873083490696e-06 pkt1=-3.3875646889063e-13
+  kt2=-0.12
+  at=416639.166937892 lat=-0.0668584012850783 wat=-0.0560647610235083 pat=1.16607975157574e-8
+  ute=-3.91515044854398 lute=7.86827016811766e-07 wute=1.60577003701783e-06 pute=-3.33980898459265e-13
+  ua1=-1.35143182854246e-10 lua1=6.25364139554892e-17 wua1=2.06528315784479e-16 pua1=-4.29554113433821e-23
+  ub1=3.7264e-19
+  uc1=2.69989354843281e-10 luc1=-5.10962777751443e-17 wuc1=-1.3249509601598e-16 puc1=2.75573900301716e-23
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=1.5e+42
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=1.0
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=8.04e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.0020386
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=5.248925e-11
+  cgso=5.248925e-11
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=9.54827175e-12
+  cgdl=9.54827175e-12
+  cf=1.2e-11
+  clc=1.0e-7
+  cle=0.6
+  dlc=-3.0e-9
+  dwc=0.0
+  vfbcv=-0.14469
+  acde=0.8
+  moin=18.13
+  noff=3.9
+  voffcv=-0.10701
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.0007380194454
+  mjs=0.34629
+  pbs=0.6587
+  cjsws=9.888892e-11
+  mjsws=0.29781
+  pbsws=0.7418
+  cjswgs=2.39155046e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.04e-6
+  sbref=1.04e-6
+  wlod={0+sky130_fd_pr__pfet_01v8__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.ends sky130_fd_pr__pfet_01v8
