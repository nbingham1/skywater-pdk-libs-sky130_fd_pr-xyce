* Capacitor value test

* Include SkyWater sky130 device models
.lib "../../../models/sky130.lib.spice" tt

.param freq=1Meg
.csparam freq={freq}

* Resistor bridge with capacitance
V1 N2 0 1.8
IAC N3 N4 dc 0 ac 1

X1 N3 N4 0 sky130_fd_pr__cap_vpp_02p7x41p1_m1m2m3m4_shieldl1_fingercap
* C34 N3 N4 50E-15

R1 N3 0 1.1Meg
R2 N4 0 1.2Meg
R3 N2 N3 1.3Meg
R4 N2 N4 1.4Meg

.ac lin 1 {freq} {freq}
.control
run
echo capacitance
print imag ( 1/v ( N4,N3 ) ) /2/PI/freq
quit
.endc

.end
