* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param sky130_fd_pr__cap_vpp_04p4x04p6_m1m2_shieldl1__slope=0.0
* statistics {
*   mismatch {
*     vary  sky130_fd_pr__cap_vpp_04p4x04p6_m1m2_shieldl1__slope dist=gauss std=0.00731
*   }
* }
.subckt sky130_fd_pr__cap_vpp_04p4x04p6_m1m2_shieldl1 c0 c1 b
.param mult=1.0
+  ctot_a={8.450e-15*sky130_fd_pr__cap_vpp_04p4x04p6_m1m2_shieldl1__cor+0.88861/sqrt(mult/0.463538)*sky130_fd_pr__cap_vpp_04p4x04p6_m1m2_shieldl1__slope*8.450e-15*sky130_fd_pr__cap_vpp_04p4x04p6_m1m2_shieldl1__cor}
+  cli2s={1.864e-15*cli2s_vpp}
+  rat_m2=0.552
+  rat_m1=0.395
+  rat_m12li=0.053
+  cap_m2={rat_m2*ctot_a}
+  cap_m1={rat_m1*ctot_a}
+  cap_m12li={rat_m12li*ctot_a}
+  lm2=1.585
+  wm2=0.140
+  nfm2=24.0
+  nvia_c0=40.0
+  nvia_c1=18.0
+  lm1=1.665
+  wm1=0.140
+  nfm1=20.0
+  nmcon=42.0
rm21 c0 a1 r={rm2*lm2/wm2*(1/3)*(1/nfm2)}
ccmvpp4p4x4p6_lishield a1 c1 c={cap_m2}
rvia1 c0 d0 r={rcvia/nvia_c0}
rvia2 c1 d1 r={rcvia/nvia_c1}
rm11 d0 b1 r={rm1*lm1/wm1*(1/3)*(1/nfm1)}
cm1 b1 d1 c={cap_m1}
rmcon d0 e0 r={rcl1/nmcon}
rliw e0 f0 r={rl1}
cli2b f0 b c={cli2s}
cm12li d1 f0 c={cap_m12li}
.ends sky130_fd_pr__cap_vpp_04p4x04p6_m1m2_shieldl1
