* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param sky130_fd_pr__nfet_03v3_nvt__toxe_slope=0.45e-2
.param sky130_fd_pr__nfet_03v3_nvt__vth0_slope=0.006 ; All devices
.param sky130_fd_pr__nfet_03v3_nvt__voff_slope=0.0065
.param sky130_fd_pr__nfet_03v3_nvt__nfactor_slope=0
.param sky130_fd_pr__nfet_03v3_nvt__lint_slope=0.0e-9 ; All devices
.param sky130_fd_pr__nfet_03v3_nvt__wint_slope=0.0e-9 ; All devices
