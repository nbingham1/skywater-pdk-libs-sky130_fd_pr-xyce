* SKY130 Spice File.
.options parser scale=1.0u
.include "parameters/lod.spice"
.param
+  lv_dlc_rotweak=.00e-9
+  lvhvt_dlc_rotweak=.00e-9
+  lvt_dlc_rotweak=.00e-9
+  hv_dlc_rotweak=.00e-9
+  sky130_fd_pr__nfet_01v8__dlc_rotweak=lv_dlc_rotweak
+  sky130_fd_pr__esd_nfet_01v8__dlc_rotweak=lv_dlc_rotweak
+  sky130_fd_pr__nfet_01v8_lvt__dlc_rotweak=lvt_dlc_rotweak
+  sky130_fd_pr__pfet_01v8__dlc_rotweak=lv_dlc_rotweak
+  sky130_fd_pr__pfet_01v8_lvt__dlc_rotweak=lvt_dlc_rotweak
+  sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak=lvhvt_dlc_rotweak
+  sky130_fd_pr__esd_nfet_g5v0d10v5__dlc_rotweak=hv_dlc_rotweak
+  sky130_fd_pr__esd_pfet_g5v0d10v5__dlc_rotweak=hv_dlc_rotweak
+  sky130_fd_pr__nfet_03v3_nvt__dlc_rotweak=hv_dlc_rotweak
+  sky130_fd_pr__nfet_05v0_nvt__dlc_rotweak=hv_dlc_rotweak
+  sky130_fd_pr__nfet_g5v0d10v5__dlc_rotweak=hv_dlc_rotweak
+  sky130_fd_pr__pfet_g5v0d10v5__dlc_rotweak=hv_dlc_rotweak
+  sky130_fd_pr__pfet_g5v0d16v0__dlc_rotweak=hv_dlc_rotweak
+  sky130_fd_pr__special_nfet_pass__dlc_rotweak=lv_dlc_rotweak
+  sky130_fd_pr__special_nfet_pass_lowleakage__dlc_rotweak=lv_dlc_rotweak
+  sky130_fd_pr__special_nfet_pass_flash__dlc_rotweak=hv_dlc_rotweak
+  sky130_fd_pr__special_nfet_latch__dlc_rotweak=lv_dlc_rotweak
+  sky130_fd_pr__special_nfet_latch_lowleakage__dlc_rotweak=lv_dlc_rotweak
+  sky130_fd_pr__special_pfet_pass__dlc_rotweak=lv_dlc_rotweak
+  sky130_fd_pr__special_pfet_pass_lowleakage__dlc_rotweak=lv_dlc_rotweak
+  sky130_fd_bs_flash__special_sonosfet_star__dlc_rotweak=hv_dlc_rotweak
+  sky130_fd_bs_flash__special_sonosfet_original__dlc_rotweak=hv_dlc_rotweak
+  sonos_eeol_dlc_rotweak=hv_dlc_rotweak
+  sonos_peol_dlc_rotweak=hv_dlc_rotweak
* include all individual diode models
.include "parasitics/sky130_fd_pr__model__parasitic__diode_ps2nw.model.spice"
.include "../cells/diode_pw2nd_05v5/sky130_fd_pr__diode_pw2nd_05v5.model.spice"
.include "../cells/diode_pd2nw_05v5/sky130_fd_pr__diode_pd2nw_05v5.model.spice"
.include "../cells/diode_pd2nw_05v5_hvt/sky130_fd_pr__diode_pd2nw_05v5_hvt.model.spice"
.include "../cells/diode_pw2nd_11v0/sky130_fd_pr__diode_pw2nd_11v0.model.spice"
.include "../cells/diode_pd2nw_11v0/sky130_fd_pr__diode_pd2nw_11v0.model.spice"
.include "../cells/diode_pw2nd_05v5_nvt/sky130_fd_pr__diode_pw2nd_05v5_nvt.model.spice"
.include "../cells/diode_pw2nd_05v5_lvt/sky130_fd_pr__diode_pw2nd_05v5_lvt.model.spice"
.include "../cells/diode_pd2nw_05v5_lvt/sky130_fd_pr__diode_pd2nw_05v5_lvt.model.spice"
.include "parasitics/sky130_fd_pr__model__parasitic__diode_pw2dn.model.spice"
.include "parasitics/sky130_fd_pr__model__parasitic__diode_ps2dn.model.spice"
.include "../cells/pfet_g5v0d16v0/sky130_fd_pr__pfet_g5v0d16v0__parasitic__diode_pw2dn.model.spice"
* call models applicable to any corner
.include "../cells/pnp_05v5/sky130_fd_pr__pnp_05v5_W0p68L0p68.model.spice"
.include "../cells/pfet_g5v0d16v0/sky130_fd_pr__pfet_g5v0d16v0.pm3.spice"
.include "../cells/pfet_g5v0d16v0/sky130_fd_pr__pfet_g5v0d16v0__subcircuit.pm3.spice"
.include "../cells/cap_var_lvt/sky130_fd_pr__cap_var_lvt.model.spice"
.include "../cells/res_iso_pw/sky130_fd_pr__res_iso_pw.model.spice"
.include "../cells/cap_vpp_08p6x07p8_l1m1m2_noshield/sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_noshield_o1.model.spice"
.include "capacitors/sky130_fd_pr__model__cap_mim.model.spice"
.include "capacitors/sky130_fd_pr__model__cap_vpp_only_mos.model.spice"
.include "sonos_p/begin_of_life/mm.spice"
.include "sonos_e/begin_of_life/mm.spice"
*.include "hspice.par"
.include "head.spice"
.include "../cells/special_nfet_pass/sky130_fd_pr__special_nfet_pass.pm3.spice"
.include "../cells/special_nfet_latch/sky130_fd_pr__special_nfet_latch.pm3.spice"
.include "../cells/special_pfet_pass/sky130_fd_pr__special_pfet_pass.pm3.spice"
.include "../cells/special_nfet_pass_flash/sky130_fd_pr__special_nfet_pass_flash.pm3.spice"
.include "capacitors/sky130_fd_pr__model__cap_vpp_only_pq.model.spice"
.include "capacitors/sky130_fd_pr__model__cap_vpp_only_p.model.spice"
.include "sky130_fd_pr__model__linear.model.spice"
.param sky130_fd_pr__rf_nfet_01v8_lvt__base__dlc_rotweak=0
.param sky130_fd_pr__pfet_01v8_lvt__rf_base_dlc_rotweak=0
.param sky130_fd_pr__rf_nfet_01v8__base__dlc_rotweak=0
.param sky130_fd_pr__rf_pfet_01v8__base__dlc_rotweak=0
.param sky130_fd_pr__rf_nfet_g5v0d10v5__base__dlc_rotweak=0
.include "../cells/rf_nfet_g5v0d10v5/sky130_fd_pr__rf_nfet_g5v0d10v5.pm3.spice"
.include "../cells/rf_nfet_01v8_lvt/sky130_fd_pr__rf_nfet_01v8_lvt.pm3.spice"
.include "../cells/rf_nfet_01v8/sky130_fd_pr__rf_nfet_01v8.pm3.spice"
.include "../cells/rf_pfet_01v8/sky130_fd_pr__rf_pfet_01v8.pm3.spice"
.include "../cells/rf_pfet_01v8_mvt/sky130_fd_pr__rf_pfet_01v8_mvt.pm3.spice"
