* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param sky130_fd_pr__cap_vpp_04p4x04p6_m1m2_noshield_o1phv__slope=0.0
* statistics {
*   mismatch {
*     vary  sky130_fd_pr__cap_vpp_04p4x04p6_m1m2_noshield_o1phv__slope dist=gauss std=0.00914
*   }
* }
.subckt sky130_fd_pr__cap_vpp_04p4x04p6_m1m2_noshield_o1phv c0 c1 b
.param mult=1.0
+  lvpp=3.6 wm1=0.14 wm2=0.14 wli=0.17
+  ctot_a={0.988e-15*lvpp*lvpp*cvpp2_phv5x4_cor+1.04204/sqrt(mult/0.35036)*sky130_fd_pr__cap_vpp_04p4x04p6_m1m2_noshield_o1phv__slope*0.988e-15*lvpp*lvpp*cvpp2_phv5x4_cor}
+  rat_m2=0.4325
+  rat_m1=0.3175
+  rat_li=0.25
+  cap_m2={rat_m2*ctot_a}
+  cap_m1={rat_m1*ctot_a}
+  cap_li={rat_li*ctot_a}
+  caps_li={cvpp2_phv5x4_sub}
+  nvia=11.0
+  ncon=10.0
+  nf=6.0
rm21 c0 a1 r={2*rm2*lvpp/wm2*(1/3)*(1/nf)}
ccmvpp2_phv5x4 a1 c1 c={cap_m2}
rvia1 c0 d0 r={rcvia/nvia}
rvia2 c1 d1 r={rcvia/nvia}
rm11 d0 b1 r={2*rm1*lvpp/wm1*(1/3)*(1/nf)}
cm1 b1 d1 c={cap_m1}
rcon1 d0 e0 r={rcl1/ncon}
rcon2 d1 e1 r={rcl1/ncon}
rli1 e0 f1 r={2*rl1*lvpp/wli*(1/3)*(1/nf)}
cli f1 e1 c={cap_li}
csli1 e0 b c={caps_li}
csli2 e1 b c={caps_li}
.ends sky130_fd_pr__cap_vpp_04p4x04p6_m1m2_noshield_o1phv
