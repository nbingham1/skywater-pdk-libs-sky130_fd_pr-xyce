* Inductor value test

* Include SkyWater sky130 device models
.include "../../../models/sky130_fd_pr__model__inductors.model.spice"

.param lofreq=1Meg
.csparam lofreq={lofreq}
.param hifreq=10G
.csparam hifreq={hifreq}

V1 N2 0 1.8
IAC N2 N3 dc 0 ac 1

* L-C tank with ideal capacitor
X1 N3 N4 mid 0 sky130_fd_pr__ind_03_90
C34 N3 N4 1.0E-10
R1 N4 0 100

.ac dec 100 {lofreq} {hifreq}
.control
run
echo inductance
let resp=mag(v(N4,N3))
meas ac ymax max_at resp
* Note: 39.478 is (2*pi)^2
let l=1/(1.0E-10*39.478*ymax*ymax)
print l
quit
.endc

.end
