* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 40
.param
+  sky130_fd_pr__pfet_01v8_lvt__toxe_mult=0.948
+  sky130_fd_pr__pfet_01v8_lvt__rshp_mult=1.0
+  sky130_fd_pr__pfet_01v8_lvt__overlap_mult=0.1
+  sky130_fd_pr__pfet_01v8_lvt__ajunction_mult=9.0161e-1
+  sky130_fd_pr__pfet_01v8_lvt__pjunction_mult=9.0587e-1
+  sky130_fd_pr__pfet_01v8_lvt__lint_diff=1.7325e-8
+  sky130_fd_pr__pfet_01v8_lvt__wint_diff=-3.2175e-8
+  sky130_fd_pr__pfet_01v8_lvt__dlc_diff=3.417e-8
+  sky130_fd_pr__pfet_01v8_lvt__dwc_diff=-3.2175e-8
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 000, W = 1.0, L = 1.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8_lvt__agidl_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_lvt__u0_diff_0=-0.00018933
+  sky130_fd_pr__pfet_01v8_lvt__pdits_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ua_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_lvt__vsat_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_lvt__b1_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_lvt__kt1_diff_0=-0.23862
+  sky130_fd_pr__pfet_01v8_lvt__pclm_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_lvt__eta0_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ub_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ags_diff_0=-0.051202
+  sky130_fd_pr__pfet_01v8_lvt__keta_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_lvt__vth0_diff_0=0.11022
+  sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_lvt__voff_diff_0=0.06319
+  sky130_fd_pr__pfet_01v8_lvt__a0_diff_0=0.13279
+  sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_0=-0.14855
+  sky130_fd_pr__pfet_01v8_lvt__b0_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_lvt__k2_diff_0=0.07564
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 001, W = 1.0, L = 2.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_1=0.10795
+  sky130_fd_pr__pfet_01v8_lvt__voff_diff_1=-0.0069915
+  sky130_fd_pr__pfet_01v8_lvt__b0_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_lvt__k2_diff_1=0.047653
+  sky130_fd_pr__pfet_01v8_lvt__agidl_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_lvt__u0_diff_1=-0.00011306
+  sky130_fd_pr__pfet_01v8_lvt__pdits_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ua_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_lvt__vsat_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_lvt__b1_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_lvt__kt1_diff_1=-0.29418
+  sky130_fd_pr__pfet_01v8_lvt__pclm_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_lvt__eta0_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ub_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ags_diff_1=-0.020877
+  sky130_fd_pr__pfet_01v8_lvt__keta_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_lvt__vth0_diff_1=0.11014
+  sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_lvt__a0_diff_1=0.11885
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 002, W = 1.0, L = 4.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_lvt__a0_diff_2=0.12779
+  sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_2=0.23595
+  sky130_fd_pr__pfet_01v8_lvt__voff_diff_2=-0.059291
+  sky130_fd_pr__pfet_01v8_lvt__b0_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_lvt__k2_diff_2=0.051303
+  sky130_fd_pr__pfet_01v8_lvt__agidl_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_lvt__u0_diff_2=-0.00019291
+  sky130_fd_pr__pfet_01v8_lvt__ua_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_lvt__vsat_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pdits_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_lvt__b1_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_lvt__kt1_diff_2=-0.29708
+  sky130_fd_pr__pfet_01v8_lvt__pclm_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_lvt__eta0_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ub_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ags_diff_2=-0.10828
+  sky130_fd_pr__pfet_01v8_lvt__keta_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_lvt__vth0_diff_2=0.1166
+  sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_2=0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 003, W = 1.0, L = 8.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_lvt__a0_diff_3=0.12606
+  sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_3=0.1086
+  sky130_fd_pr__pfet_01v8_lvt__voff_diff_3=-0.033808
+  sky130_fd_pr__pfet_01v8_lvt__b0_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_lvt__k2_diff_3=0.053159
+  sky130_fd_pr__pfet_01v8_lvt__agidl_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_lvt__u0_diff_3=-0.0001103
+  sky130_fd_pr__pfet_01v8_lvt__ua_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_lvt__vsat_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pdits_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_lvt__b1_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_lvt__kt1_diff_3=-0.40981
+  sky130_fd_pr__pfet_01v8_lvt__pclm_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_lvt__eta0_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ub_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ags_diff_3=-0.062196
+  sky130_fd_pr__pfet_01v8_lvt__keta_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_lvt__vth0_diff_3=0.11157
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 004, W = 1.0, L = 0.35
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_lvt__vth0_diff_4=0.23648
+  sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_lvt__a0_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_4=8.0
+  sky130_fd_pr__pfet_01v8_lvt__voff_diff_4=-0.45
+  sky130_fd_pr__pfet_01v8_lvt__b0_diff_4=4.3243e-8
+  sky130_fd_pr__pfet_01v8_lvt__k2_diff_4=0.11582
+  sky130_fd_pr__pfet_01v8_lvt__agidl_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_lvt__u0_diff_4=-0.00095521
+  sky130_fd_pr__pfet_01v8_lvt__ua_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_lvt__vsat_diff_4=51751.0
+  sky130_fd_pr__pfet_01v8_lvt__pdits_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_lvt__b1_diff_4=2.0324e-7
+  sky130_fd_pr__pfet_01v8_lvt__kt1_diff_4=-0.52086
+  sky130_fd_pr__pfet_01v8_lvt__pclm_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_lvt__eta0_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ub_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ags_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_lvt__keta_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_4=0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 005, W = 1.0, L = 0.5
* ---------------------------------
+  sky130_fd_pr__pfet_01v8_lvt__keta_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_lvt__vth0_diff_5=0.1966
+  sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_lvt__a0_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_5=-0.80325
+  sky130_fd_pr__pfet_01v8_lvt__voff_diff_5=0.081339
+  sky130_fd_pr__pfet_01v8_lvt__b0_diff_5=4.3678e-7
+  sky130_fd_pr__pfet_01v8_lvt__k2_diff_5=0.060869
+  sky130_fd_pr__pfet_01v8_lvt__agidl_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_lvt__u0_diff_5=-0.00037073
+  sky130_fd_pr__pfet_01v8_lvt__ua_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_lvt__vsat_diff_5=-32446.0
+  sky130_fd_pr__pfet_01v8_lvt__pdits_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_lvt__b1_diff_5=4.8211e-7
+  sky130_fd_pr__pfet_01v8_lvt__kt1_diff_5=-0.52796
+  sky130_fd_pr__pfet_01v8_lvt__pclm_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_lvt__eta0_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ub_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ags_diff_5=0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 006, W = 3.0, L = 1.5
* ---------------------------------
+  sky130_fd_pr__pfet_01v8_lvt__eta0_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ags_diff_6=0.12095
+  sky130_fd_pr__pfet_01v8_lvt__keta_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_lvt__vth0_diff_6=0.090316
+  sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_lvt__a0_diff_6=0.092751
+  sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_6=0.05588
+  sky130_fd_pr__pfet_01v8_lvt__voff_diff_6=0.019108
+  sky130_fd_pr__pfet_01v8_lvt__b0_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_lvt__k2_diff_6=0.045543
+  sky130_fd_pr__pfet_01v8_lvt__agidl_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_lvt__u0_diff_6=-0.00041554
+  sky130_fd_pr__pfet_01v8_lvt__ua_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_lvt__vsat_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pdits_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_lvt__b1_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_lvt__kt1_diff_6=-0.2147
+  sky130_fd_pr__pfet_01v8_lvt__pclm_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ub_diff_6=0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 007, W = 3.0, L = 1.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8_lvt__pclm_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ub_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_lvt__eta0_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ags_diff_7=0.058371
+  sky130_fd_pr__pfet_01v8_lvt__keta_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_lvt__vth0_diff_7=0.080156
+  sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_lvt__a0_diff_7=0.10788
+  sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_7=-0.090095
+  sky130_fd_pr__pfet_01v8_lvt__voff_diff_7=0.021242
+  sky130_fd_pr__pfet_01v8_lvt__b0_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_lvt__k2_diff_7=0.073455
+  sky130_fd_pr__pfet_01v8_lvt__agidl_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_lvt__u0_diff_7=-0.0003142
+  sky130_fd_pr__pfet_01v8_lvt__ua_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_lvt__uc_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_lvt__vsat_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pdits_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_lvt__b1_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_lvt__kt1_diff_7=-0.35565
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 008, W = 3.0, L = 2.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8_lvt__kt1_diff_8=-0.24421
+  sky130_fd_pr__pfet_01v8_lvt__pclm_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ub_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_lvt__eta0_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ags_diff_8=0.070133
+  sky130_fd_pr__pfet_01v8_lvt__keta_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_lvt__vth0_diff_8=0.13775
+  sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_lvt__a0_diff_8=0.099781
+  sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_8=-0.022398
+  sky130_fd_pr__pfet_01v8_lvt__voff_diff_8=0.047981
+  sky130_fd_pr__pfet_01v8_lvt__b0_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_lvt__k2_diff_8=0.054904
+  sky130_fd_pr__pfet_01v8_lvt__agidl_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_lvt__u0_diff_8=-0.00047282
+  sky130_fd_pr__pfet_01v8_lvt__ua_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_lvt__vsat_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pdits_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_lvt__b1_diff_8=0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 009, W = 3.0, L = 4.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8_lvt__pdits_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_lvt__b1_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_lvt__kt1_diff_9=-0.25403
+  sky130_fd_pr__pfet_01v8_lvt__pclm_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ub_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_lvt__eta0_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ags_diff_9=0.076884
+  sky130_fd_pr__pfet_01v8_lvt__keta_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_lvt__vth0_diff_9=0.12658
+  sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_lvt__a0_diff_9=0.098398
+  sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_9=0.020287
+  sky130_fd_pr__pfet_01v8_lvt__voff_diff_9=0.013952
+  sky130_fd_pr__pfet_01v8_lvt__b0_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_lvt__k2_diff_9=0.057134
+  sky130_fd_pr__pfet_01v8_lvt__agidl_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_lvt__u0_diff_9=-0.0004462
+  sky130_fd_pr__pfet_01v8_lvt__ua_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_lvt__vsat_diff_9=0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 010, W = 3.0, L = 8.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8_lvt__u0_diff_10=-0.00043243
+  sky130_fd_pr__pfet_01v8_lvt__vsat_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_lvt__vth0_diff_10=0.12893
+  sky130_fd_pr__pfet_01v8_lvt__keta_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ua_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pclm_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_lvt__kt1_diff_10=-0.32854
+  sky130_fd_pr__pfet_01v8_lvt__b0_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pdits_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_lvt__b1_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_lvt__agidl_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_10=0.074913
+  sky130_fd_pr__pfet_01v8_lvt__ub_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_lvt__k2_diff_10=0.046913
+  sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_lvt__voff_diff_10=-0.00058355
+  sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_lvt__eta0_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ags_diff_10=0.023555
+  sky130_fd_pr__pfet_01v8_lvt__a0_diff_10=0.10527
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 011, W = 3.0, L = 0.35
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_lvt__eta0_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ags_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_lvt__a0_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_lvt__u0_diff_11=-0.0011267
+  sky130_fd_pr__pfet_01v8_lvt__vsat_diff_11=96214.0
+  sky130_fd_pr__pfet_01v8_lvt__vth0_diff_11=0.17584
+  sky130_fd_pr__pfet_01v8_lvt__keta_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ua_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pclm_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_lvt__kt1_diff_11=-0.60261
+  sky130_fd_pr__pfet_01v8_lvt__b0_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pdits_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_lvt__b1_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_lvt__agidl_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_11=8.0
+  sky130_fd_pr__pfet_01v8_lvt__ub_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_lvt__k2_diff_11=0.091919
+  sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_lvt__voff_diff_11=-0.45
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 012, W = 3.0, L = 0.5
* ---------------------------------
+  sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_lvt__voff_diff_12=-0.025789
+  sky130_fd_pr__pfet_01v8_lvt__k2_diff_12=0.035523
+  sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_lvt__eta0_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ags_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_lvt__a0_diff_12=0.095072
+  sky130_fd_pr__pfet_01v8_lvt__u0_diff_12=-0.00054776
+  sky130_fd_pr__pfet_01v8_lvt__vsat_diff_12=-19485.0
+  sky130_fd_pr__pfet_01v8_lvt__vth0_diff_12=0.098837
+  sky130_fd_pr__pfet_01v8_lvt__keta_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ua_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pclm_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_lvt__kt1_diff_12=-0.63957
+  sky130_fd_pr__pfet_01v8_lvt__b0_diff_12=-2.1123e-7
+  sky130_fd_pr__pfet_01v8_lvt__pdits_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_lvt__b1_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_lvt__agidl_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_12=0.055068
+  sky130_fd_pr__pfet_01v8_lvt__ub_diff_12=0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 013, W = 5.0, L = 1.5
* ---------------------------------
+  sky130_fd_pr__pfet_01v8_lvt__agidl_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_13=-0.064147
+  sky130_fd_pr__pfet_01v8_lvt__ub_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_lvt__voff_diff_13=0.035765
+  sky130_fd_pr__pfet_01v8_lvt__k2_diff_13=0.053005
+  sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_lvt__eta0_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ags_diff_13=-0.095668
+  sky130_fd_pr__pfet_01v8_lvt__a0_diff_13=0.10862
+  sky130_fd_pr__pfet_01v8_lvt__u0_diff_13=-0.00037409
+  sky130_fd_pr__pfet_01v8_lvt__vsat_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_lvt__vth0_diff_13=0.12353
+  sky130_fd_pr__pfet_01v8_lvt__keta_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ua_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pclm_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_lvt__kt1_diff_13=-0.21665
+  sky130_fd_pr__pfet_01v8_lvt__b0_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pdits_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_lvt__b1_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_13=0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 014, W = 5.0, L = 1.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_lvt__agidl_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_14=0.04799
+  sky130_fd_pr__pfet_01v8_lvt__ub_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_lvt__voff_diff_14=0.0090418
+  sky130_fd_pr__pfet_01v8_lvt__k2_diff_14=0.048649
+  sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_lvt__eta0_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ags_diff_14=-0.11234
+  sky130_fd_pr__pfet_01v8_lvt__a0_diff_14=0.12656
+  sky130_fd_pr__pfet_01v8_lvt__u0_diff_14=-0.00026832
+  sky130_fd_pr__pfet_01v8_lvt__vsat_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_lvt__vth0_diff_14=0.088094
+  sky130_fd_pr__pfet_01v8_lvt__keta_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ua_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pclm_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_lvt__kt1_diff_14=-0.27128
+  sky130_fd_pr__pfet_01v8_lvt__b0_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pdits_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_lvt__b1_diff_14=0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 015, W = 5.0, L = 2.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8_lvt__pdits_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_lvt__b1_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_lvt__agidl_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_15=-0.18945
+  sky130_fd_pr__pfet_01v8_lvt__ub_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_lvt__voff_diff_15=0.071071
+  sky130_fd_pr__pfet_01v8_lvt__k2_diff_15=0.061291
+  sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_lvt__eta0_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ags_diff_15=-0.07987
+  sky130_fd_pr__pfet_01v8_lvt__a0_diff_15=0.11171
+  sky130_fd_pr__pfet_01v8_lvt__u0_diff_15=-0.00044527
+  sky130_fd_pr__pfet_01v8_lvt__vsat_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_lvt__vth0_diff_15=0.15954
+  sky130_fd_pr__pfet_01v8_lvt__keta_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ua_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pclm_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_lvt__kt1_diff_15=-0.24517
+  sky130_fd_pr__pfet_01v8_lvt__b0_diff_15=0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 016, W = 5.0, L = 4.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8_lvt__kt1_diff_16=-0.25356
+  sky130_fd_pr__pfet_01v8_lvt__b0_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pdits_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_lvt__b1_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_lvt__agidl_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ub_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_16=0.037134
+  sky130_fd_pr__pfet_01v8_lvt__voff_diff_16=0.015802
+  sky130_fd_pr__pfet_01v8_lvt__k2_diff_16=0.062116
+  sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_lvt__eta0_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ags_diff_16=-0.017309
+  sky130_fd_pr__pfet_01v8_lvt__a0_diff_16=0.10722
+  sky130_fd_pr__pfet_01v8_lvt__u0_diff_16=-0.00035119
+  sky130_fd_pr__pfet_01v8_lvt__vsat_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_lvt__vth0_diff_16=0.13305
+  sky130_fd_pr__pfet_01v8_lvt__keta_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ua_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pclm_diff_16=0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 017, W = 5.0, L = 8.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8_lvt__pclm_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_lvt__kt1_diff_17=-0.41635
+  sky130_fd_pr__pfet_01v8_lvt__b0_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pdits_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_lvt__b1_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_lvt__agidl_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ub_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_17=0.062702
+  sky130_fd_pr__pfet_01v8_lvt__voff_diff_17=0.00095753
+  sky130_fd_pr__pfet_01v8_lvt__k2_diff_17=0.051507
+  sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_lvt__eta0_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ags_diff_17=0.0039705
+  sky130_fd_pr__pfet_01v8_lvt__a0_diff_17=0.10653
+  sky130_fd_pr__pfet_01v8_lvt__u0_diff_17=-0.00035511
+  sky130_fd_pr__pfet_01v8_lvt__vsat_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_lvt__vth0_diff_17=0.13008
+  sky130_fd_pr__pfet_01v8_lvt__keta_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ua_diff_17=0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 018, W = 5.0, L = 0.35
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_lvt__ua_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pclm_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_lvt__kt1_diff_18=-0.43258
+  sky130_fd_pr__pfet_01v8_lvt__b0_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pdits_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_lvt__b1_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_lvt__agidl_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ub_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_18=8.0
+  sky130_fd_pr__pfet_01v8_lvt__voff_diff_18=-0.45
+  sky130_fd_pr__pfet_01v8_lvt__k2_diff_18=0.072545
+  sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_lvt__eta0_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ags_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_lvt__a0_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_lvt__u0_diff_18=-0.00086413
+  sky130_fd_pr__pfet_01v8_lvt__vsat_diff_18=8387.2
+  sky130_fd_pr__pfet_01v8_lvt__vth0_diff_18=0.12199
+  sky130_fd_pr__pfet_01v8_lvt__keta_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_18=0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 019, W = 5.0, L = 0.5
* ---------------------------------
+  sky130_fd_pr__pfet_01v8_lvt__keta_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ua_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pclm_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_lvt__kt1_diff_19=-0.53131
+  sky130_fd_pr__pfet_01v8_lvt__b0_diff_19=4.4057e-7
+  sky130_fd_pr__pfet_01v8_lvt__pdits_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_lvt__b1_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_lvt__agidl_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ub_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_19=0.078897
+  sky130_fd_pr__pfet_01v8_lvt__voff_diff_19=-0.021945
+  sky130_fd_pr__pfet_01v8_lvt__k2_diff_19=0.035497
+  sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_lvt__eta0_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ags_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_lvt__a0_diff_19=0.11429
+  sky130_fd_pr__pfet_01v8_lvt__u0_diff_19=-0.00039722
+  sky130_fd_pr__pfet_01v8_lvt__vsat_diff_19=-23382.0
+  sky130_fd_pr__pfet_01v8_lvt__vth0_diff_19=0.083283
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 020, W = 7.0, L = 1.5
* ---------------------------------
+  sky130_fd_pr__pfet_01v8_lvt__keta_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ua_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pclm_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_lvt__kt1_diff_20=-0.25477
+  sky130_fd_pr__pfet_01v8_lvt__b0_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pdits_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_lvt__b1_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_lvt__agidl_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_20=0.088389
+  sky130_fd_pr__pfet_01v8_lvt__ub_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_lvt__k2_diff_20=0.039247
+  sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_lvt__voff_diff_20=0.0063659
+  sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_lvt__eta0_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ags_diff_20=0.0051686
+  sky130_fd_pr__pfet_01v8_lvt__a0_diff_20=0.12399
+  sky130_fd_pr__pfet_01v8_lvt__u0_diff_20=-0.0003164
+  sky130_fd_pr__pfet_01v8_lvt__vsat_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_lvt__vth0_diff_20=0.089169
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 021, W = 7.0, L = 1.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8_lvt__u0_diff_21=-0.00034756
+  sky130_fd_pr__pfet_01v8_lvt__vsat_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_lvt__vth0_diff_21=0.08408
+  sky130_fd_pr__pfet_01v8_lvt__keta_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ua_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_lvt__uc_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pclm_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_lvt__kt1_diff_21=-0.32092
+  sky130_fd_pr__pfet_01v8_lvt__b0_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pdits_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_lvt__b1_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_lvt__agidl_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_21=0.085842
+  sky130_fd_pr__pfet_01v8_lvt__ub_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_lvt__k2_diff_21=0.063334
+  sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_lvt__voff_diff_21=0.0086499
+  sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_lvt__eta0_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ags_diff_21=-0.029768
+  sky130_fd_pr__pfet_01v8_lvt__a0_diff_21=0.12577
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 022, W = 7.0, L = 2.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_lvt__eta0_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ags_diff_22=0.090995
+  sky130_fd_pr__pfet_01v8_lvt__a0_diff_22=0.099945
+  sky130_fd_pr__pfet_01v8_lvt__u0_diff_22=-0.00026521
+  sky130_fd_pr__pfet_01v8_lvt__vsat_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_lvt__vth0_diff_22=0.085914
+  sky130_fd_pr__pfet_01v8_lvt__keta_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ua_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pclm_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_lvt__kt1_diff_22=-0.21994
+  sky130_fd_pr__pfet_01v8_lvt__b0_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pdits_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_lvt__b1_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_lvt__agidl_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_22=0.07581
+  sky130_fd_pr__pfet_01v8_lvt__ub_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_lvt__uc_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_lvt__k2_diff_22=0.069356
+  sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_lvt__voff_diff_22=-0.010347
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 023, W = 7.0, L = 4.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_lvt__voff_diff_23=0.012934
+  sky130_fd_pr__pfet_01v8_lvt__k2_diff_23=0.053103
+  sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_lvt__eta0_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ags_diff_23=-0.057499
+  sky130_fd_pr__pfet_01v8_lvt__a0_diff_23=0.11225
+  sky130_fd_pr__pfet_01v8_lvt__u0_diff_23=-0.00030034
+  sky130_fd_pr__pfet_01v8_lvt__vsat_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_lvt__vth0_diff_23=0.12349
+  sky130_fd_pr__pfet_01v8_lvt__keta_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ua_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pclm_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_lvt__kt1_diff_23=-0.27418
+  sky130_fd_pr__pfet_01v8_lvt__b0_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pdits_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_lvt__b1_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_lvt__agidl_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_23=0.072834
+  sky130_fd_pr__pfet_01v8_lvt__ub_diff_23=0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 024, W = 7.0, L = 8.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8_lvt__agidl_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_24=0.0038305
+  sky130_fd_pr__pfet_01v8_lvt__ub_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_lvt__voff_diff_24=0.027527
+  sky130_fd_pr__pfet_01v8_lvt__k2_diff_24=0.050677
+  sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_lvt__eta0_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ags_diff_24=-0.037406
+  sky130_fd_pr__pfet_01v8_lvt__a0_diff_24=0.10942
+  sky130_fd_pr__pfet_01v8_lvt__u0_diff_24=-0.00027269
+  sky130_fd_pr__pfet_01v8_lvt__vsat_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_lvt__vth0_diff_24=0.12024
+  sky130_fd_pr__pfet_01v8_lvt__keta_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ua_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pclm_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_lvt__kt1_diff_24=-0.37048
+  sky130_fd_pr__pfet_01v8_lvt__b0_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pdits_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_lvt__b1_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_24=0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 025, W = 7.0, L = 0.35
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_lvt__agidl_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_25=8.0
+  sky130_fd_pr__pfet_01v8_lvt__ub_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_lvt__voff_diff_25=-0.45
+  sky130_fd_pr__pfet_01v8_lvt__k2_diff_25=0.078624
+  sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_lvt__eta0_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ags_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_lvt__a0_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_lvt__u0_diff_25=-0.0010475
+  sky130_fd_pr__pfet_01v8_lvt__vsat_diff_25=65650.0
+  sky130_fd_pr__pfet_01v8_lvt__vth0_diff_25=0.12236
+  sky130_fd_pr__pfet_01v8_lvt__keta_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ua_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pclm_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_lvt__kt1_diff_25=-0.41395
+  sky130_fd_pr__pfet_01v8_lvt__b0_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pdits_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_lvt__b1_diff_25=0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 026, W = 7.0, L = 0.5
* ---------------------------------
+  sky130_fd_pr__pfet_01v8_lvt__pdits_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_lvt__b1_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_lvt__agidl_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_26=0.1125
+  sky130_fd_pr__pfet_01v8_lvt__ub_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_lvt__voff_diff_26=-0.057692
+  sky130_fd_pr__pfet_01v8_lvt__k2_diff_26=0.037596
+  sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_lvt__eta0_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ags_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_lvt__a0_diff_26=0.09606
+  sky130_fd_pr__pfet_01v8_lvt__u0_diff_26=-0.00035609
+  sky130_fd_pr__pfet_01v8_lvt__vsat_diff_26=-19372.0
+  sky130_fd_pr__pfet_01v8_lvt__vth0_diff_26=0.071633
+  sky130_fd_pr__pfet_01v8_lvt__keta_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ua_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pclm_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_lvt__kt1_diff_26=-0.54124
+  sky130_fd_pr__pfet_01v8_lvt__b0_diff_26=-7.8239e-8
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 027, W = 0.42, L = 1.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_lvt__kt1_diff_27=-0.20686
+  sky130_fd_pr__pfet_01v8_lvt__b0_diff_27=1.8119e-7
+  sky130_fd_pr__pfet_01v8_lvt__pdits_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_lvt__b1_diff_27=3.2805e-7
+  sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_lvt__agidl_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ub_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_27=-0.14655
+  sky130_fd_pr__pfet_01v8_lvt__voff_diff_27=0.06188
+  sky130_fd_pr__pfet_01v8_lvt__k2_diff_27=0.07356
+  sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_lvt__eta0_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ags_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_lvt__a0_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_lvt__u0_diff_27=5.4948e-5
+  sky130_fd_pr__pfet_01v8_lvt__vsat_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_lvt__vth0_diff_27=0.091519
+  sky130_fd_pr__pfet_01v8_lvt__keta_diff_27=-0.008
+  sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ua_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pclm_diff_27=0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 028, W = 0.42, L = 20.0
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_lvt__pclm_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_lvt__kt1_diff_28=-0.40367
+  sky130_fd_pr__pfet_01v8_lvt__b0_diff_28=-2.5405e-8
+  sky130_fd_pr__pfet_01v8_lvt__pdits_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_lvt__b1_diff_28=4.753e-7
+  sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_lvt__agidl_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ub_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_28=4.1916
+  sky130_fd_pr__pfet_01v8_lvt__voff_diff_28=-0.24899
+  sky130_fd_pr__pfet_01v8_lvt__k2_diff_28=0.024556
+  sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_lvt__eta0_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ags_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_lvt__a0_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_lvt__u0_diff_28=-0.00024467
+  sky130_fd_pr__pfet_01v8_lvt__vsat_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_lvt__vth0_diff_28=0.069986
+  sky130_fd_pr__pfet_01v8_lvt__keta_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ua_diff_28=0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 029, W = 0.42, L = 2.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_lvt__ua_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pclm_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_lvt__kt1_diff_29=-0.26031
+  sky130_fd_pr__pfet_01v8_lvt__b0_diff_29=1.0733e-7
+  sky130_fd_pr__pfet_01v8_lvt__pdits_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_lvt__b1_diff_29=1.6884e-7
+  sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_lvt__agidl_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ub_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_29=0.082548
+  sky130_fd_pr__pfet_01v8_lvt__voff_diff_29=0.0083437
+  sky130_fd_pr__pfet_01v8_lvt__k2_diff_29=0.042789
+  sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_lvt__eta0_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ags_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_lvt__a0_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_lvt__u0_diff_29=-0.00026374
+  sky130_fd_pr__pfet_01v8_lvt__vsat_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_lvt__vth0_diff_29=0.13606
+  sky130_fd_pr__pfet_01v8_lvt__keta_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_29=0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 030, W = 0.42, L = 4.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ua_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pclm_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_lvt__kt1_diff_30=-0.19799
+  sky130_fd_pr__pfet_01v8_lvt__b0_diff_30=6.0837e-8
+  sky130_fd_pr__pfet_01v8_lvt__pdits_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_lvt__b1_diff_30=1.8757e-7
+  sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_lvt__agidl_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_30=0.063904
+  sky130_fd_pr__pfet_01v8_lvt__ub_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_lvt__k2_diff_30=0.045861
+  sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_lvt__voff_diff_30=-0.0051189
+  sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_lvt__eta0_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ags_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_lvt__a0_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_lvt__u0_diff_30=-0.00025436
+  sky130_fd_pr__pfet_01v8_lvt__vsat_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_lvt__vth0_diff_30=0.10358
+  sky130_fd_pr__pfet_01v8_lvt__keta_diff_30=0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 031, W = 0.42, L = 8.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_lvt__keta_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ua_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pclm_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_lvt__kt1_diff_31=-0.29664
+  sky130_fd_pr__pfet_01v8_lvt__b0_diff_31=1.0853e-7
+  sky130_fd_pr__pfet_01v8_lvt__pdits_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_lvt__b1_diff_31=1.6602e-8
+  sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_lvt__agidl_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_31=0.022441
+  sky130_fd_pr__pfet_01v8_lvt__ub_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_lvt__k2_diff_31=0.04913
+  sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_lvt__voff_diff_31=-0.01143
+  sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_lvt__eta0_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ags_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_lvt__a0_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_lvt__u0_diff_31=-0.00032262
+  sky130_fd_pr__pfet_01v8_lvt__vsat_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_lvt__vth0_diff_31=0.1471
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 032, W = 0.42, L = 0.35
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_lvt__u0_diff_32=-0.00080392
+  sky130_fd_pr__pfet_01v8_lvt__vsat_diff_32=73141.0
+  sky130_fd_pr__pfet_01v8_lvt__vth0_diff_32=0.29494
+  sky130_fd_pr__pfet_01v8_lvt__keta_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ua_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pclm_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_lvt__kt1_diff_32=-1.12
+  sky130_fd_pr__pfet_01v8_lvt__b0_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pdits_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_lvt__b1_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_lvt__agidl_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_32=8.0
+  sky130_fd_pr__pfet_01v8_lvt__ub_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_lvt__k2_diff_32=0.11361
+  sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_lvt__voff_diff_32=-0.45
+  sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_lvt__eta0_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_32=0.006
+  sky130_fd_pr__pfet_01v8_lvt__ags_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_lvt__a0_diff_32=0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 033, W = 0.42, L = 0.5
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_lvt__eta0_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ags_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_lvt__a0_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_lvt__u0_diff_33=-0.00040451
+  sky130_fd_pr__pfet_01v8_lvt__vsat_diff_33=-26432.0
+  sky130_fd_pr__pfet_01v8_lvt__vth0_diff_33=0.14117
+  sky130_fd_pr__pfet_01v8_lvt__keta_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ua_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pclm_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_lvt__kt1_diff_33=-0.593
+  sky130_fd_pr__pfet_01v8_lvt__b0_diff_33=1.4751e-7
+  sky130_fd_pr__pfet_01v8_lvt__pdits_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_lvt__b1_diff_33=2.0999e-7
+  sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_lvt__agidl_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_33=-0.38541
+  sky130_fd_pr__pfet_01v8_lvt__ub_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_lvt__k2_diff_33=0.049869
+  sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_lvt__voff_diff_33=0.05919
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 034, W = 0.55, L = 1.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_lvt__voff_diff_34=0.052219
+  sky130_fd_pr__pfet_01v8_lvt__k2_diff_34=0.074745
+  sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_lvt__eta0_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ags_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_lvt__a0_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_lvt__u0_diff_34=-0.00027176
+  sky130_fd_pr__pfet_01v8_lvt__vsat_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_lvt__vth0_diff_34=0.15751
+  sky130_fd_pr__pfet_01v8_lvt__keta_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ua_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pclm_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_lvt__kt1_diff_34=-0.24322
+  sky130_fd_pr__pfet_01v8_lvt__b0_diff_34=2.8632e-7
+  sky130_fd_pr__pfet_01v8_lvt__pdits_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_lvt__b1_diff_34=3.5539e-7
+  sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_lvt__agidl_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_34=-0.022927
+  sky130_fd_pr__pfet_01v8_lvt__ub_diff_34=0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 035, W = 0.55, L = 2.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_lvt__agidl_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_35=-0.03773
+  sky130_fd_pr__pfet_01v8_lvt__ub_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_lvt__voff_diff_35=0.033552
+  sky130_fd_pr__pfet_01v8_lvt__k2_diff_35=0.064877
+  sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_lvt__eta0_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ags_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_lvt__a0_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_lvt__u0_diff_35=-0.00019897
+  sky130_fd_pr__pfet_01v8_lvt__vsat_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_lvt__vth0_diff_35=0.13136
+  sky130_fd_pr__pfet_01v8_lvt__keta_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ua_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pclm_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_lvt__kt1_diff_35=-0.17416
+  sky130_fd_pr__pfet_01v8_lvt__b0_diff_35=1.9722e-7
+  sky130_fd_pr__pfet_01v8_lvt__pdits_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_lvt__b1_diff_35=2.3556e-7
+  sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_35=0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 036, W = 0.55, L = 4.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_lvt__agidl_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_36=0.027543
+  sky130_fd_pr__pfet_01v8_lvt__ub_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_lvt__voff_diff_36=0.014621
+  sky130_fd_pr__pfet_01v8_lvt__k2_diff_36=0.069899
+  sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_lvt__eta0_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ags_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_lvt__a0_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_lvt__u0_diff_36=-0.00022057
+  sky130_fd_pr__pfet_01v8_lvt__vsat_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_lvt__vth0_diff_36=0.12913
+  sky130_fd_pr__pfet_01v8_lvt__keta_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ua_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pclm_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_lvt__kt1_diff_36=-0.23093
+  sky130_fd_pr__pfet_01v8_lvt__b0_diff_36=2.4068e-7
+  sky130_fd_pr__pfet_01v8_lvt__pdits_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_lvt__b1_diff_36=2.4974e-7
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 037, W = 0.55, L = 8.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_lvt__pdits_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_lvt__b1_diff_37=1.6808e-7
+  sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_lvt__agidl_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_37=0.058378
+  sky130_fd_pr__pfet_01v8_lvt__ub_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_lvt__voff_diff_37=-0.063832
+  sky130_fd_pr__pfet_01v8_lvt__k2_diff_37=0.051472
+  sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_lvt__eta0_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ags_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_lvt__a0_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_lvt__u0_diff_37=-0.00025453
+  sky130_fd_pr__pfet_01v8_lvt__vsat_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_lvt__vth0_diff_37=0.10671
+  sky130_fd_pr__pfet_01v8_lvt__keta_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ua_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pclm_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_lvt__kt1_diff_37=-0.28348
+  sky130_fd_pr__pfet_01v8_lvt__b0_diff_37=1.6138e-7
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 038, W = 0.55, L = 0.35
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_lvt__kt1_diff_38=-0.67185
+  sky130_fd_pr__pfet_01v8_lvt__b0_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pdits_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_lvt__b1_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_lvt__agidl_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ub_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_38=8.0
+  sky130_fd_pr__pfet_01v8_lvt__voff_diff_38=-0.45
+  sky130_fd_pr__pfet_01v8_lvt__k2_diff_38=0.10349
+  sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_lvt__eta0_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ags_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_lvt__a0_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_lvt__u0_diff_38=-0.00081189
+  sky130_fd_pr__pfet_01v8_lvt__vsat_diff_38=43431.0
+  sky130_fd_pr__pfet_01v8_lvt__vth0_diff_38=0.17921
+  sky130_fd_pr__pfet_01v8_lvt__keta_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ua_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_lvt__pclm_diff_38=0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 039, W = 0.55, L = 0.5
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_lvt__pclm_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_lvt__kt1_diff_39=-0.67864
+  sky130_fd_pr__pfet_01v8_lvt__b0_diff_39=2.3872e-7
+  sky130_fd_pr__pfet_01v8_lvt__pdits_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_lvt__b1_diff_39=3.8314e-7
+  sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_lvt__agidl_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ub_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_39=-0.15511
+  sky130_fd_pr__pfet_01v8_lvt__voff_diff_39=0.051343
+  sky130_fd_pr__pfet_01v8_lvt__k2_diff_39=0.045998
+  sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_lvt__eta0_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ags_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_lvt__a0_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_lvt__u0_diff_39=-0.0001216
+  sky130_fd_pr__pfet_01v8_lvt__vsat_diff_39=-28361.0
+  sky130_fd_pr__pfet_01v8_lvt__vth0_diff_39=0.081136
+  sky130_fd_pr__pfet_01v8_lvt__keta_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_lvt__ua_diff_39=0.0
.include "sky130_fd_pr__pfet_01v8_lvt.pm3.spice"
