* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 18
.param
+  sky130_fd_pr__rf_nfet_01v8_b__toxe_mult=1.052
+  sky130_fd_pr__rf_nfet_01v8_b__rbpb_mult=1.2
+  sky130_fd_pr__rf_nfet_01v8_b__overlap_mult=0.9600
+  sky130_fd_pr__rf_nfet_01v8_b__ajunction_mult=1.2169
+  sky130_fd_pr__rf_nfet_01v8_b__pjunction_mult=1.2474
+  sky130_fd_pr__rf_nfet_01v8_b__lint_diff=-1.7325e-8
+  sky130_fd_pr__rf_nfet_01v8_b__wint_diff=3.2175e-8
+  sky130_fd_pr__rf_nfet_01v8_b__rshg_diff=7.0
+  sky130_fd_pr__rf_nfet_01v8_b__dlc_diff=-17.422e-9
+  sky130_fd_pr__rf_nfet_01v8_b__dwc_diff=0.0
+  sky130_fd_pr__rf_nfet_01v8_b__xgw_diff=6.4250e-8
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 000, W = 1.65, L = 0.15
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_bM02__ags_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__vth0_diff_0=0.032714
+  sky130_fd_pr__rf_nfet_01v8_bM02__vsat_diff_0=20474.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__a0_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__b0_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__k2_diff_0=0.0083532
+  sky130_fd_pr__rf_nfet_01v8_bM02__nfactor_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__u0_diff_0=0.00017601
+  sky130_fd_pr__rf_nfet_01v8_bM02__rdsw_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__ua_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__voff_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__b1_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__kt1_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__ub_diff_0=0.0
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 001, W = 1.65, L = 0.18
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_bM02__ags_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__vth0_diff_1=0.032194
+  sky130_fd_pr__rf_nfet_01v8_bM02__vsat_diff_1=21175.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__a0_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__b0_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__k2_diff_1=0.014272
+  sky130_fd_pr__rf_nfet_01v8_bM02__nfactor_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__u0_diff_1=-0.00050746
+  sky130_fd_pr__rf_nfet_01v8_bM02__rdsw_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__ua_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__voff_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__b1_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__kt1_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__ub_diff_1=0.0
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 002, W = 1.65, L = 0.25
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_bM02__kt1_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__ub_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__ags_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__vth0_diff_2=0.018697
+  sky130_fd_pr__rf_nfet_01v8_bM02__vsat_diff_2=32392.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__a0_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__b0_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__k2_diff_2=0.031744
+  sky130_fd_pr__rf_nfet_01v8_bM02__nfactor_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__u0_diff_2=-0.0018379
+  sky130_fd_pr__rf_nfet_01v8_bM02__rdsw_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__ua_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__voff_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__b1_diff_2=0.0
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 003, W = 3.01, L = 0.15
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_bM02__kt1_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__ub_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__ags_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__vth0_diff_3=0.036104
+  sky130_fd_pr__rf_nfet_01v8_bM02__vsat_diff_3=12645.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__a0_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__b0_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__k2_diff_3=0.0022323
+  sky130_fd_pr__rf_nfet_01v8_bM02__nfactor_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__u0_diff_3=-0.0069942
+  sky130_fd_pr__rf_nfet_01v8_bM02__rdsw_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__ua_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__voff_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__b1_diff_3=0.0
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 004, W = 3.01, L = 0.18
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_bM02__voff_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__b1_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__rdsw_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__kt1_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__ub_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__ags_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__vth0_diff_4=0.0098858
+  sky130_fd_pr__rf_nfet_01v8_bM02__vsat_diff_4=23380.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__a0_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__b0_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__k2_diff_4=0.0131
+  sky130_fd_pr__rf_nfet_01v8_bM02__nfactor_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__u0_diff_4=-0.0040868
+  sky130_fd_pr__rf_nfet_01v8_bM02__ua_diff_4=0.0
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 005, W = 3.01, L = 0.25
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_bM02__nfactor_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__ua_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__voff_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__b1_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__rdsw_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__kt1_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__ub_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__ags_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__vth0_diff_5=0.0085637
+  sky130_fd_pr__rf_nfet_01v8_bM02__vsat_diff_5=21055.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__a0_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__b0_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__k2_diff_5=0.032731
+  sky130_fd_pr__rf_nfet_01v8_bM02__u0_diff_5=-0.0019994
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 006, W = 5.05, L = 0.15
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_bM02__u0_diff_6=-0.0048122
+  sky130_fd_pr__rf_nfet_01v8_bM02__nfactor_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__ua_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__voff_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__b1_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__rdsw_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__kt1_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__ub_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__ags_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__vth0_diff_6=0.015103
+  sky130_fd_pr__rf_nfet_01v8_bM02__vsat_diff_6=4095.2
+  sky130_fd_pr__rf_nfet_01v8_bM02__a0_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__b0_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__k2_diff_6=0.0010067
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 007, W = 5.05, L = 0.18
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_bM02__b0_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__k2_diff_7=0.011492
+  sky130_fd_pr__rf_nfet_01v8_bM02__u0_diff_7=-0.0042353
+  sky130_fd_pr__rf_nfet_01v8_bM02__nfactor_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__ua_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__b1_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__rdsw_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__voff_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__kt1_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__ub_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__ags_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__vth0_diff_7=0.0051454
+  sky130_fd_pr__rf_nfet_01v8_bM02__vsat_diff_7=18771.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__a0_diff_7=0.0
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 008, W = 5.05, L = 0.25
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_bM02__a0_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__b0_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__k2_diff_8=0.030405
+  sky130_fd_pr__rf_nfet_01v8_bM02__u0_diff_8=-0.0042395
+  sky130_fd_pr__rf_nfet_01v8_bM02__nfactor_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__ua_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__b1_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__rdsw_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__voff_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__kt1_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__ub_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__ags_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__vth0_diff_8=0.0015836
+  sky130_fd_pr__rf_nfet_01v8_bM02__vsat_diff_8=20830.0
*
* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 000, W = 1.65, L = 0.15
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_bM04__rdsw_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__ua_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__k2_diff_0=0.0072696
+  sky130_fd_pr__rf_nfet_01v8_bM04__u0_diff_0=-0.0014397
+  sky130_fd_pr__rf_nfet_01v8_bM04__vth0_diff_0=0.057292
+  sky130_fd_pr__rf_nfet_01v8_bM04__voff_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__b1_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__kt1_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__nfactor_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__ub_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__vsat_diff_0=10629.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__ags_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__a0_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__b0_diff_0=0.0
*
* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 001, W = 1.65, L = 0.18
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_bM04__b0_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__rdsw_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__ua_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__k2_diff_1=0.018201
+  sky130_fd_pr__rf_nfet_01v8_bM04__u0_diff_1=-0.0021915
+  sky130_fd_pr__rf_nfet_01v8_bM04__vth0_diff_1=0.020199
+  sky130_fd_pr__rf_nfet_01v8_bM04__voff_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__b1_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__kt1_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__nfactor_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__ub_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__vsat_diff_1=24240.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__ags_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__a0_diff_1=0.0
*
* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 002, W = 1.65, L = 0.25
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_bM04__ags_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__a0_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__b0_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__ua_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__rdsw_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__k2_diff_2=0.033909
+  sky130_fd_pr__rf_nfet_01v8_bM04__u0_diff_2=-0.0024784
+  sky130_fd_pr__rf_nfet_01v8_bM04__vth0_diff_2=0.01762
+  sky130_fd_pr__rf_nfet_01v8_bM04__voff_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__b1_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__kt1_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__nfactor_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__ub_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__vsat_diff_2=39930.0
*
* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 003, W = 3.01, L = 0.15
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_bM04__vsat_diff_3=11859.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__ags_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__a0_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__b0_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__ua_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__rdsw_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__k2_diff_3=0.0020408
+  sky130_fd_pr__rf_nfet_01v8_bM04__u0_diff_3=-0.0072915
+  sky130_fd_pr__rf_nfet_01v8_bM04__vth0_diff_3=0.030316
+  sky130_fd_pr__rf_nfet_01v8_bM04__voff_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__b1_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__kt1_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__nfactor_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__ub_diff_3=0.0
*
* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 004, W = 3.01, L = 0.18
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_bM04__kt1_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__nfactor_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__ub_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__vsat_diff_4=27029.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__ags_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__a0_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__b0_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__ua_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__rdsw_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__k2_diff_4=0.015422
+  sky130_fd_pr__rf_nfet_01v8_bM04__u0_diff_4=-0.0070125
+  sky130_fd_pr__rf_nfet_01v8_bM04__vth0_diff_4=0.0054988
+  sky130_fd_pr__rf_nfet_01v8_bM04__voff_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__b1_diff_4=0.0
*
* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 005, W = 3.01, L = 0.25
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_bM04__voff_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__kt1_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__nfactor_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__ub_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__vsat_diff_5=55116.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__ags_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__a0_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__b0_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__ua_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__rdsw_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__k2_diff_5=0.034152
+  sky130_fd_pr__rf_nfet_01v8_bM04__u0_diff_5=-0.0062872
+  sky130_fd_pr__rf_nfet_01v8_bM04__vth0_diff_5=0.0021981
+  sky130_fd_pr__rf_nfet_01v8_bM04__b1_diff_5=0.0
*
* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 006, W = 5.05, L = 0.15
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_bM04__b1_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__voff_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__kt1_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__nfactor_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__ub_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__vsat_diff_6=4091.9
+  sky130_fd_pr__rf_nfet_01v8_bM04__ags_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__a0_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__b0_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__ua_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__rdsw_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__k2_diff_6=0.0010631
+  sky130_fd_pr__rf_nfet_01v8_bM04__u0_diff_6=-0.0047075
+  sky130_fd_pr__rf_nfet_01v8_bM04__vth0_diff_6=0.015982
*
* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 007, W = 5.05, L = 0.18
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_bM04__u0_diff_7=-0.0056998
+  sky130_fd_pr__rf_nfet_01v8_bM04__b1_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__voff_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__kt1_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__ub_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__nfactor_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__vsat_diff_7=12177.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__ags_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__a0_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__b0_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__ua_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__rdsw_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__k2_diff_7=0.014379
+  sky130_fd_pr__rf_nfet_01v8_bM04__vth0_diff_7=-0.0040004
*
* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 008, W = 5.05, L = 0.25
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_bM04__vth0_diff_8=-0.0017169
+  sky130_fd_pr__rf_nfet_01v8_bM04__u0_diff_8=-0.0057354
+  sky130_fd_pr__rf_nfet_01v8_bM04__b1_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__voff_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__kt1_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__ub_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__nfactor_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__vsat_diff_8=47784.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__ags_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__a0_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__b0_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__ua_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__rdsw_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__k2_diff_8=0.03191
.include "sky130_fd_pr__rf_nfet_01v8_b.pm3.spice"
