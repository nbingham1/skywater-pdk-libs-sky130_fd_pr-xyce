* Transistor Vth and I-V characteristic

* Include SkyWater sky130 device models
.include "../sky130_fd_pr__rf_pfet_01v8_hcM04W3p00L0p15.spice"
.lib "../../../models/sky130.lib.spice" tt

* Gate bias
Rg 1 2 680
X1 3 2 5 5 sky130_fd_pr__rf_pfet_01v8_hcM04W3p00L0p15
Rd 3 4 100

* DC source for current measure
Vid 4 0 DC 0V
Vgb 5 1 DC 0V
Vdd 5 0 DC 3.3V

.control
* Sweep Vds from 0 to 1.8V
dc Vdd 0 1.8 0.01 Vgb 0 1.2 0.01
let vgs=V(5) - V ( 1 )
let vds=V(5) - V ( 3 )
wrdata sky130_fd_pr__rf_pfet_01v8_hcM04W3p00L0p15__iv.data Vid#branch vgs vds

* Sweep Vgs from 0 to 1.2V
dc Vgb 0 1.2 0.01
+ # Find threshold
let ih=Vid#branch[98]
let il=Vid#branch[85]
let vh=V(5)[98] - V ( 2 ) [98]
let vl=V(5)[98] - V ( 2 ) [85]
let vth=((vl - vh ) / ( ih - il ) ) * ih vh
echo threshold voltage
print vth
quit
.endc
.end
