* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre=0.0
* statistics {
*   process {
*   }
*   mismatch {
*     vary sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre dist=gauss std = 1.0
*   }
* }
.subckt sky130_fd_pr__pfet_01v8_lvt d g s b
.param l=1 w=1 ad=0 as=0 pd=0 ps=0 nrd=0 nrs=0 sa=0 sb=0 sd=0 mult=1 nf=1.0
msky130_fd_pr__pfet_01v8_lvt d g s b sky130_fd_pr__pfet_01v8_lvt__model l={l} w={w} ad={ad} as={as} pd={pd} ps={ps} nrd={nrd} nrs={nrs} sa={sa} sb={sb} sd={sd} nf={nf}
.model sky130_fd_pr__pfet_01v8_lvt__model.0 pmos
* DC IV MOS Parameters
+  lmin=2.0e-05 lmax=1.0e-04 wmin=7e-06 wmax=1.0e-4
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.4525e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=3.9651e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-7.916e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.44996e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.44996e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.58924+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}
+  k1=0.64774
+  k2=-0.087544
+  k3=3.39
+  dvt0=2.4422
+  dvt1=0.16136
+  dvt2=0.026237
+  dvt0w=0.5
+  dvt1w=1928100.0
+  dvt2w=-0.032
+  w0=1.0e-8
+  k3b=1.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=123760.0
+  ua=-3.0054e-9
+  ub=3.0419e-18
+  uc=4.9353e-11
+  rdsw=484.7
+  prwb=0.1
+  prwg=0.052
+  wr=1.0
+  u0=0.00283229
+  a0=1.74243
+  keta=-0.01258
+  a1=0.0
+  a2=0.46703705
+  ags=0.49444
+  b0=0.0
+  b1=2.1073e-24
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-6.393105e-11
+  cdsc=2.8125e-7
+  cdscb=1.0e-4
+  cdscd=1.0e-10
+  eta0=0.2
+  etab=-0.00025
+  dsub=1.0
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.030097
+  pdiblc1=0.0
+  pdiblc2=0.0018466
+  pdiblcb=-0.025
+  drout=0.43496
+  pscbe1=800000000.0
+  pscbe2=8.6797e-9
+  pvag=0.0
+  delta=0.01363
+  alpha0=5.0449517e-13
+  alpha1=-4.0583656e-18
+  beta0=6.2016506
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=2300000000.0
+  cgidl=0.5
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.60135
+  kt2=-0.055045
+  at=285600.0
+  ute=-0.22271
+  ua1=6.8217e-10
+  ub1=-1.4864e-19
+  uc1=-9.961e-12
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+41
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=1.4472e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=1.0e-11
+  cgso=1.0e-11
+  cgbo=1.0e-13
+  capmod=2.0
+  xpart=0.0
+  cgsl=0.0
+  cgdl=0.0
+  cf=0.0
+  clc=7.0e-8
+  cle=0.492
+  dlc=-5.9781e-8
+  dwc=3.2175e-8
+  vfbcv=-1.0
+  acde=0.44
+  moin=8.7
+  noff=2.6123
+  voffcv=0.112
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000838062107
+  mjs=0.3362
+  pbs=0.6587
+  cjsws=9.9839168e-11
+  mjsws=0.2659
+  pbsws=0.7418
+  cjswgs=2.60659646e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.1 pmos
* DC IV MOS Parameters
+  lmin=8e-06 lmax=2.0e-05 wmin=7e-06 wmax=1.0e-4
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.4525e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=3.9651e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-7.916e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.44996e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.44996e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-0.58924+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}
+  k1=0.64774
+  k2=-0.087544
+  k3=3.39
+  dvt0=2.4422
+  dvt1=0.16136
+  dvt2=0.026237
+  dvt0w=0.5
+  dvt1w=1928100.0
+  dvt2w=-0.032
+  w0=1.0e-8
+  k3b=1.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=123760.0
+  ua=-3.0054e-9
+  ub=3.0419e-18
+  uc=4.9353e-11
+  rdsw=484.7
+  prwb=0.1
+  prwg=0.052
+  wr=1.0
+  u0=0.00283229
+  a0=1.74243
+  keta=-0.01258
+  a1=0.0
+  a2=0.46703705
+  ags=0.49444
+  b0=0.0
+  b1=2.1073e-24
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-6.393105e-11
+  cdsc=2.8125e-7
+  cdscb=1.0e-4
+  cdscd=1.0e-10
+  eta0=0.2
+  etab=-0.00025
+  dsub=1.0
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.030097
+  pdiblc1=0.0
+  pdiblc2=0.0018466
+  pdiblcb=-0.025
+  drout=0.43496
+  pscbe1=800000000.0
+  pscbe2=8.6797e-9
+  pvag=0.0
+  delta=0.01363
+  alpha0=5.0449517e-13
+  alpha1=-4.0583656e-18
+  beta0=6.2016506
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=2300000000.0
+  cgidl=0.5
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.60135
+  kt2=-0.055045
+  at=285600.0
+  ute=-0.22271
+  ua1=6.8217e-10
+  ub1=-1.4864e-19
+  uc1=-9.961e-12
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+41
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=1.4472e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=1.0e-11
+  cgso=1.0e-11
+  cgbo=1.0e-13
+  capmod=2.0
+  xpart=0.0
+  cgsl=0.0
+  cgdl=0.0
+  cf=0.0
+  clc=7.0e-8
+  cle=0.492
+  dlc=-5.9781e-8
+  dwc=3.2175e-8
+  vfbcv=-1.0
+  acde=0.44
+  moin=8.7
+  noff=2.6123
+  voffcv=0.112
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000838062107
+  mjs=0.3362
+  pbs=0.6587
+  cjsws=9.9839168e-11
+  mjsws=0.2659
+  pbsws=0.7418
+  cjswgs=2.60659646e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.2 pmos
* DC IV MOS Parameters
+  lmin=4e-06 lmax=8e-06 wmin=7e-06 wmax=1.0e-4
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.4525e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=3.9651e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-7.916e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.44996e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.44996e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-6.022739767e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0=1.046504510e-7
+  k1=0.64774
+  k2=-8.706152126e-02 lk2=-3.873845907e-9
+  k3=3.39
+  dvt0=2.4422
+  dvt1=0.16136
+  dvt2=0.026237
+  dvt0w=0.5
+  dvt1w=1928100.0
+  dvt2w=-0.032
+  w0=1.0e-8
+  k3b=1.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=123760.0
+  ua=-3.064727761e-09 lua=4.763455615e-16
+  ub=3.131747815e-18 lub=-7.213925990e-25
+  uc=3.769192204e-11 luc=9.362737801e-17
+  rdsw=484.7
+  prwb=0.1
+  prwg=0.052
+  wr=1.0
+  u0=2.744013514e-03 lu0=7.087763159e-10
+  a0=1.827301938e+00 la0=-6.814410358e-7
+  keta=-0.01258
+  a1=0.0
+  a2=0.46703705
+  ags=4.754732471e-01 lags=1.522850072e-7
+  b0=0.0
+  b1=2.1073e-24
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-6.393105e-11
+  cdsc=2.8125e-7
+  cdscb=1.0e-4
+  cdscd=1.0e-10
+  eta0=0.2
+  etab=-0.00025
+  dsub=1.0
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.030097
+  pdiblc1=0.0
+  pdiblc2=5.951487250e-05 lpdiblc2=1.434859584e-8
+  pdiblcb=-0.025
+  drout=0.43496
+  pscbe1=800000000.0
+  pscbe2=8.6797e-9
+  pvag=0.0
+  delta=5.792490487e-03 ldelta=6.292775575e-8
+  alpha0=5.0449517e-13
+  alpha1=-4.0583656e-18
+  beta0=6.2016506
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=2300000000.0
+  cgidl=0.5
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-6.114226250e-01 lkt1=8.087360976e-8
+  kt2=-0.055045
+  at=2.992886974e+05 lat=-1.099072357e-1
+  ute=-3.130916641e-01 lute=7.256789003e-07 wute=4.235164736e-22
+  ua1=6.681489060e-10 lua1=1.125760648e-16
+  ub1=-1.755943445e-19 lub1=2.164177797e-25
+  uc1=-9.961e-12
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+41
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=1.4472e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=1.0e-11
+  cgso=1.0e-11
+  cgbo=1.0e-13
+  capmod=2.0
+  xpart=0.0
+  cgsl=0.0
+  cgdl=0.0
+  cf=0.0
+  clc=7.0e-8
+  cle=0.492
+  dlc=-5.9781e-8
+  dwc=3.2175e-8
+  vfbcv=-1.0
+  acde=0.44
+  moin=8.7
+  noff=2.6123
+  voffcv=0.112
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000838062107
+  mjs=0.3362
+  pbs=0.6587
+  cjsws=9.9839168e-11
+  mjsws=0.2659
+  pbsws=0.7418
+  cjswgs=2.60659646e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.3 pmos
* DC IV MOS Parameters
+  lmin=2e-06 lmax=4e-06 wmin=7e-06 wmax=1.0e-4
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.4525e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=3.9651e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-7.916e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.44996e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.44996e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-5.654750182e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0=-4.361439272e-8
+  k1=0.64774
+  k2=-5.867482080e-02 lk2=-1.182452814e-7
+  k3=3.39
+  dvt0=2.4422
+  dvt1=0.16136
+  dvt2=0.026237
+  dvt0w=0.5
+  dvt1w=1928100.0
+  dvt2w=-0.032
+  w0=1.0e-8
+  k3b=1.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=1.572514993e+05 lvsat=-1.349389253e-1
+  ua=-3.116027127e-09 lua=6.830332731e-16
+  ub=3.179750695e-18 lub=-9.147986027e-25
+  uc=7.050407242e-11 luc=-3.857441650e-17
+  rdsw=484.7
+  prwb=0.1
+  prwg=0.052
+  wr=1.0
+  u0=2.640966061e-03 lu0=1.123959659e-9
+  a0=2.325843537e+00 la0=-2.690090064e-6
+  keta=-0.01258
+  a1=0.0
+  a2=0.46703705
+  ags=4.838792107e-01 lags=1.184169594e-7
+  b0=0.0
+  b1=2.1073e-24
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-6.393105e-11
+  cdsc=2.8125e-7
+  cdscb=1.0e-4
+  cdscd=1.0e-10
+  eta0=0.2
+  etab=-0.00025
+  dsub=1.0
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.030097
+  pdiblc1=0.0
+  pdiblc2=2.055030400e-04 lpdiblc2=1.376040222e-8
+  pdiblcb=-0.025
+  drout=0.43496
+  pscbe1=800000000.0
+  pscbe2=8.6797e-9
+  pvag=0.0
+  delta=1.964978460e-02 ldelta=7.096024907e-9
+  alpha0=5.0449517e-13
+  alpha1=-4.0583656e-18
+  beta0=6.2016506
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=2300000000.0
+  cgidl=0.5
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.59135
+  kt2=-0.055045
+  at=3.798742980e+05 lat=-4.345906499e-1
+  ute=-0.13298
+  ua1=6.9609e-10
+  ub1=-1.577383861e-19 lub1=1.444752306e-25
+  uc1=-9.961e-12
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+41
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=1.4472e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=1.0e-11
+  cgso=1.0e-11
+  cgbo=1.0e-13
+  capmod=2.0
+  xpart=0.0
+  cgsl=0.0
+  cgdl=0.0
+  cf=0.0
+  clc=7.0e-8
+  cle=0.492
+  dlc=-5.9781e-8
+  dwc=3.2175e-8
+  vfbcv=-1.0
+  acde=0.44
+  moin=8.7
+  noff=2.6123
+  voffcv=0.112
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000838062107
+  mjs=0.3362
+  pbs=0.6587
+  cjsws=9.9839168e-11
+  mjsws=0.2659
+  pbsws=0.7418
+  cjswgs=2.60659646e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.4 pmos
* DC IV MOS Parameters
+  lmin=1.5e-06 lmax=2e-06 wmin=7e-06 wmax=1.0e-4
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.4525e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=3.9651e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-7.916e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.44996e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.44996e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-5.958690710e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0=1.805666001e-8
+  k1=0.64774
+  k2=-1.861894421e-01 lk2=1.404882609e-7
+  k3=3.39
+  dvt0=2.4422
+  dvt1=0.16136
+  dvt2=0.026237
+  dvt0w=0.5
+  dvt1w=1928100.0
+  dvt2w=-0.032
+  w0=1.0e-8
+  k3b=1.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=90748.0
+  ua=-2.222214180e-09 lua=-1.130557888e-15
+  ub=1.811164190e-18 lub=1.862131845e-24
+  uc=-9.800498300e-12 luc=1.243675727e-16
+  rdsw=484.7
+  prwb=0.1
+  prwg=0.052
+  wr=1.0
+  u0=3.397162734e-03 lu0=-4.104012004e-10
+  a0=1.275301624e+00 la0=-5.584879955e-7
+  keta=-0.01258
+  a1=0.0
+  a2=0.46703705
+  ags=2.616899060e-01 lags=5.692501682e-7
+  b0=0.0
+  b1=2.1073e-24
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-6.393105e-11
+  cdsc=2.8125e-7
+  cdscb=1.0e-4
+  cdscd=1.0e-10
+  eta0=0.2
+  etab=-0.00025
+  dsub=1.0
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.030097
+  pdiblc1=0.0
+  pdiblc2=-3.516761880e-03 lpdiblc2=2.131306385e-8
+  pdiblcb=-0.025
+  drout=0.43496
+  pscbe1=800000000.0
+  pscbe2=8.6797e-9
+  pvag=0.0
+  delta=1.682590730e-02 ldelta=1.282581314e-8
+  alpha0=5.0449517e-13
+  alpha1=-4.0583656e-18
+  beta0=6.2016506
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=2300000000.0
+  cgidl=0.5
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.59135
+  kt2=-0.055045
+  at=2.067602830e+05 lat=-8.333365772e-2
+  ute=-0.13298
+  ua1=8.025118800e-10 lua1=-2.159353156e-16
+  ub1=-3.177120695e-19 lub1=4.690698329e-25
+  uc1=-9.961e-12
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+41
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=1.4472e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=1.0e-11
+  cgso=1.0e-11
+  cgbo=1.0e-13
+  capmod=2.0
+  xpart=0.0
+  cgsl=0.0
+  cgdl=0.0
+  cf=0.0
+  clc=7.0e-8
+  cle=0.492
+  dlc=-5.9781e-8
+  dwc=3.2175e-8
+  vfbcv=-1.0
+  acde=0.44
+  moin=8.7
+  noff=2.6123
+  voffcv=0.112
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000838062107
+  mjs=0.3362
+  pbs=0.6587
+  cjsws=9.9839168e-11
+  mjsws=0.2659
+  pbsws=0.7418
+  cjswgs=2.60659646e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.5 pmos
* DC IV MOS Parameters
+  lmin=1e-06 lmax=1.5e-06 wmin=7e-06 wmax=1.0e-4
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.4525e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=3.9651e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-7.916e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.44996e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.44996e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-5.762392200e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0=-1.195836366e-8
+  k1=0.64774
+  k2=-5.284545930e-02 lk2=-6.340135596e-8
+  k3=3.39
+  dvt0=2.4422
+  dvt1=0.16136
+  dvt2=0.026237
+  dvt0w=0.5
+  dvt1w=1928100.0
+  dvt2w=-0.032
+  w0=1.0e-8
+  k3b=1.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=9.000090970e+04 lvsat=1.142338423e-3
+  ua=-3.159795030e-09 lua=3.030501106e-16
+  ub=3.144871030e-18 lub=-1.771725984e-25
+  uc=8.781968720e-11 luc=-2.489857191e-17
+  rdsw=484.7
+  prwb=0.1
+  prwg=0.052
+  wr=1.0
+  u0=2.260077152e-03 lu0=1.328259509e-9
+  a0=6.360654375e-01 la0=4.189360953e-7
+  keta=-0.01258
+  a1=0.0
+  a2=0.46703705
+  ags=-1.257058720e-01 lags=1.161597683e-6
+  b0=0.0
+  b1=2.1073e-24
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-1.519546450e-01+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff=-4.578794506e-8
+  nfactor={2.599866240e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-9.566690927e-8
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-6.393105e-11
+  cdsc=2.8125e-7
+  cdscb=1.0e-4
+  cdscd=1.0e-10
+  eta0=0.2
+  etab=-0.00025
+  dsub=1.0
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.030097
+  pdiblc1=0.0
+  pdiblc2=2.549860000e-04 lpdiblc2=1.554587276e-8
+  pdiblcb=-0.025
+  drout=0.43496
+  pscbe1=800000000.0
+  pscbe2=8.6797e-9
+  pvag=0.0
+  delta=9.714448900e-03 ldelta=2.369958861e-8
+  alpha0=5.0449517e-13
+  alpha1=-4.0583656e-18
+  beta0=6.2016506
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=2300000000.0
+  cgidl=0.5
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-6.530930000e-01 lkt1=9.440813415e-8
+  kt2=-9.469635460e-02 lkt2=6.062890375e-8
+  at=2.061616390e+05 lat=-8.241830111e-2
+  ute=6.274531000e-02 lute=-2.992737853e-7
+  ua1=6.6129e-10
+  ub1=-1.048927610e-20 lub1=-6.891793793e-28
+  uc1=-9.961e-12
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+41
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=1.4472e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=1.0e-11
+  cgso=1.0e-11
+  cgbo=1.0e-13
+  capmod=2.0
+  xpart=0.0
+  cgsl=0.0
+  cgdl=0.0
+  cf=0.0
+  clc=7.0e-8
+  cle=0.492
+  dlc=-5.9781e-8
+  dwc=3.2175e-8
+  vfbcv=-1.0
+  acde=0.44
+  moin=8.7
+  noff=2.6123
+  voffcv=0.112
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000838062107
+  mjs=0.3362
+  pbs=0.6587
+  cjsws=9.9839168e-11
+  mjsws=0.2659
+  pbsws=0.7418
+  cjswgs=2.60659646e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=2.74e-6
+  sbref=2.74e-6
+  wlod={0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.6 pmos
* DC IV MOS Parameters
+  lmin=5e-07 lmax=1e-06 wmin=7e-06 wmax=1.0e-4
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.4525e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=3.9651e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-7.916e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.44996e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.44996e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-6.007476580e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0=1.326204446e-8
+  k1=0.64774
+  k2=-1.417083655e-01 lk2=2.804301767e-08 wk2=2.117582368e-22
+  k3=3.39
+  dvt0=2.4422
+  dvt1=0.16136
+  dvt2=0.026237
+  dvt0w=0.5
+  dvt1w=1928100.0
+  dvt2w=-0.032
+  w0=1.0e-8
+  k3b=1.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=1.979082760e+04 lvsat=7.339202341e-2
+  ua=-2.784566970e-09 lua=-8.307832452e-17
+  ub=2.814725670e-18 lub=1.625634843e-25
+  uc=5.745739320e-11 luc=6.345746728e-18
+  rdsw=484.7
+  prwb=0.1
+  prwg=0.052
+  wr=1.0
+  u0=3.601967392e-03 lu0=-5.261264274e-11
+  a0=1.074211189e+00 la0=-3.193779050e-8
+  keta=-0.01258
+  a1=0.0
+  a2=0.46703705
+  ags=1.619157563e+00 lags=-6.339540352e-7
+  b0=2.017161840e-06 lb0=-2.075760391e-12
+  b1=2.1073e-24
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-2.118453550e-01+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff=1.584259006e-8
+  nfactor={2.474733760e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=3.310066927e-8
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-6.393105e-11
+  cdsc=2.8125e-7
+  cdscb=1.0e-4
+  cdscd=1.0e-10
+  eta0=0.2
+  etab=-0.00025
+  dsub=1.0
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.030097
+  pdiblc1=0.0
+  pdiblc2=-2.541823210e-02 lpdiblc2=4.196489784e-8
+  pdiblcb=-0.025
+  drout=0.43496
+  pscbe1=800000000.0
+  pscbe2=8.6797e-9
+  pvag=0.0
+  delta=2.057155950e-02 ldelta=1.252707895e-8
+  alpha0=5.0449517e-13
+  alpha1=-4.0583656e-18
+  beta0=6.2016506
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=2300000000.0
+  cgidl=0.5
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-4.866375590e-01 lkt1=-7.688283741e-8
+  kt2=-1.436728840e-02 lkt2=-2.203372182e-8
+  at=1.966812454e+05 lat=-7.266250208e-2
+  ute=-4.777976000e-02 lute=-1.855379620e-7
+  ua1=4.125730140e-10 lua1=2.559422144e-16
+  ub1=6.110683441e-19 lub1=-6.403030484e-25 wub1=3.443831106e-40 pub1=-1.423193753e-46
+  uc1=-2.375269864e-11 luc1=1.419234749e-17
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+41
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=1.4472e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=1.0e-11
+  cgso=1.0e-11
+  cgbo=1.0e-13
+  capmod=2.0
+  xpart=0.0
+  cgsl=0.0
+  cgdl=0.0
+  cf=0.0
+  clc=7.0e-8
+  cle=0.492
+  dlc=-5.9781e-8
+  dwc=3.2175e-8
+  vfbcv=-1.0
+  acde=0.44
+  moin=8.7
+  noff=2.6123
+  voffcv=0.112
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000838062107
+  mjs=0.3362
+  pbs=0.6587
+  cjsws=9.9839168e-11
+  mjsws=0.2659
+  pbsws=0.7418
+  cjswgs=2.60659646e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.74e-6
+  sbref=1.74e-6
+  wlod={0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.7 pmos
* DC IV MOS Parameters
+  lmin=3.5e-07 lmax=5e-07 wmin=7e-06 wmax=1.0e-4
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.4525e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=3.9651e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-7.916e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.44996e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.44996e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope3/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-5.845497700e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0=4.692551819e-9
+  k1=0.64774
+  k2=-9.621982500e-02 lk2=3.977305316e-9
+  k3=3.39
+  dvt0=2.4422
+  dvt1=0.16136
+  dvt2=0.026237
+  dvt0w=0.5
+  dvt1w=1928100.0
+  dvt2w=-0.032
+  w0=1.0e-8
+  k3b=1.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=2.357679170e+05 lvsat=-4.087065574e-2
+  ua=-3.087407900e-09 lua=7.713966950e-17
+  ub=3.020920000e-18 lub=5.347637400e-26
+  uc=8.540747800e-11 luc=-8.441245636e-18
+  rdsw=484.7
+  prwb=0.1
+  prwg=0.052
+  wr=1.0
+  u0=2.489799480e-03 lu0=5.357797911e-10
+  a0=1.048824261e+00 la0=-1.850683613e-8
+  keta=-0.01258
+  a1=0.0
+  a2=0.46703705
+  ags=4.101302500e-01 lags=5.681864738e-9
+  b0=-6.723872800e-06 lb0=2.548683985e-12
+  b1=2.1073e-24
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-6.393105e-11
+  cdsc=2.8125e-7
+  cdscb=1.0e-4
+  cdscd=1.0e-10
+  eta0=0.2
+  etab=-0.00025
+  dsub=1.0
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.030097
+  pdiblc1=0.0
+  pdiblc2=-1.028139590e-01 lpdiblc2=8.291110716e-8
+  pdiblcb=-0.025
+  drout=0.43496
+  pscbe1=800000000.0
+  pscbe2=8.6797e-9
+  pvag=0.0
+  delta=2.294991700e-02 ldelta=1.126880891e-8
+  alpha0=5.0449517e-13
+  alpha1=-4.0583656e-18
+  beta0=6.2016506
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=2300000000.0
+  cgidl=0.5
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-6.572300000e-01 lkt1=1.336909350e-8
+  kt2=-0.056015
+  at=1.455597670e+05 lat=-4.561668393e-2
+  ute=-0.39848
+  ua1=8.9635e-10
+  ub1=-5.9922e-19
+  uc1=3.0734e-12
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+41
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=1.4472e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=1.0e-11
+  cgso=1.0e-11
+  cgbo=1.0e-13
+  capmod=2.0
+  xpart=0.0
+  cgsl=0.0
+  cgdl=0.0
+  cf=0.0
+  clc=7.0e-8
+  cle=0.492
+  dlc=-5.9781e-8
+  dwc=3.2175e-8
+  vfbcv=-1.0
+  acde=0.44
+  moin=8.7
+  noff=2.6123
+  voffcv=0.112
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000838062107
+  mjs=0.3362
+  pbs=0.6587
+  cjsws=9.9839168e-11
+  mjsws=0.2659
+  pbsws=0.7418
+  cjswgs=2.60659646e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.44e-6
+  sbref=1.44e-6
+  wlod={0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.8 pmos
* DC IV MOS Parameters
+  lmin=2.0e-05 lmax=1.0e-04 wmin=5.0e-06 wmax=7.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.4525e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=3.9651e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-7.916e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.44996e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.44996e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-6.373398229e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0=3.328843485e-7
+  k1=0.64774
+  k2=-9.397781263e-02 wk2=4.452647424e-8
+  k3=3.39
+  dvt0=2.4422
+  dvt1=0.16136
+  dvt2=0.026237
+  dvt0w=0.5
+  dvt1w=1928100.0
+  dvt2w=-0.032
+  w0=1.0e-8
+  k3b=1.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=123760.0
+  ua=-3.120298298e-09 wua=7.951764232e-16
+  ub=3.229624629e-18 wub=-1.299185462e-24
+  uc=5.085135254e-11 wuc=-1.036964543e-17
+  rdsw=484.7
+  prwb=0.1
+  prwg=0.052
+  wr=1.0
+  u0=2.960203545e-03 wu0=-8.852510117e-10
+  a0=1.719794789e+00 wa0=1.566514581e-7
+  keta=-0.01258
+  a1=0.0
+  a2=0.46703705
+  ags=5.828649431e-01 wags=-6.119623266e-7
+  b0=0.0
+  b1=2.1073e-24
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-6.393105e-11
+  cdsc=2.8125e-7
+  cdscb=1.0e-4
+  cdscd=1.0e-10
+  eta0=0.2
+  etab=-0.00025
+  dsub=1.0
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.030097
+  pdiblc1=0.0
+  pdiblc2=2.344328603e-03 wpdiblc2=-3.444629345e-9
+  pdiblcb=-0.025
+  drout=0.43496
+  pscbe1=800000000.0
+  pscbe2=8.6797e-9
+  pvag=0.0
+  delta=3.616379570e-03 wdelta=6.930124288e-8
+  alpha0=5.0449517e-13
+  alpha1=-4.0583656e-18
+  beta0=6.2016506
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=2300000000.0
+  cgidl=0.5
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.60135
+  kt2=-0.055045
+  at=285600.0
+  ute=-0.22271
+  ua1=6.8217e-10
+  ub1=-1.4864e-19
+  uc1=-9.961e-12
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+41
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=1.4472e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=1.0e-11
+  cgso=1.0e-11
+  cgbo=1.0e-13
+  capmod=2.0
+  xpart=0.0
+  cgsl=0.0
+  cgdl=0.0
+  cf=0.0
+  clc=7.0e-8
+  cle=0.492
+  dlc=-5.9781e-8
+  dwc=3.2175e-8
+  vfbcv=-1.0
+  acde=0.44
+  moin=8.7
+  noff=2.6123
+  voffcv=0.112
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000838062107
+  mjs=0.3362
+  pbs=0.6587
+  cjsws=9.9839168e-11
+  mjsws=0.2659
+  pbsws=0.7418
+  cjswgs=2.60659646e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.9 pmos
* DC IV MOS Parameters
+  lmin=8e-06 lmax=2.0e-05 wmin=5.0e-06 wmax=7.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.4525e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=3.9651e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-7.916e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.44996e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.44996e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-6.373398230e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0=3.328843485e-7
+  k1=0.64774
+  k2=-9.397781264e-02 wk2=4.452647424e-8
+  k3=3.39
+  dvt0=2.4422
+  dvt1=0.16136
+  dvt2=0.026237
+  dvt0w=0.5
+  dvt1w=1928100.0
+  dvt2w=-0.032
+  w0=1.0e-8
+  k3b=1.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=123760.0
+  ua=-3.120298298e-09 wua=7.951764232e-16
+  ub=3.229624629e-18 wub=-1.299185462e-24
+  uc=5.085135254e-11 wuc=-1.036964543e-17
+  rdsw=484.7
+  prwb=0.1
+  prwg=0.052
+  wr=1.0
+  u0=2.960203545e-03 wu0=-8.852510117e-10
+  a0=1.719794789e+00 wa0=1.566514581e-7
+  keta=-0.01258
+  a1=0.0
+  a2=0.46703705
+  ags=5.828649431e-01 wags=-6.119623266e-7
+  b0=0.0
+  b1=2.1073e-24
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-6.393105e-11
+  cdsc=2.8125e-7
+  cdscb=1.0e-4
+  cdscd=1.0e-10
+  eta0=0.2
+  etab=-0.00025
+  dsub=1.0
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.030097
+  pdiblc1=0.0
+  pdiblc2=2.344328603e-03 wpdiblc2=-3.444629345e-9
+  pdiblcb=-0.025
+  drout=0.43496
+  pscbe1=800000000.0
+  pscbe2=8.6797e-9
+  pvag=0.0
+  delta=3.616379570e-03 wdelta=6.930124288e-8
+  alpha0=5.0449517e-13
+  alpha1=-4.0583656e-18
+  beta0=6.2016506
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=2300000000.0
+  cgidl=0.5
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.60135
+  kt2=-0.055045
+  at=285600.0
+  ute=-0.22271
+  ua1=6.8217e-10
+  ub1=-1.4864e-19
+  uc1=-9.961e-12
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+41
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=1.4472e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=1.0e-11
+  cgso=1.0e-11
+  cgbo=1.0e-13
+  capmod=2.0
+  xpart=0.0
+  cgsl=0.0
+  cgdl=0.0
+  cf=0.0
+  clc=7.0e-8
+  cle=0.492
+  dlc=-5.9781e-8
+  dwc=3.2175e-8
+  vfbcv=-1.0
+  acde=0.44
+  moin=8.7
+  noff=2.6123
+  voffcv=0.112
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000838062107
+  mjs=0.3362
+  pbs=0.6587
+  cjsws=9.9839168e-11
+  mjsws=0.2659
+  pbsws=0.7418
+  cjswgs=2.60659646e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.10 pmos
* DC IV MOS Parameters
+  lmin=4e-06 lmax=8e-06 wmin=5.0e-06 wmax=7.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.4525e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=3.9651e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-7.916e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.44996e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.44996e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-6.797902389e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0=3.408365119e-07 wvth0=5.364666402e-07 pvth0=-1.634572399e-12
+  k1=0.64774
+  k2=-1.161065884e-01 lk2=1.776730471e-07 wk2=2.010121381e-07 pk2=-1.256431219e-12
+  k3=3.39
+  dvt0=2.4422
+  dvt1=0.16136
+  dvt2=0.026237
+  dvt0w=0.5
+  dvt1w=1928100.0
+  dvt2w=-0.032
+  w0=1.0e-8
+  k3b=1.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=123760.0
+  ua=-3.325593058e-09 lua=1.648321887e-15 wua=1.805369935e-15 pua=-8.110894214e-21
+  ub=3.540529425e-18 lub=-2.496270159e-24 wub=-2.829054074e-24 pub=1.228339158e-29
+  uc=1.049995307e-11 luc=3.239834039e-16 wuc=1.881874052e-16 puc=-1.594224488e-21
+  rdsw=484.7
+  prwb=0.1
+  prwg=0.052
+  wr=1.0
+  u0=2.762811152e-03 lu0=1.584873389e-09 wu0=-1.300927720e-10 pu0=-6.063203264e-15
+  a0=2.026714996e+00 la0=-2.464277688e-06 wa0=-1.380077551e-06 pa0=1.233847405e-11
+  keta=-0.01258
+  a1=0.0
+  a2=0.46703705
+  ags=6.601273673e-01 lags=-6.203438677e-07 wags=-1.277935401e-06 pags=5.347131109e-12
+  b0=0.0
+  b1=2.1073e-24
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-6.393105e-11
+  cdsc=2.8125e-7
+  cdscb=1.0e-4
+  cdscd=1.0e-10
+  eta0=0.2
+  etab=-0.00025
+  dsub=1.0
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.030097
+  pdiblc1=0.0
+  pdiblc2=-1.458267684e-04 lpdiblc2=1.999358198e-08 wpdiblc2=1.421107484e-09 ppdiblc2=-3.906724429e-14
+  pdiblcb=-0.025
+  drout=0.43496
+  pscbe1=800000000.0
+  pscbe2=8.6797e-9
+  pvag=0.0
+  delta=-1.183421344e-02 ldelta=1.240535838e-07 wdelta=1.219890946e-07 pdelta=-4.230333960e-13
+  alpha0=5.0449517e-13
+  alpha1=-4.0583656e-18
+  beta0=6.2016506
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=2300000000.0
+  cgidl=0.5
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-6.114226250e-01 lkt1=8.087360976e-8
+  kt2=-0.055045
+  at=2.992886974e+05 lat=-1.099072357e-1
+  ute=-3.130916641e-01 lute=7.256789003e-7
+  ua1=6.681489060e-10 lua1=1.125760648e-16
+  ub1=-1.755943445e-19 lub1=2.164177797e-25
+  uc1=-9.961e-12
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+41
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=1.4472e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=1.0e-11
+  cgso=1.0e-11
+  cgbo=1.0e-13
+  capmod=2.0
+  xpart=0.0
+  cgsl=0.0
+  cgdl=0.0
+  cf=0.0
+  clc=7.0e-8
+  cle=0.492
+  dlc=-5.9781e-8
+  dwc=3.2175e-8
+  vfbcv=-1.0
+  acde=0.44
+  moin=8.7
+  noff=2.6123
+  voffcv=0.112
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000838062107
+  mjs=0.3362
+  pbs=0.6587
+  cjsws=9.9839168e-11
+  mjsws=0.2659
+  pbsws=0.7418
+  cjswgs=2.60659646e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.11 pmos
* DC IV MOS Parameters
+  lmin=2e-06 lmax=4e-06 wmin=5.0e-06 wmax=7.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.4525e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=3.9651e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-7.916e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.44996e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.44996e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-6.096308845e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0=5.816096533e-08 wvth0=3.055894155e-07 pvth0=-7.043565169e-13
+  k1=0.64774
+  k2=3.042248022e-02 lk2=-4.126998969e-07 wk2=-6.166155130e-07 pk2=2.037831468e-12
+  k3=3.39
+  dvt0=2.4422
+  dvt1=0.16136
+  dvt2=0.026237
+  dvt0w=0.5
+  dvt1w=1928100.0
+  dvt2w=-0.032
+  w0=1.0e-8
+  k3b=1.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=2.396522761e+05 lvsat=-4.669357751e-01 wvsat=-5.702708913e-01 pvsat=2.297649934e-6
+  ua=-3.650875034e-09 lua=2.958899234e-15 wua=3.701520837e-15 pua=-1.575058101e-20
+  ub=4.002671892e-18 lub=-4.358265263e-24 wub=-5.695189081e-24 pub=2.383119283e-29
+  uc=1.422928225e-10 luc=-2.070166568e-16 wuc=-4.968282593e-16 puc=1.165737876e-21
+  rdsw=484.7
+  prwb=0.1
+  prwg=0.052
+  wr=1.0
+  u0=2.552667726e-03 lu0=2.431551760e-09 wu0=6.110861086e-10 pu0=-9.049450033e-15
+  a0=3.633417835e+00 la0=-8.937763762e-06 wa0=-9.049326831e-06 pa0=4.323826286e-11
+  keta=-0.01258
+  a1=0.0
+  a2=0.46703705
+  ags=9.156305669e-01 lags=-1.649779034e-06 wags=-2.988020747e-06 pags=1.223715048e-11
+  b0=0.0
+  b1=2.1073e-24
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-6.393105e-11
+  cdsc=2.8125e-7
+  cdscb=1.0e-4
+  cdscd=1.0e-10
+  eta0=0.2
+  etab=-0.00025
+  dsub=1.0
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.030097
+  pdiblc1=0.0
+  pdiblc2=2.305065239e-03 lpdiblc2=1.011881554e-08 wpdiblc2=-1.453043591e-08 ppdiblc2=2.520232162e-14
+  pdiblcb=-0.025
+  drout=0.43496
+  pscbe1=800000000.0
+  pscbe2=8.6797e-9
+  pvag=0.0
+  delta=3.353622852e-02 ldelta=-5.874619537e-08 wdelta=-9.610388466e-08 pdelta=4.556741222e-13
+  alpha0=5.0449517e-13
+  alpha1=-4.0583656e-18
+  beta0=6.2016506
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=2300000000.0
+  cgidl=0.5
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.59135
+  kt2=-0.055045
+  at=5.841539410e+05 lat=-1.257643545e+00 wat=-1.413757717e+00 pat=5.696100528e-6
+  ute=-0.13298
+  ua1=6.9609e-10
+  ub1=-2.459625306e-19 lub1=4.999347198e-25 wub1=6.105726600e-25 pub1=-2.460027776e-30
+  uc1=-9.961e-12
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+41
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=1.4472e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=1.0e-11
+  cgso=1.0e-11
+  cgbo=1.0e-13
+  capmod=2.0
+  xpart=0.0
+  cgsl=0.0
+  cgdl=0.0
+  cf=0.0
+  clc=7.0e-8
+  cle=0.492
+  dlc=-5.9781e-8
+  dwc=3.2175e-8
+  vfbcv=-1.0
+  acde=0.44
+  moin=8.7
+  noff=2.6123
+  voffcv=0.112
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000838062107
+  mjs=0.3362
+  pbs=0.6587
+  cjsws=9.9839168e-11
+  mjsws=0.2659
+  pbsws=0.7418
+  cjswgs=2.60659646e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.12 pmos
* DC IV MOS Parameters
+  lmin=1.5e-06 lmax=2e-06 wmin=5.0e-06 wmax=7.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.4525e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=3.9651e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-7.916e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.44996e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.44996e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-3.958220328e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0=-3.756678852e-07 wvth0=-1.384465137e-06 pvth0=2.724848673e-12
+  k1=0.64774
+  k2=-3.768684965e-01 lk2=4.137138595e-07 wk2=1.319632150e-06 pk2=-1.890911853e-12
+  k3=3.39
+  dvt0=2.4422
+  dvt1=0.16136
+  dvt2=0.026237
+  dvt0w=0.5
+  dvt1w=1928100.0
+  dvt2w=-0.032
+  w0=1.0e-8
+  k3b=1.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=-3.905839557e+05 lvsat=8.118450510e-01 wvsat=3.331153103e+00 pvsat=-5.618534421e-6
+  ua=-4.737163815e-10 lua=-3.487714530e-15 wua=-1.210082522e-14 pua=1.631316925e-20
+  ub=-8.431746190e-19 lub=5.474199600e-24 wub=1.836987729e-23 pub=-2.499803009e-29
+  uc=-7.410884336e-11 luc=2.320731434e-16 wuc=4.450586350e-16 puc=-7.453977272e-22
+  rdsw=484.7
+  prwb=0.1
+  prwg=0.052
+  wr=1.0
+  u0=3.763996351e-03 lu0=-2.629458709e-11 wu0=-2.538744680e-09 pu0=-2.658285871e-15
+  a0=2.447259018e+00 la0=-6.530988214e-06 wa0=-8.110763195e-06 pa0=4.133387031e-11
+  keta=-0.01258
+  a1=0.0
+  a2=0.46703705
+  ags=2.798359271e-01 lags=-3.597199201e-07 wags=-1.255831320e-07 pags=6.429121432e-12
+  b0=0.0
+  b1=2.1073e-24
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-6.393105e-11
+  cdsc=2.8125e-7
+  cdscb=1.0e-4
+  cdscd=1.0e-10
+  eta0=0.2
+  etab=-0.00025
+  dsub=1.0
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.030097
+  pdiblc1=0.0
+  pdiblc2=-7.034865623e-03 lpdiblc2=2.907000226e-08 wpdiblc2=2.434773354e-08 ppdiblc2=-5.368342810e-14
+  pdiblcb=-0.025
+  drout=0.43496
+  pscbe1=800000000.0
+  pscbe2=8.6797e-9
+  pvag=0.0
+  delta=-6.342109790e-03 ldelta=2.216894698e-08 wdelta=1.603388495e-07 pdelta=-6.466100766e-14
+  alpha0=5.0449517e-13
+  alpha1=-4.0583656e-18
+  beta0=6.2016506
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=2300000000.0
+  cgidl=0.5
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-8.170697983e-01 lkt1=4.579967568e-07 wkt1=1.562138557e-06 pkt1=-3.169657238e-12
+  kt2=-2.082861711e-01 lkt2=3.109339982e-07 wkt2=1.060535866e-06 pkt2=-2.151880299e-12
+  at=-8.509003540e+05 lat=1.654153372e+00 wat=7.319749855e+00 pat=-1.202462301e-5
+  ute=-0.13298
+  ua1=8.493111182e-10 lua1=-3.108933098e-16 wua1=-3.238833941e-16 pua1=6.571756008e-22
+  ub1=3.518450828e-20 lub1=-7.052667938e-26 wub1=-2.442290640e-24 pub1=3.734384503e-30
+  uc1=-9.961e-12
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+41
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=1.4472e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=1.0e-11
+  cgso=1.0e-11
+  cgbo=1.0e-13
+  capmod=2.0
+  xpart=0.0
+  cgsl=0.0
+  cgdl=0.0
+  cf=0.0
+  clc=7.0e-8
+  cle=0.492
+  dlc=-5.9781e-8
+  dwc=3.2175e-8
+  vfbcv=-1.0
+  acde=0.44
+  moin=8.7
+  noff=2.6123
+  voffcv=0.112
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000838062107
+  mjs=0.3362
+  pbs=0.6587
+  cjsws=9.9839168e-11
+  mjsws=0.2659
+  pbsws=0.7418
+  cjswgs=2.60659646e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.13 pmos
* DC IV MOS Parameters
+  lmin=1e-06 lmax=1.5e-06 wmin=5.0e-06 wmax=7.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.4525e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=3.9651e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-7.916e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.44996e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.44996e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-5.591515254e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0=-1.259289246e-07 wvth0=-1.182587739e-07 pvth0=7.887558332e-13
+  k1=0.64774
+  k2=4.328419262e-02 lk2=-2.287206098e-07 wk2=-6.652842898e-07 pk2=1.144124630e-12
+  k3=3.39
+  dvt0=2.4422
+  dvt1=0.16136
+  dvt2=0.026237
+  dvt0w=0.5
+  dvt1w=1928100.0
+  dvt2w=-0.032
+  w0=1.0e-8
+  k3b=1.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=4.301935345e+05 lvsat=-4.431647703e-01 wvsat=-2.354370418e+00 pvsat=3.074915318e-6
+  ua=-3.237962852e-09 lua=7.389565360e-16 wua=5.409758886e-16 pua=-3.016776726e-21
+  ub=3.137910776e-18 lub=-6.130790238e-25 wub=4.816981255e-26 pub=3.016776726e-30
+  uc=1.685889935e-10 luc=-1.390239842e-16 wuc=-5.589799769e-16 puc=7.898275123e-22
+  rdsw=484.7
+  prwb=0.1
+  prwg=0.052
+  wr=1.0
+  u0=2.008992917e-03 lu0=2.657193414e-09 wu0=1.737678162e-09 pu0=-9.197150218e-15
+  a0=-5.608885275e+00 la0=5.787259218e-06 wa0=4.321941791e-05 pa0=-3.715254310e-11
+  keta=-0.01258
+  a1=0.0
+  a2=0.46703705
+  ags=-2.907209322e+00 lags=4.513431619e-06 wags=1.924994537e-05 pags=-2.319703042e-11
+  b0=0.0
+  b1=2.1073e-24
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-7.827862077e-02+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff=-1.584422699e-07 wvoff=-5.098895135e-07 pvoff=7.796465607e-13
+  nfactor={2.753801026e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-3.310408938e-07 wnfactor=-1.065336166e-06 pnfactor=1.628952264e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-6.393105e-11
+  cdsc=2.8125e-7
+  cdscb=1.0e-4
+  cdscd=1.0e-10
+  eta0=0.2
+  etab=-0.00025
+  dsub=1.0
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.030097
+  pdiblc1=0.0
+  pdiblc2=1.735531450e-02 lpdiblc2=-8.223802658e-09 wpdiblc2=-1.183462092e-07 ppdiblc2=1.645027451e-13
+  pdiblcb=-0.025
+  drout=0.43496
+  pscbe1=800000000.0
+  pscbe2=8.6797e-9
+  pvag=0.0
+  delta=5.472932948e-03 ldelta=4.103155882e-09 wdelta=2.935425097e-08 pdelta=1.356209928e-13
+  alpha0=5.0449517e-13
+  alpha1=-4.0583656e-18
+  beta0=6.2016506
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=2300000000.0
+  cgidl=0.5
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-6.299189728e-01 lkt1=1.718337870e-07 wkt1=-1.603804439e-07 pkt1=-5.358395606e-13
+  kt2=5.854481647e-02 lkt2=-9.706392334e-08 wkt2=-1.060535866e-06 pkt2=1.091344433e-12
+  at=9.520047665e+05 lat=-1.102578703e+00 wat=-5.161755040e+00 pat=7.060222050e-6
+  ute=3.557784043e-01 lute=-7.473360381e-07 wute=-2.027993550e-06 pute=3.100903537e-12
+  ua1=5.140280594e-10 lua1=2.017712512e-16 wua1=1.019155418e-15 pua1=-1.396397895e-21
+  ub1=-9.380338003e-21 lub1=-2.384801176e-27 wub1=-7.674625668e-27 pub1=1.173488638e-32
+  uc1=-9.961e-12
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+41
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=1.4472e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=1.0e-11
+  cgso=1.0e-11
+  cgbo=1.0e-13
+  capmod=2.0
+  xpart=0.0
+  cgsl=0.0
+  cgdl=0.0
+  cf=0.0
+  clc=7.0e-8
+  cle=0.492
+  dlc=-5.9781e-8
+  dwc=3.2175e-8
+  vfbcv=-1.0
+  acde=0.44
+  moin=8.7
+  noff=2.6123
+  voffcv=0.112
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000838062107
+  mjs=0.3362
+  pbs=0.6587
+  cjsws=9.9839168e-11
+  mjsws=0.2659
+  pbsws=0.7418
+  cjswgs=2.60659646e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=2.74e-6
+  sbref=2.74e-6
+  wlod={0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.14 pmos
* DC IV MOS Parameters
+  lmin=5e-07 lmax=1e-06 wmin=5.0e-06 wmax=7.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.4525e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=3.9651e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-7.916e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.44996e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.44996e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-7.903706083e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0=1.120070727e-07 wvth0=1.312323173e-06 pvth0=-6.833845194e-13
+  k1=0.64774
+  k2=-2.634852910e-01 lk2=8.696052732e-08 wk2=8.427813251e-07 pk2=-4.077502912e-13
+  k3=3.39
+  dvt0=2.4422
+  dvt1=0.16136
+  dvt2=0.026237
+  dvt0w=0.5
+  dvt1w=1928100.0
+  dvt2w=-0.032
+  w0=1.0e-8
+  k3b=1.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=-1.028507103e+05 lvsat=1.053644098e-01 wvsat=8.487650461e-01 pvsat=-2.212712307e-7
+  ua=-1.737285564e-09 lua=-8.053154274e-16 wua=-7.247918334e-15 pua=4.998384873e-21
+  ub=1.433180830e-18 lub=1.141173327e-24 wub=9.561254609e-24 pub=-6.772663183e-30
+  uc=-2.900706455e-11 luc=6.431223943e-17 wuc=5.983943998e-16 puc=-4.011685901e-22
+  rdsw=484.7
+  prwb=0.1
+  prwg=0.052
+  wr=1.0
+  u0=6.111080558e-03 lu0=-1.564059874e-09 wu0=-1.736481447e-08 pu0=1.046026983e-14
+  a0=6.204592231e-01 la0=-6.230477378e-07 wa0=3.140280325e-06 pa0=4.090893430e-12
+  keta=-0.01258
+  a1=0.0
+  a2=0.46703705
+  ags=2.389767331e+00 lags=-9.374222066e-07 wags=-5.333157481e-06 pags=2.100211567e-12
+  b0=-5.004850223e-07 lb0=5.150241122e-13 wb0=1.742387360e-11 pb0=-1.793003713e-17
+  b1=2.1073e-24
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-2.855213792e-01+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff=5.482089068e-08 wvoff=5.098895135e-07 pvoff=-2.697570471e-13
+  nfactor={2.320798974e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.145398678e-07 wnfactor=1.065336166e-06 pnfactor=-5.636160985e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-6.393105e-11
+  cdsc=2.8125e-7
+  cdscb=1.0e-4
+  cdscd=1.0e-10
+  eta0=0.2
+  etab=-0.00025
+  dsub=1.0
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.030097
+  pdiblc1=0.0
+  pdiblc2=-4.484436000e-02 lpdiblc2=5.578277238e-08 wpdiblc2=1.344423645e-07 ppdiblc2=-9.562933671e-14
+  pdiblcb=-0.025
+  drout=0.43496
+  pscbe1=800000000.0
+  pscbe2=8.6797e-9
+  pvag=0.0
+  delta=3.969475540e-03 ldelta=5.650288727e-09 wdelta=1.148980093e-07 pdelta=4.759218832e-14
+  alpha0=5.0449517e-13
+  alpha1=-4.0583656e-18
+  beta0=6.2016506
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=2300000000.0
+  cgidl=0.5
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-3.005446141e-01 lkt1=-1.671088968e-07 wkt1=-1.287893072e-06 pkt1=6.244273091e-13
+  kt2=-1.436728840e-02 lkt2=-2.203372182e-8
+  at=-3.086198170e+05 lat=1.946670250e-01 wat=3.497036052e+00 pat=-1.850106923e-6
+  ute=-3.408128543e-01 lute=-3.050880343e-08 wute=2.027993550e-06 pute=-1.072909987e-12
+  ua1=5.130357165e-10 lua1=2.027924217e-16 wua1=-6.952720239e-16 pua1=3.678336643e-22
+  ub1=6.099594060e-19 lub1=-6.397163647e-25 wub1=7.674625668e-27 pub1=-4.060260709e-33
+  uc1=-2.375269864e-11 luc1=1.419234749e-17 puc1=-2.350988702e-38
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+41
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=1.4472e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=1.0e-11
+  cgso=1.0e-11
+  cgbo=1.0e-13
+  capmod=2.0
+  xpart=0.0
+  cgsl=0.0
+  cgdl=0.0
+  cf=0.0
+  clc=7.0e-8
+  cle=0.492
+  dlc=-5.9781e-8
+  dwc=3.2175e-8
+  vfbcv=-1.0
+  acde=0.44
+  moin=8.7
+  noff=2.6123
+  voffcv=0.112
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000838062107
+  mjs=0.3362
+  pbs=0.6587
+  cjsws=9.9839168e-11
+  mjsws=0.2659
+  pbsws=0.7418
+  cjswgs=2.60659646e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.74e-6
+  sbref=1.74e-6
+  wlod={0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.15 pmos
* DC IV MOS Parameters
+  lmin=3.5e-07 lmax=5e-07 wmin=5.0e-06 wmax=7.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.4525e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=3.9651e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-7.916e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.44996e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.44996e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope3/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-6.077951966e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0=1.541555110e-08 wvth0=1.608745771e-07 pvth0=-7.421063966e-14
+  k1=0.64774
+  k2=-1.258932233e-01 lk2=1.416744389e-08 wk2=2.053606284e-07 pk2=-7.052287168e-14
+  k3=3.39
+  dvt0=2.4422
+  dvt1=0.16136
+  dvt2=0.026237
+  dvt0w=0.5
+  dvt1w=1928100.0
+  dvt2w=-0.032
+  w0=1.0e-8
+  k3b=1.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=3.175514299e+05 lvsat=-1.170493425e-01 wvsat=-5.659989941e-01 pvsat=5.272096848e-7
+  ua=-4.208560399e-09 lua=5.021125243e-16 wua=7.759157859e-15 pua=-2.941108787e-21
+  ub=4.672276971e-18 lub=-5.724704857e-25 wub=-1.142854288e-23 pub=4.331989180e-30
+  uc=1.668906202e-10 luc=-3.932743067e-17 wuc=-5.639202190e-16 puc=2.137539590e-22
+  rdsw=484.7
+  prwb=0.1
+  prwg=0.052
+  wr=1.0
+  u0=2.561725261e-04 lu0=1.533479221e-09 wu0=1.545825759e-08 pu0=-6.904776448e-15
+  a0=-4.492291905e+00 la0=2.081853247e-06 wa0=3.834839157e-05 pa0=-1.453595782e-11
+  keta=-0.01258
+  a1=0.0
+  a2=0.46703705
+  ags=1.131621985e+00 lags=-2.718004111e-07 wags=-4.993226405e-06 pags=1.920371031e-12
+  b0=1.668283408e-06 lb0=-6.323628257e-13 wb0=-5.807957868e-11 pb0=2.201506430e-17
+  b1=2.1073e-24
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-6.393105e-11
+  cdsc=2.8125e-7
+  cdscb=1.0e-4
+  cdscd=1.0e-10
+  eta0=0.2
+  etab=-0.00025
+  dsub=1.0
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.030097
+  pdiblc1=0.0
+  pdiblc2=-1.785943197e-01 lpdiblc2=1.265431886e-07 wpdiblc2=5.244529909e-07 ppdiblc2=-3.019644586e-13
+  pdiblcb=-0.025
+  drout=0.43496
+  pscbe1=800000000.0
+  pscbe2=8.6797e-9
+  pvag=0.0
+  delta=4.309650713e-04 ldelta=7.522337691e-09 wdelta=1.558468656e-07 pdelta=2.592819588e-14
+  alpha0=5.0449517e-13
+  alpha1=-4.0583656e-18
+  beta0=6.2016506
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=2300000000.0
+  cgidl=0.5
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-6.023872462e-01 lkt1=-7.419052341e-09 wkt1=-3.795501368e-07 pkt1=1.438684793e-13
+  kt2=-0.056015
+  at=1.455597670e+05 lat=-4.561668393e-2
+  ute=-0.39848
+  ua1=8.9635e-10
+  ub1=-5.9922e-19
+  uc1=3.0734e-12
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+41
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=1.4472e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=1.0e-11
+  cgso=1.0e-11
+  cgbo=1.0e-13
+  capmod=2.0
+  xpart=0.0
+  cgsl=0.0
+  cgdl=0.0
+  cf=0.0
+  clc=7.0e-8
+  cle=0.492
+  dlc=-5.9781e-8
+  dwc=3.2175e-8
+  vfbcv=-1.0
+  acde=0.44
+  moin=8.7
+  noff=2.6123
+  voffcv=0.112
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000838062107
+  mjs=0.3362
+  pbs=0.6587
+  cjsws=9.9839168e-11
+  mjsws=0.2659
+  pbsws=0.7418
+  cjswgs=2.60659646e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.44e-6
+  sbref=1.44e-6
+  wlod={0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.16 pmos
* DC IV MOS Parameters
+  lmin=2.0e-05 lmax=1.0e-04 wmin=3.0e-06 wmax=5.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.4525e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=3.9651e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-7.916e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.44996e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.44996e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-5.804381686e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0=5.288849193e-8
+  k1=0.64774
+  k2=-8.666535496e-02 wk2=8.544078384e-9
+  k3=3.39
+  dvt0=2.4422
+  dvt1=0.16136
+  dvt2=0.026237
+  dvt0w=0.5
+  dvt1w=1928100.0
+  dvt2w=-0.032
+  w0=1.0e-8
+  k3b=1.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=123760.0
+  ua=-3.104734900e-09 wua=7.185936404e-16
+  ub=3.067824430e-18 wub=-5.030155483e-25
+  uc=3.094818709e-11 wuc=8.756782101e-17
+  rdsw=484.7
+  prwb=0.1
+  prwg=0.052
+  wr=1.0
+  u0=2.418031224e-03 wu0=1.782615244e-9
+  a0=1.774741483e+00 wa0=-1.137246295e-7
+  keta=-0.01258
+  a1=0.0
+  a2=0.46703705
+  ags=4.556815264e-01 wags=1.386885726e-8
+  b0=0.0
+  b1=2.1073e-24
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-6.393105e-11
+  cdsc=2.8125e-7
+  cdscb=1.0e-4
+  cdscd=1.0e-10
+  eta0=0.2
+  etab=-0.00025
+  dsub=1.0
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.030097
+  pdiblc1=0.0
+  pdiblc2=7.632714483e-04 wpdiblc2=4.335275432e-9
+  pdiblcb=-0.025
+  drout=0.43496
+  pscbe1=800000000.0
+  pscbe2=8.6797e-9
+  pvag=0.0
+  delta=1.336714452e-02 wdelta=2.132067331e-8
+  alpha0=5.0449517e-13
+  alpha1=-4.0583656e-18
+  beta0=6.2016506
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=2300000000.0
+  cgidl=0.5
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.60135
+  kt2=-0.055045
+  at=2.897765981e+05 wat=-2.055177811e-2
+  ute=-1.218875050e-01 wute=-4.961170493e-7
+  ua1=6.8217e-10
+  ub1=-1.464640800e-19 wub1=-1.070704524e-26
+  uc1=-9.961e-12
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+41
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=1.4472e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=1.0e-11
+  cgso=1.0e-11
+  cgbo=1.0e-13
+  capmod=2.0
+  xpart=0.0
+  cgsl=0.0
+  cgdl=0.0
+  cf=0.0
+  clc=7.0e-8
+  cle=0.492
+  dlc=-5.9781e-8
+  dwc=3.2175e-8
+  vfbcv=-1.0
+  acde=0.44
+  moin=8.7
+  noff=2.6123
+  voffcv=0.112
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000838062107
+  mjs=0.3362
+  pbs=0.6587
+  cjsws=9.9839168e-11
+  mjsws=0.2659
+  pbsws=0.7418
+  cjswgs=2.60659646e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.17 pmos
* DC IV MOS Parameters
+  lmin=8e-06 lmax=2.0e-05 wmin=3.0e-06 wmax=5.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.4525e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=3.9651e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-7.916e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.44996e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.44996e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-5.804381686e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0=5.288849193e-8
+  k1=0.64774
+  k2=-8.666535496e-02 wk2=8.544078384e-9
+  k3=3.39
+  dvt0=2.4422
+  dvt1=0.16136
+  dvt2=0.026237
+  dvt0w=0.5
+  dvt1w=1928100.0
+  dvt2w=-0.032
+  w0=1.0e-8
+  k3b=1.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=123760.0
+  ua=-3.104734900e-09 wua=7.185936404e-16
+  ub=3.067824430e-18 wub=-5.030155483e-25
+  uc=3.094818709e-11 wuc=8.756782101e-17
+  rdsw=484.7
+  prwb=0.1
+  prwg=0.052
+  wr=1.0
+  u0=2.418031224e-03 wu0=1.782615244e-9
+  a0=1.774741483e+00 wa0=-1.137246295e-7
+  keta=-0.01258
+  a1=0.0
+  a2=0.46703705
+  ags=4.556815264e-01 wags=1.386885726e-8
+  b0=0.0
+  b1=2.1073e-24
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-6.393105e-11
+  cdsc=2.8125e-7
+  cdscb=1.0e-4
+  cdscd=1.0e-10
+  eta0=0.2
+  etab=-0.00025
+  dsub=1.0
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.030097
+  pdiblc1=0.0
+  pdiblc2=7.632714483e-04 wpdiblc2=4.335275432e-9
+  pdiblcb=-0.025
+  drout=0.43496
+  pscbe1=800000000.0
+  pscbe2=8.6797e-9
+  pvag=0.0
+  delta=1.336714452e-02 wdelta=2.132067331e-8
+  alpha0=5.0449517e-13
+  alpha1=-4.0583656e-18
+  beta0=6.2016506
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=2300000000.0
+  cgidl=0.5
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.60135
+  kt2=-0.055045
+  at=2.897765981e+05 wat=-2.055177811e-2
+  ute=-1.218875050e-01 wute=-4.961170493e-7
+  ua1=6.8217e-10
+  ub1=-1.464640800e-19 wub1=-1.070704524e-26
+  uc1=-9.961e-12
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+41
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=1.4472e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=1.0e-11
+  cgso=1.0e-11
+  cgbo=1.0e-13
+  capmod=2.0
+  xpart=0.0
+  cgsl=0.0
+  cgdl=0.0
+  cf=0.0
+  clc=7.0e-8
+  cle=0.492
+  dlc=-5.9781e-8
+  dwc=3.2175e-8
+  vfbcv=-1.0
+  acde=0.44
+  moin=8.7
+  noff=2.6123
+  voffcv=0.112
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000838062107
+  mjs=0.3362
+  pbs=0.6587
+  cjsws=9.9839168e-11
+  mjsws=0.2659
+  pbsws=0.7418
+  cjswgs=2.60659646e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.18 pmos
* DC IV MOS Parameters
+  lmin=4e-06 lmax=8e-06 wmin=3.0e-06 wmax=5.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.4525e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=3.9651e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-7.916e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.44996e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.44996e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-5.660267856e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0=-1.157097147e-07 wvth0=-2.332895660e-08 pvth0=6.119537051e-13
+  k1=0.64774
+  k2=-6.409969449e-02 lk2=-1.811808162e-07 wk2=-5.489808081e-08 pk2=5.093802683e-13
+  k3=3.39
+  dvt0=2.4422
+  dvt1=0.16136
+  dvt2=0.026237
+  dvt0w=0.5
+  dvt1w=1928100.0
+  dvt2w=-0.032
+  w0=1.0e-8
+  k3b=1.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=123760.0
+  ua=-3.148863544e-09 lua=3.543110854e-16 wua=9.357373684e-16 pua=-1.743457849e-21
+  ub=3.067824430e-18 wub=-5.030155483e-25
+  uc=3.094818709e-11 wuc=8.756782101e-17
+  rdsw=484.7
+  prwb=0.1
+  prwg=0.052
+  wr=1.0
+  u0=2.070331750e-03 lu0=2.791696462e-09 wu0=3.277389238e-09 pu0=-1.200161514e-14
+  a0=1.802267960e+00 la0=-2.210114584e-07 wa0=-2.756414694e-07 pa0=1.300038403e-12
+  keta=-0.01258
+  a1=0.0
+  a2=0.46703705
+  ags=4.038249094e-01 lags=4.163593708e-07 wags=-1.674840839e-08 pags=2.458275568e-13
+  b0=0.0
+  b1=2.1073e-24
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-6.393105e-11
+  cdsc=2.8125e-7
+  cdscb=1.0e-4
+  cdscd=1.0e-10
+  eta0=0.2
+  etab=-0.00025
+  dsub=1.0
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.030097
+  pdiblc1=0.0
+  pdiblc2=-1.481179665e-03 lpdiblc2=1.802081021e-08 wpdiblc2=7.991975812e-09 ppdiblc2=-2.935983018e-14
+  pdiblcb=-0.025
+  drout=0.43496
+  pscbe1=800000000.0
+  pscbe2=8.6797e-9
+  pvag=0.0
+  delta=1.183062683e-02 ldelta=1.233677730e-08 wdelta=5.541562408e-09 pdelta=1.266912704e-13
+  alpha0=5.0449517e-13
+  alpha1=-4.0583656e-18
+  beta0=6.2016506
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=2300000000.0
+  cgidl=0.5
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-6.114226250e-01 lkt1=8.087360976e-8
+  kt2=-0.055045
+  at=3.076722262e+05 lat=-1.436848925e-01 wat=-4.125281352e-02 pat=1.662096483e-7
+  ute=-1.107144508e-01 lute=-8.970901086e-08 wute=-9.958371487e-07 pute=4.012277664e-12
+  ua1=6.681489060e-10 lua1=1.125760648e-16
+  ub1=-1.712267019e-19 lub1=1.988203291e-25 wub1=-2.149185040e-26 pub1=8.659173985e-32
+  uc1=-9.961e-12
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+41
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=1.4472e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=1.0e-11
+  cgso=1.0e-11
+  cgbo=1.0e-13
+  capmod=2.0
+  xpart=0.0
+  cgsl=0.0
+  cgdl=0.0
+  cf=0.0
+  clc=7.0e-8
+  cle=0.492
+  dlc=-5.9781e-8
+  dwc=3.2175e-8
+  vfbcv=-1.0
+  acde=0.44
+  moin=8.7
+  noff=2.6123
+  voffcv=0.112
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000838062107
+  mjs=0.3362
+  pbs=0.6587
+  cjsws=9.9839168e-11
+  mjsws=0.2659
+  pbsws=0.7418
+  cjswgs=2.60659646e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.19 pmos
* DC IV MOS Parameters
+  lmin=2e-06 lmax=4e-06 wmin=3.0e-06 wmax=5.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.4525e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=3.9651e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-7.916e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.44996e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.44996e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-5.355479310e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0=-2.385105439e-07 wvth0=-5.895042572e-08 pvth0=7.554743853e-13
+  k1=0.64774
+  k2=-1.178826415e-01 lk2=3.551336647e-08 wk2=1.131492029e-07 pk2=-1.676906402e-13
+  k3=3.39
+  dvt0=2.4422
+  dvt1=0.16136
+  dvt2=0.026237
+  dvt0w=0.5
+  dvt1w=1928100.0
+  dvt2w=-0.032
+  w0=1.0e-8
+  k3b=1.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=123760.0
+  ua=-2.913156164e-09 lua=-5.953657309e-16 wua=7.142907016e-17 pua=1.738883500e-21
+  ub=2.771788681e-18 lub=1.192742833e-24 wub=3.616154703e-25 pub=-3.483641605e-30
+  uc=-1.746924586e-12 luc=1.317302397e-16 wuc=2.119478363e-16 puc=-5.011333004e-22
+  rdsw=484.7
+  prwb=0.1
+  prwg=0.052
+  wr=1.0
+  u0=2.426467841e-03 lu0=1.356806341e-09 wu0=1.232077629e-09 pu0=-3.760952401e-15
+  a0=1.483877856e+00 la0=1.061798189e-06 wa0=1.527910245e-06 pa0=-5.966561632e-12
+  keta=-0.01258
+  a1=0.0
+  a2=0.46703705
+  ags=4.966782586e-02 lags=1.843275968e-06 wags=1.273120381e-06 pags=-4.951118289e-12
+  b0=0.0
+  b1=2.1073e-24
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-6.393105e-11
+  cdsc=2.8125e-7
+  cdscb=1.0e-4
+  cdscd=1.0e-10
+  eta0=0.2
+  etab=-0.00025
+  dsub=1.0
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.030097
+  pdiblc1=0.0
+  pdiblc2=-1.525378118e-03 lpdiblc2=1.819888799e-08 wpdiblc2=4.318019053e-09 ppdiblc2=-1.455727470e-14
+  pdiblcb=-0.025
+  drout=0.43496
+  pscbe1=800000000.0
+  pscbe2=8.6797e-9
+  pvag=0.0
+  delta=1.265404665e-02 ldelta=9.019177687e-09 wdelta=6.651025897e-09 pdelta=1.222211865e-13
+  alpha0=5.0449517e-13
+  alpha1=-4.0583656e-18
+  beta0=6.2016506
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=2300000000.0
+  cgidl=0.5
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.59135
+  kt2=-0.055045
+  at=2.858375770e+05 lat=-5.571199899e-02 wat=5.416701912e-02 pat=-2.182416284e-7
+  ute=-0.13298
+  ua1=6.9609e-10
+  ub1=-1.2188e-19
+  uc1=-9.961e-12
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+41
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=1.4472e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=1.0e-11
+  cgso=1.0e-11
+  cgbo=1.0e-13
+  capmod=2.0
+  xpart=0.0
+  cgsl=0.0
+  cgdl=0.0
+  cf=0.0
+  clc=7.0e-8
+  cle=0.492
+  dlc=-5.9781e-8
+  dwc=3.2175e-8
+  vfbcv=-1.0
+  acde=0.44
+  moin=8.7
+  noff=2.6123
+  voffcv=0.112
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000838062107
+  mjs=0.3362
+  pbs=0.6587
+  cjsws=9.9839168e-11
+  mjsws=0.2659
+  pbsws=0.7418
+  cjswgs=2.60659646e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.20 pmos
* DC IV MOS Parameters
+  lmin=1.5e-06 lmax=2e-06 wmin=3.0e-06 wmax=5.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.4525e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=3.9651e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-7.916e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.44996e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.44996e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-8.408099814e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0=3.808814195e-07 wvth0=8.051861717e-07 pvth0=-9.979019777e-13
+  k1=0.64774
+  k2=-1.325280863e-01 lk2=6.522970632e-08 wk2=1.173067829e-07 pk2=-1.761265778e-13
+  k3=3.39
+  dvt0=2.4422
+  dvt1=0.16136
+  dvt2=0.026237
+  dvt0w=0.5
+  dvt1w=1928100.0
+  dvt2w=-0.032
+  w0=1.0e-8
+  k3b=1.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=5.238709145e+05 lvsat=-8.118450510e-01 wvsat=-1.168603148e+00 pvsat=2.371154217e-6
+  ua=-2.997410078e-09 lua=-4.244103279e-16 wua=3.175093065e-16 pua=1.239574396e-21
+  ub=2.881848248e-18 lub=9.694264685e-25 wub=4.016471364e-26 pub=-2.831401948e-30
+  uc=-3.454642331e-11 luc=1.982820626e-16 wuc=2.503839138e-16 puc=-5.791220235e-22
+  rdsw=484.7
+  prwb=0.1
+  prwg=0.052
+  wr=1.0
+  u0=3.713007035e-03 lu0=-1.253646009e-09 wu0=-2.287841652e-09 pu0=3.381139815e-15
+  a0=-8.087779112e-01 la0=5.713711374e-06 wa0=7.911211212e-06 pa0=-1.891859846e-11
+  keta=-0.01258
+  a1=0.0
+  a2=0.46703705
+  ags=1.375084975e-01 lags=1.665042854e-06 wags=5.747671664e-07 pags=-3.534124699e-12
+  b0=0.0
+  b1=2.1073e-24
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-6.393105e-11
+  cdsc=2.8125e-7
+  cdscb=1.0e-4
+  cdscd=1.0e-10
+  eta0=0.2
+  etab=-0.00025
+  dsub=1.0
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.030097
+  pdiblc1=0.0
+  pdiblc2=-7.646509209e-03 lpdiblc2=3.061896903e-08 wpdiblc2=2.735744691e-08 ppdiblc2=-6.130542579e-14
+  pdiblcb=-0.025
+  drout=0.43496
+  pscbe1=800000000.0
+  pscbe2=8.6797e-9
+  pvag=0.0
+  delta=-1.423514152e-02 ldelta=6.357868494e-08 wdelta=1.991780750e-07 pdelta=-2.684258224e-13
+  alpha0=5.0449517e-13
+  alpha1=-4.0583656e-18
+  beta0=6.2016506
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=2300000000.0
+  cgidl=0.5
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-3.656302017e-01 lkt1=-4.579967568e-07 wkt1=-6.592593635e-07 pkt1=1.337670211e-12
+  kt2=9.819617107e-02 lkt2=-3.109339982e-07 wkt2=-4.475711819e-07 pkt2=9.081443066e-13
+  at=1.119225344e+06 lat=-1.746697447e+00 wat=-2.374643726e+00 pat=4.709936815e-6
+  ute=-0.13298
+  ua1=9.111257279e-10 lua1=-4.363182436e-16 wua1=-6.280544203e-16 pua1=1.274353821e-21
+  ub1=-9.565918141e-19 lub1=1.693672006e-24 wub1=2.437941126e-24 pub1=-4.946704442e-30
+  uc1=-9.961e-12
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+41
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=1.4472e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=1.0e-11
+  cgso=1.0e-11
+  cgbo=1.0e-13
+  capmod=2.0
+  xpart=0.0
+  cgsl=0.0
+  cgdl=0.0
+  cf=0.0
+  clc=7.0e-8
+  cle=0.492
+  dlc=-5.9781e-8
+  dwc=3.2175e-8
+  vfbcv=-1.0
+  acde=0.44
+  moin=8.7
+  noff=2.6123
+  voffcv=0.112
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000838062107
+  mjs=0.3362
+  pbs=0.6587
+  cjsws=9.9839168e-11
+  mjsws=0.2659
+  pbsws=0.7418
+  cjswgs=2.60659646e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.21 pmos
* DC IV MOS Parameters
+  lmin=1e-06 lmax=1.5e-06 wmin=3.0e-06 wmax=5.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.4525e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=3.9651e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-7.916e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.44996e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.44996e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-6.504345252e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0=8.978782820e-08 wvth0=3.309173009e-07 pvth0=-2.727211609e-13
+  k1=0.64774
+  k2=-1.536999888e-01 lk2=9.760260373e-08 wk2=3.040153777e-07 pk2=-4.616133547e-13
+  k3=3.39
+  dvt0=2.4422
+  dvt1=0.16136
+  dvt2=0.026237
+  dvt0w=0.5
+  dvt1w=1928100.0
+  dvt2w=-0.032
+  w0=1.0e-8
+  k3b=1.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=-2.994917688e+05 lvsat=4.471176599e-01 wvsat=1.236190595e+00 pvsat=-1.305895655e-6
+  ua=-3.156828990e-09 lua=-1.806508405e-16 wua=1.417406554e-16 pua=1.508333452e-21
+  ub=3.624354131e-18 lub=-1.659021519e-25 wub=-2.345471031e-24 pub=8.163543871e-31
+  uc=1.316998896e-10 luc=-5.591686226e-17 wuc=-3.774598371e-16 puc=3.808824638e-22
+  rdsw=484.7
+  prwb=0.1
+  prwg=0.052
+  wr=1.0
+  u0=3.880060310e-03 lu0=-1.509078820e-09 wu0=-7.469279418e-09 pu0=1.130381723e-14
+  a0=5.345603572e+00 la0=-3.696645632e-06 wa0=-1.068431345e-05 pa0=9.514888530e-12
+  keta=-0.01258
+  a1=0.0
+  a2=0.46703705
+  ags=1.841386323e+00 lags=-9.402715361e-07 wags=-4.116459731e-06 pags=3.638995789e-12
+  b0=0.0
+  b1=2.1073e-24
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={6.826812792e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-6.558879535e-06 wnfactor=-2.110739702e-05 pnfactor=3.227426541e-11
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-6.393105e-11
+  cdsc=2.8125e-7
+  cdscb=1.0e-4
+  cdscd=1.0e-10
+  eta0=0.2
+  etab=-0.00025
+  dsub=1.0
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.030097
+  pdiblc1=0.0
+  pdiblc2=-1.559004090e-02 lpdiblc2=4.276502616e-08 wpdiblc2=4.376793516e-08 ppdiblc2=-8.639788286e-14
+  pdiblcb=-0.025
+  drout=0.43496
+  pscbe1=800000000.0
+  pscbe2=8.6797e-9
+  pvag=0.0
+  delta=3.753677100e-02 ldelta=-1.558315789e-08 wdelta=-1.284222128e-07 pdelta=2.324913976e-13
+  alpha0=5.0449517e-13
+  alpha1=-4.0583656e-18
+  beta0=6.2016506
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=2300000000.0
+  cgidl=0.5
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-8.565996838e-01 lkt1=2.927201299e-07 wkt1=9.550468777e-07 pkt1=-1.130684747e-12
+  kt2=-2.479375257e-01 lkt2=2.183217308e-07 wkt2=4.475711819e-07 pkt2=-4.605731247e-13
+  at=-6.550948881e+05 lat=9.663269033e-01 wat=2.746297016e+00 pat=-3.120237627e-6
+  ute=-6.742667849e-01 lute=8.276545584e-07 wute=3.040547753e-06 pute=-4.649149541e-12
+  ua1=5.935088561e-10 lua1=4.933383408e-17 wua1=6.280544203e-16 pua1=-6.462994012e-22
+  ub1=4.845062001e-19 lub1=-5.098389123e-25 wub1=-2.437941126e-24 pub1=2.508763316e-30
+  uc1=-9.961e-12
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+41
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=1.4472e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=1.0e-11
+  cgso=1.0e-11
+  cgbo=1.0e-13
+  capmod=2.0
+  xpart=0.0
+  cgsl=0.0
+  cgdl=0.0
+  cf=0.0
+  clc=7.0e-8
+  cle=0.492
+  dlc=-5.9781e-8
+  dwc=3.2175e-8
+  vfbcv=-1.0
+  acde=0.44
+  moin=8.7
+  noff=2.6123
+  voffcv=0.112
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000838062107
+  mjs=0.3362
+  pbs=0.6587
+  cjsws=9.9839168e-11
+  mjsws=0.2659
+  pbsws=0.7418
+  cjswgs=2.60659646e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=2.74e-6
+  sbref=2.74e-6
+  wlod={0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.22 pmos
* DC IV MOS Parameters
+  lmin=5e-07 lmax=1e-06 wmin=3.0e-06 wmax=5.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.4525e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=3.9651e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-7.916e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.44996e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.44996e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-4.997046705e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0=-6.532072880e-08 wvth0=-1.179561257e-07 pvth0=1.891920388e-13
+  k1=0.64774
+  k2=-2.388971445e-02 lk2=-3.597865906e-08 wk2=-3.361961495e-07 pk2=1.971963173e-13
+  k3=3.39
+  dvt0=2.4422
+  dvt1=0.16136
+  dvt2=0.026237
+  dvt0w=0.5
+  dvt1w=1928100.0
+  dvt2w=-0.032
+  w0=1.0e-8
+  k3b=1.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=-5.318514276e+03 lvsat=1.443986723e-01 wvsat=3.688385642e-01 pvsat=-4.133470479e-7
+  ua=-3.881952907e-09 lua=5.655379262e-16 wua=3.305341971e-15 pua=-1.747170482e-21
+  ub=4.025447164e-18 lub=-5.786469370e-25 wub=-3.194505154e-24 pub=1.690052952e-30
+  uc=1.029317244e-10 luc=-2.631298177e-17 wuc=-5.083653486e-17 puc=4.477075458e-23
+  rdsw=484.7
+  prwb=0.1
+  prwg=0.052
+  wr=1.0
+  u0=7.528886426e-04 lu0=1.708937185e-09 wu0=9.001229771e-09 pu0=-5.645160250e-15
+  a0=1.706751038e+00 la0=4.791556771e-08 wa0=-2.205033636e-06 pa0=7.892856345e-13
+  keta=-0.01258
+  a1=0.0
+  a2=0.46703705
+  ags=1.494686325e+00 lags=-5.834999025e-07 wags=-9.287341631e-07 pags=3.586667931e-13
+  b0=4.389714866e-06 lb0=-4.517236083e-12 wb0=-6.639323204e-12 pb0=6.832195543e-18
+  b1=2.1073e-24
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={4.530899072e-01+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor=1.025576844e-5
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-6.393105e-11
+  cdsc=2.8125e-7
+  cdscb=1.0e-4
+  cdscd=1.0e-10
+  eta0=0.2
+  etab=-0.00025
+  dsub=1.0
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.030097
+  pdiblc1=0.0
+  pdiblc2=-1.243593973e-02 lpdiblc2=3.951929834e-08 wpdiblc2=-2.502968432e-08 ppdiblc2=-1.560169253e-14
+  pdiblcb=-0.025
+  drout=0.43496
+  pscbe1=800000000.0
+  pscbe2=8.6797e-9
+  pvag=0.0
+  delta=2.176107904e-03 ldelta=2.080473246e-08 wdelta=1.237226298e-07 pdelta=-2.697825267e-14
+  alpha0=5.0449517e-13
+  alpha1=-4.0583656e-18
+  beta0=6.2016506
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=2300000000.0
+  cgidl=0.5
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-5.330673870e-01 lkt1=-4.021078014e-08 wkt1=-1.437187281e-07 pkt1=-8.077935669e-28
+  kt2=-6.577959009e-03 lkt2=-3.004933123e-08 wkt2=-3.832893755e-08 pkt2=3.944239319e-14
+  at=5.271204909e+05 lat=-2.502318325e-01 wat=-6.153896098e-01 pat=3.391059950e-7
+  ute=6.338216323e-01 lute=-5.184338272e-07 wute=-2.767888419e-06 pute=1.328021701e-12
+  ua1=3.717403100e-10 lua1=2.775447565e-16
+  ub1=5.559692978e-19 lub1=-5.833780129e-25 wub1=2.733436431e-25 pub1=-2.812842760e-31
+  uc1=-2.375269864e-11 luc1=1.419234749e-17
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+41
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=1.4472e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=1.0e-11
+  cgso=1.0e-11
+  cgbo=1.0e-13
+  capmod=2.0
+  xpart=0.0
+  cgsl=0.0
+  cgdl=0.0
+  cf=0.0
+  clc=7.0e-8
+  cle=0.492
+  dlc=-5.9781e-8
+  dwc=3.2175e-8
+  vfbcv=-1.0
+  acde=0.44
+  moin=8.7
+  noff=2.6123
+  voffcv=0.112
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000838062107
+  mjs=0.3362
+  pbs=0.6587
+  cjsws=9.9839168e-11
+  mjsws=0.2659
+  pbsws=0.7418
+  cjswgs=2.60659646e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.74e-6
+  sbref=1.74e-6
+  wlod={0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.23 pmos
* DC IV MOS Parameters
+  lmin=3.5e-07 lmax=5e-07 wmin=3.0e-06 wmax=5.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.4525e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=3.9651e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-7.916e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.44996e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.44996e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope3/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-5.894845813e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0=-1.782266702e-08 wvth0=7.077356905e-08 pvth0=8.934459377e-14
+  k1=0.64774
+  k2=-8.549974579e-02 lk2=-3.383871979e-09 wk2=6.596524342e-09 pk2=1.584185324e-14
+  k3=3.39
+  dvt0=2.4422
+  dvt1=0.16136
+  dvt2=0.026237
+  dvt0w=0.5
+  dvt1w=1928100.0
+  dvt2w=-0.032
+  w0=1.0e-8
+  k3b=1.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=4.448863602e+05 lvsat=-9.378221657e-02 wvsat=-1.192575731e+00 pvsat=4.127191850e-7
+  ua=-2.885089321e-09 lua=3.814724639e-17 wua=1.246756373e-15 pua=-6.580757713e-22
+  ub=2.697358341e-18 lub=1.239784546e-25 wub=-1.710564734e-24 pub=9.049742724e-31
+  uc=-1.850840351e-11 luc=3.793491788e-17 wuc=3.483723860e-16 puc=-1.664307250e-22
+  rdsw=484.7
+  prwb=0.1
+  prwg=0.052
+  wr=1.0
+  u0=4.093263195e-03 lu0=-5.828797234e-11 wu0=-3.422906787e-09 pu0=9.278291959e-16
+  a0=5.635157179e+00 la0=-2.030407701e-06 wa0=-1.148572688e-05 pa0=5.699236397e-12
+  keta=-0.01258
+  a1=0.0
+  a2=0.46703705
+  ags=-1.591489433e-01 lags=2.914616460e-07 wags=1.358267519e-06 pags=-8.512714466e-13
+  b0=-1.463238289e-05 lb0=5.546404733e-12 wb0=2.213107735e-11 pb0=-8.388784869e-18
+  b1=2.1073e-24
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={4.530899072e-01+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor=1.025576844e-5
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-6.393105e-11
+  cdsc=2.8125e-7
+  cdscb=1.0e-4
+  cdscd=1.0e-10
+  eta0=0.2
+  etab=-0.00025
+  dsub=1.0
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.030097
+  pdiblc1=0.0
+  pdiblc2=-4.106505058e-02 lpdiblc2=5.466552944e-08 wpdiblc2=-1.522870087e-07 ppdiblc2=5.172379493e-14
+  pdiblcb=-0.025
+  drout=0.43496
+  pscbe1=800000000.0
+  pscbe2=8.6797e-9
+  pvag=0.0
+  delta=6.042888853e-02 ldelta=-1.001390113e-08 wdelta=-1.393847964e-07 pdelta=1.122187312e-13
+  alpha0=5.0449517e-13
+  alpha1=-4.0583656e-18
+  beta0=6.2016506
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=2300000000.0
+  cgidl=0.5
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-6.872166792e-01 lkt1=4.134190292e-08 wkt1=3.786988485e-08 pkt1=-9.606945566e-14
+  kt2=-8.197943130e-02 lkt2=9.841817685e-09 wkt2=1.277631252e-07 pkt2=-4.842861260e-14
+  at=1.272234497e+05 lat=-3.866630286e-02 wat=9.022747980e-02 pat=-3.420072622e-8
+  ute=-2.137776579e-01 lute=-7.001142277e-08 wute=-9.088644454e-07 pute=3.445050680e-13
+  ua1=8.9635e-10
+  ub1=-4.140540993e-19 lub1=-7.018713465e-26 wub1=-9.111454772e-25 pub1=3.453696931e-31
+  uc1=3.0734e-12
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+41
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=1.4472e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=1.0e-11
+  cgso=1.0e-11
+  cgbo=1.0e-13
+  capmod=2.0
+  xpart=0.0
+  cgsl=0.0
+  cgdl=0.0
+  cf=0.0
+  clc=7.0e-8
+  cle=0.492
+  dlc=-5.9781e-8
+  dwc=3.2175e-8
+  vfbcv=-1.0
+  acde=0.44
+  moin=8.7
+  noff=2.6123
+  voffcv=0.112
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000838062107
+  mjs=0.3362
+  pbs=0.6587
+  cjsws=9.9839168e-11
+  mjsws=0.2659
+  pbsws=0.7418
+  cjswgs=2.60659646e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.44e-6
+  sbref=1.44e-6
+  wlod={0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.24 pmos
* DC IV MOS Parameters
+  lmin=2.0e-05 lmax=1.0e-04 wmin=1e-06 wmax=3.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.4525e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=3.9651e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-7.916e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.44996e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.44996e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-5.789992373e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0=4.868580801e-8
+  k1=0.64774
+  k2=-8.380721095e-02 wk2=1.963028989e-10
+  k3=3.39
+  dvt0=2.4422
+  dvt1=0.16136
+  dvt2=0.026237
+  dvt0w=0.5
+  dvt1w=1928100.0
+  dvt2w=-0.032
+  w0=1.0e-8
+  k3b=1.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=123760.0
+  ua=-2.845994368e-09 wua=-3.710931514e-17
+  ub=2.875160504e-18 wub=5.969759392e-26
+  uc=5.924696406e-11 wuc=4.915639716e-18
+  rdsw=484.7
+  prwb=0.1
+  prwg=0.052
+  wr=1.0
+  u0=3.232196885e-03 wu0=-5.953167763e-10
+  a0=1.892252227e+00 wa0=-4.569380225e-7
+  keta=-0.01258
+  a1=0.0
+  a2=0.46703705
+  ags=4.306730406e-01 wags=8.691109169e-8
+  b0=0.0
+  b1=2.1073e-24
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-6.393105e-11
+  cdsc=2.8125e-7
+  cdscb=1.0e-4
+  cdscd=1.0e-10
+  eta0=0.2
+  etab=-0.00025
+  dsub=1.0
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.030097
+  pdiblc1=0.0
+  pdiblc2=2.641382535e-03 wpdiblc2=-1.150119861e-9
+  pdiblcb=-0.025
+  drout=0.43496
+  pscbe1=800000000.0
+  pscbe2=8.6797e-9
+  pvag=0.0
+  delta=2.423930824e-02 wdelta=-1.043363353e-8
+  alpha0=5.0449517e-13
+  alpha1=-4.0583656e-18
+  beta0=6.2016506
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=2300000000.0
+  cgidl=0.5
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-5.921430200e-01 wkt1=-2.689080807e-8
+  kt2=-0.055045
+  at=2.866437595e+05 wat=-1.140170262e-2
+  ute=-0.29175
+  ua1=6.8217e-10
+  ub1=-1.5013e-19
+  uc1=-9.961e-12
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+41
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=1.4472e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=1.0e-11
+  cgso=1.0e-11
+  cgbo=1.0e-13
+  capmod=2.0
+  xpart=0.0
+  cgsl=0.0
+  cgdl=0.0
+  cf=0.0
+  clc=7.0e-8
+  cle=0.492
+  dlc=-5.9781e-8
+  dwc=3.2175e-8
+  vfbcv=-1.0
+  acde=0.44
+  moin=8.7
+  noff=2.6123
+  voffcv=0.112
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000838062107
+  mjs=0.3362
+  pbs=0.6587
+  cjsws=9.9839168e-11
+  mjsws=0.2659
+  pbsws=0.7418
+  cjswgs=2.60659646e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.25 pmos
* DC IV MOS Parameters
+  lmin=8e-06 lmax=2.0e-05 wmin=1e-06 wmax=3.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.4525e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=3.9651e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-7.916e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.44996e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.44996e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-5.789992373e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0=4.868580801e-8
+  k1=0.64774
+  k2=-8.380721095e-02 wk2=1.963028989e-10
+  k3=3.39
+  dvt0=2.4422
+  dvt1=0.16136
+  dvt2=0.026237
+  dvt0w=0.5
+  dvt1w=1928100.0
+  dvt2w=-0.032
+  w0=1.0e-8
+  k3b=1.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=123760.0
+  ua=-2.845994368e-09 wua=-3.710931514e-17
+  ub=2.875160504e-18 wub=5.969759392e-26
+  uc=5.924696406e-11 wuc=4.915639716e-18
+  rdsw=484.7
+  prwb=0.1
+  prwg=0.052
+  wr=1.0
+  u0=3.232196885e-03 wu0=-5.953167763e-10
+  a0=1.892252227e+00 wa0=-4.569380225e-7
+  keta=-0.01258
+  a1=0.0
+  a2=0.46703705
+  ags=4.306730406e-01 wags=8.691109169e-8
+  b0=0.0
+  b1=2.1073e-24
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-6.393105e-11
+  cdsc=2.8125e-7
+  cdscb=1.0e-4
+  cdscd=1.0e-10
+  eta0=0.2
+  etab=-0.00025
+  dsub=1.0
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.030097
+  pdiblc1=0.0
+  pdiblc2=2.641382535e-03 wpdiblc2=-1.150119861e-9
+  pdiblcb=-0.025
+  drout=0.43496
+  pscbe1=800000000.0
+  pscbe2=8.6797e-9
+  pvag=0.0
+  delta=2.423930824e-02 wdelta=-1.043363353e-8
+  alpha0=5.0449517e-13
+  alpha1=-4.0583656e-18
+  beta0=6.2016506
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=2300000000.0
+  cgidl=0.5
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-5.921430200e-01 wkt1=-2.689080807e-8
+  kt2=-0.055045
+  at=2.866437595e+05 wat=-1.140170262e-2
+  ute=-0.29175
+  ua1=6.8217e-10
+  ub1=-1.5013e-19
+  uc1=-9.961e-12
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+41
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=1.4472e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=1.0e-11
+  cgso=1.0e-11
+  cgbo=1.0e-13
+  capmod=2.0
+  xpart=0.0
+  cgsl=0.0
+  cgdl=0.0
+  cf=0.0
+  clc=7.0e-8
+  cle=0.492
+  dlc=-5.9781e-8
+  dwc=3.2175e-8
+  vfbcv=-1.0
+  acde=0.44
+  moin=8.7
+  noff=2.6123
+  voffcv=0.112
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000838062107
+  mjs=0.3362
+  pbs=0.6587
+  cjsws=9.9839168e-11
+  mjsws=0.2659
+  pbsws=0.7418
+  cjswgs=2.60659646e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.26 pmos
* DC IV MOS Parameters
+  lmin=4e-06 lmax=8e-06 wmin=1e-06 wmax=3.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.4525e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=3.9651e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-7.916e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.44996e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.44996e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-5.854252118e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0=5.159447050e-08 wvth0=3.332798786e-08 pvth0=1.233087059e-13
+  k1=0.64774
+  k2=-7.884924703e-02 lk2=-3.980774024e-08 wk2=-1.181909220e-08 pk2=9.647220801e-14
+  k3=3.39
+  dvt0=2.4422
+  dvt1=0.16136
+  dvt2=0.026237
+  dvt0w=0.5
+  dvt1w=1928100.0
+  dvt2w=-0.032
+  w0=1.0e-8
+  k3b=1.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=123760.0
+  ua=-2.825050338e-09 lua=-1.681606585e-16 wua=-1.002321257e-17 pua=-2.174756718e-22
+  ub=2.913646964e-18 lub=-3.090097086e-25 wub=-5.270973173e-26 pub=9.025240380e-31
+  uc=5.924696406e-11 wuc=4.915639716e-18
+  rdsw=484.7
+  prwb=0.1
+  prwg=0.052
+  wr=1.0
+  u0=3.468090899e-03 lu0=-1.894004832e-09 wu0=-8.050431142e-10 pu0=1.683903253e-15
+  a0=1.901743330e+00 la0=-7.620454204e-08 wa0=-5.661789828e-07 pa0=8.771011320e-13
+  keta=-0.01258
+  a1=0.0
+  a2=0.46703705
+  ags=3.462015318e-01 lags=6.782259683e-07 wags=1.515520755e-07 pags=-5.190056908e-13
+  b0=0.0
+  b1=2.1073e-24
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-6.393105e-11
+  cdsc=2.8125e-7
+  cdscb=1.0e-4
+  cdscd=1.0e-10
+  eta0=0.2
+  etab=-0.00025
+  dsub=1.0
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.030097
+  pdiblc1=0.0
+  pdiblc2=2.669930835e-03 lpdiblc2=-2.292157300e-10 wpdiblc2=-4.132164323e-09 ppdiblc2=2.394298409e-14
+  pdiblcb=-0.025
+  drout=0.43496
+  pscbe1=800000000.0
+  pscbe2=8.6797e-9
+  pvag=0.0
+  delta=1.862458204e-02 ldelta=4.508091738e-08 wdelta=-1.430152898e-08 pdelta=3.105552593e-14
+  alpha0=5.0449517e-13
+  alpha1=-4.0583656e-18
+  beta0=6.2016506
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=2300000000.0
+  cgidl=0.5
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-5.929417993e-01 lkt1=6.413439001e-09 wkt1=-5.397691064e-08 pkt1=2.174756718e-13
+  kt2=-0.055045
+  at=3.013837967e+05 lat=-1.183484957e-01 wat=-2.288621011e-02 pat=9.220968485e-8
+  ute=-4.516730671e-01 lute=1.284030302e-6
+  ua1=6.681489060e-10 lua1=1.125760648e-16
+  ub1=-1.554139985e-19 lub1=4.242548792e-26 wub1=-6.767598157e-26 pub1=5.433738398e-31
+  uc1=-9.961e-12
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+41
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=1.4472e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=1.0e-11
+  cgso=1.0e-11
+  cgbo=1.0e-13
+  capmod=2.0
+  xpart=0.0
+  cgsl=0.0
+  cgdl=0.0
+  cf=0.0
+  clc=7.0e-8
+  cle=0.492
+  dlc=-5.9781e-8
+  dwc=3.2175e-8
+  vfbcv=-1.0
+  acde=0.44
+  moin=8.7
+  noff=2.6123
+  voffcv=0.112
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000838062107
+  mjs=0.3362
+  pbs=0.6587
+  cjsws=9.9839168e-11
+  mjsws=0.2659
+  pbsws=0.7418
+  cjswgs=2.60659646e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.27 pmos
* DC IV MOS Parameters
+  lmin=2e-06 lmax=4e-06 wmin=1e-06 wmax=3.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.4525e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=3.9651e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-7.916e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.44996e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.44996e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-5.797602261e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0=2.876995996e-08 wvth0=7.018033612e-08 pvth0=-2.517124784e-14
+  k1=0.64774
+  k2=-8.352011458e-02 lk2=-2.098858133e-08 wk2=1.278663924e-08 pk2=-2.665514236e-15
+  k3=3.39
+  dvt0=2.4422
+  dvt1=0.16136
+  dvt2=0.026237
+  dvt0w=0.5
+  dvt1w=1928100.0
+  dvt2w=-0.032
+  w0=1.0e-8
+  k3b=1.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=123760.0
+  ua=-2.843435609e-09 lua=-9.408548301e-17 wua=-1.322036159e-16 pua=2.747952821e-22
+  ub=2.808695885e-18 lub=1.138434344e-25 wub=2.538206735e-25 pub=-3.325022913e-31
+  uc=7.369069805e-11 luc=-5.819452643e-17 wuc=-8.382677281e-18 puc=5.357958409e-23
+  rdsw=484.7
+  prwb=0.1
+  prwg=0.052
+  wr=1.0
+  u0=3.027707242e-03 lu0=-1.196770578e-10 wu0=-5.239610864e-10 pu0=5.514097089e-16
+  a0=2.191899704e+00 la0=-1.245259083e-06 wa0=-5.400077507e-07 pa0=7.716559291e-13
+  keta=-0.01258
+  a1=0.0
+  a2=0.46703705
+  ags=4.529002729e-01 lags=2.483314054e-07 wags=9.540017929e-08 pags=-2.927668935e-13
+  b0=0.0
+  b1=2.1073e-24
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-6.393105e-11
+  cdsc=2.8125e-7
+  cdscb=1.0e-4
+  cdscd=1.0e-10
+  eta0=0.2
+  etab=-0.00025
+  dsub=1.0
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.030097
+  pdiblc1=0.0
+  pdiblc2=-3.795440704e-05 lpdiblc2=1.068098930e-08 wpdiblc2=-2.629640357e-11 ppdiblc2=7.400236946e-15
+  pdiblcb=-0.025
+  drout=0.43496
+  pscbe1=800000000.0
+  pscbe2=8.6797e-9
+  pvag=0.0
+  delta=1.203272971e-02 ldelta=7.163982001e-08 wdelta=8.465705037e-09 pdelta=-6.067479828e-14
+  alpha0=5.0449517e-13
+  alpha1=-4.0583656e-18
+  beta0=6.2016506
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=2300000000.0
+  cgidl=0.5
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.59135
+  kt2=-0.055045
+  at=3.043834928e+05 lat=-1.304344210e-1
+  ute=-1.429185169e-01 lute=4.004278157e-08 wute=2.902740647e-08 pute=-1.169528720e-13
+  ua1=6.9609e-10
+  ub1=-1.682223343e-19 lub1=9.403091343e-26 wub1=1.353519631e-25 pub1=-2.746359008e-31
+  uc1=-9.961e-12
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+41
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=1.4472e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=1.0e-11
+  cgso=1.0e-11
+  cgbo=1.0e-13
+  capmod=2.0
+  xpart=0.0
+  cgsl=0.0
+  cgdl=0.0
+  cf=0.0
+  clc=7.0e-8
+  cle=0.492
+  dlc=-5.9781e-8
+  dwc=3.2175e-8
+  vfbcv=-1.0
+  acde=0.44
+  moin=8.7
+  noff=2.6123
+  voffcv=0.112
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000838062107
+  mjs=0.3362
+  pbs=0.6587
+  cjsws=9.9839168e-11
+  mjsws=0.2659
+  pbsws=0.7418
+  cjswgs=2.60659646e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.28 pmos
* DC IV MOS Parameters
+  lmin=1.5e-06 lmax=2e-06 wmin=1e-06 wmax=3.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.4525e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=3.9651e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-7.916e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.44996e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.44996e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-5.938056420e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0=5.726881116e-08 wvth0=8.376109167e-08 pvth0=-5.272727990e-14
+  k1=0.64774
+  k2=-9.741007728e-02 lk2=7.194847478e-09 wk2=1.473768404e-08 pk2=-6.624281684e-15
+  k3=3.39
+  dvt0=2.4422
+  dvt1=0.16136
+  dvt2=0.026237
+  dvt0w=0.5
+  dvt1w=1928100.0
+  dvt2w=-0.032
+  w0=1.0e-8
+  k3b=1.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=123760.0
+  ua=-2.889804838e-09 wua=3.226896969e-18
+  ub=2.864802652e-18 wub=8.994975300e-26
+  uc=4.501002165e-11 wuc=1.802356411e-17
+  rdsw=484.7
+  prwb=0.1
+  prwg=0.052
+  wr=1.0
+  u0=3.037817259e-03 lu0=-1.401907876e-10 wu0=-3.158162249e-10 pu0=1.290733777e-16
+  a0=2.127843843e+00 la0=-1.115286537e-06 wa0=-6.657740725e-07 pa0=1.026842084e-12
+  keta=-0.01258
+  a1=0.0
+  a2=0.46703705
+  ags=2.478043356e-01 lags=6.644813169e-07 wags=2.526263324e-07 pags=-6.117866195e-13
+  b0=0.0
+  b1=2.1073e-24
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-6.393105e-11
+  cdsc=2.8125e-7
+  cdscb=1.0e-4
+  cdscd=1.0e-10
+  eta0=0.2
+  etab=-0.00025
+  dsub=1.0
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.030097
+  pdiblc1=0.0
+  pdiblc2=-1.704093044e-03 lpdiblc2=1.406166791e-08 wpdiblc2=1.000144390e-08 ppdiblc2=-1.294654952e-14
+  pdiblcb=-0.025
+  drout=0.43496
+  pscbe1=800000000.0
+  pscbe2=8.6797e-9
+  pvag=0.0
+  delta=6.772660727e-02 ldelta=-4.136584224e-08 wdelta=-4.020744077e-08 pdelta=3.808544822e-14
+  alpha0=5.0449517e-13
+  alpha1=-4.0583656e-18
+  beta0=6.2016506
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=2300000000.0
+  cgidl=0.5
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-0.59135
+  kt2=-0.055045
+  at=3.366079537e+05 lat=-1.958194635e-01 wat=-8.885467997e-02 pat=1.802905884e-7
+  ute=-1.231837733e-01 wute=-2.861181979e-8
+  ua1=6.9609e-10
+  ub1=-1.2188e-19
+  uc1=-9.961e-12
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+41
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=1.4472e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=1.0e-11
+  cgso=1.0e-11
+  cgbo=1.0e-13
+  capmod=2.0
+  xpart=0.0
+  cgsl=0.0
+  cgdl=0.0
+  cf=0.0
+  clc=7.0e-8
+  cle=0.492
+  dlc=-5.9781e-8
+  dwc=3.2175e-8
+  vfbcv=-1.0
+  acde=0.44
+  moin=8.7
+  noff=2.6123
+  voffcv=0.112
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000838062107
+  mjs=0.3362
+  pbs=0.6587
+  cjsws=9.9839168e-11
+  mjsws=0.2659
+  pbsws=0.7418
+  cjswgs=2.60659646e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.29 pmos
* DC IV MOS Parameters
+  lmin=1e-06 lmax=1.5e-06 wmin=1e-06 wmax=3.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.4525e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=3.9651e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-7.916e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.44996e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.44996e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-5.501399842e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0=-9.498162958e-09 wvth0=3.798723549e-08 pvth0=1.726323491e-14
+  k1=0.64774
+  k2=-4.471292616e-02 lk2=-7.338173144e-08 wk2=-1.430291816e-08 pk2=3.778025110e-14
+  k3=3.39
+  dvt0=2.4422
+  dvt1=0.16136
+  dvt2=0.026237
+  dvt0w=0.5
+  dvt1w=1928100.0
+  dvt2w=-0.032
+  w0=1.0e-8
+  k3b=1.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=123760.0
+  ua=-3.210496412e-09 lua=4.903534518e-16 wua=2.984869881e-16 pua=-4.514674423e-22
+  ub=2.756302504e-18 lub=1.659021519e-25 wub=1.898456226e-25 pub=-1.527457795e-31
+  uc=-2.613421692e-11 luc=1.087830980e-16 wuc=8.352592228e-17 puc=-1.001563808e-22
+  rdsw=484.7
+  prwb=0.1
+  prwg=0.052
+  wr=1.0
+  u0=7.730282867e-04 lu0=3.322784790e-09 wu0=1.605422800e-09 pu0=-2.808597153e-15
+  a0=1.666148017e+00 la0=-4.093305343e-07 wa0=6.226502821e-08 pa0=-8.636610252e-14
+  keta=-0.01258
+  a1=0.0
+  a2=0.46703705
+  ags=5.392527643e-01 lags=2.188420970e-07 wags=-3.133208492e-07 pags=2.535749186e-13
+  b0=0.0
+  b1=2.1073e-24
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={-1.752212792e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=6.558879535e-06 wnfactor=3.949345849e-06 pnfactor=-6.038747270e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-6.393105e-11
+  cdsc=2.8125e-7
+  cdscb=1.0e-4
+  cdscd=1.0e-10
+  eta0=0.2
+  etab=-0.00025
+  dsub=1.0
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.030097
+  pdiblc1=0.0
+  pdiblc2=3.057559796e-03 lpdiblc2=6.780862630e-09 wpdiblc2=-1.069607488e-08 ppdiblc2=1.870099158e-14
+  pdiblcb=-0.025
+  drout=0.43496
+  pscbe1=800000000.0
+  pscbe2=8.6797e-9
+  pvag=0.0
+  delta=1.039456576e-03 ldelta=6.060214552e-08 wdelta=-2.182457956e-08 pdelta=9.977134292e-15
+  alpha0=5.0449517e-13
+  alpha1=-4.0583656e-18
+  beta0=6.2016506
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=2300000000.0
+  cgidl=0.5
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-5.257414274e-01 lkt1=-1.003187880e-07 wkt1=-1.129017031e-08 pkt1=1.726323491e-14
+  kt2=-9.469635460e-02 lkt2=6.062890375e-8
+  at=2.342394908e+05 lat=-3.929296527e-02 wat=1.488198737e-01 pat=-1.831256879e-7
+  ute=6.022737188e-01 lute=-1.109260778e-06 wute=-6.878415434e-07 pute=1.007995209e-12
+  ua1=8.085445840e-10 lua1=-1.719486817e-16
+  ub1=-3.502056140e-19 lub1=3.491212801e-25
+  uc1=-9.961e-12
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+41
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=1.4472e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=1.0e-11
+  cgso=1.0e-11
+  cgbo=1.0e-13
+  capmod=2.0
+  xpart=0.0
+  cgsl=0.0
+  cgdl=0.0
+  cf=0.0
+  clc=7.0e-8
+  cle=0.492
+  dlc=-5.9781e-8
+  dwc=3.2175e-8
+  vfbcv=-1.0
+  acde=0.44
+  moin=8.7
+  noff=2.6123
+  voffcv=0.112
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000838062107
+  mjs=0.3362
+  pbs=0.6587
+  cjsws=9.9839168e-11
+  mjsws=0.2659
+  pbsws=0.7418
+  cjswgs=2.60659646e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=2.74e-6
+  sbref=2.74e-6
+  wlod={0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.30 pmos
* DC IV MOS Parameters
+  lmin=5e-07 lmax=1e-06 wmin=1e-06 wmax=3.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.4525e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=3.9651e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-7.916e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.44996e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.44996e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-5.842527254e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0=2.560555334e-08 wvth0=1.289832090e-07 pvth0=-7.637617162e-14
+  k1=0.64774
+  k2=-1.600758257e-01 lk2=4.533246028e-08 wk2=6.156235314e-08 pk2=-4.028890633e-14
+  k3=3.39
+  dvt0=2.4422
+  dvt1=0.16136
+  dvt2=0.026237
+  dvt0w=0.5
+  dvt1w=1928100.0
+  dvt2w=-0.032
+  w0=1.0e-8
+  k3b=1.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=1.122854965e+05 lvsat=1.180783780e-02 wvsat=2.535276500e-02 pvsat=-2.608926283e-8
+  ua=-2.707113552e-09 lua=-2.765268020e-17 wua=-1.260089821e-16 pua=-1.463986422e-23
+  ub=2.956488873e-18 lub=-4.009963158e-26 wub=-7.240081165e-26 pub=1.171189137e-31
+  uc=9.139088439e-11 luc=-1.215610751e-17 wuc=-1.712922666e-17 puc=3.422800254e-24
+  rdsw=484.7
+  prwb=0.1
+  prwg=0.052
+  wr=1.0
+  u0=4.405587208e-03 lu0=-4.152999672e-10 wu0=-1.667199622e-09 pu0=5.590949505e-16
+  a0=7.768607084e-01 la0=5.057905703e-07 wa0=5.108951894e-07 pa0=-5.480289699e-13
+  keta=-0.01258
+  a1=0.0
+  a2=0.46703705
+  ags=1.200009075e+00 lags=-4.611091849e-07 wags=-6.807091021e-08 pags=1.200468866e-15
+  b0=2.724792270e-06 lb0=-2.803947485e-12 wb0=-1.776587108e-12 pb0=1.828196964e-18
+  b1=2.366065308e-07 lb1=-2.434799505e-13 wb1=-6.910562212e-13 pb1=7.111314044e-19
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={4.621510093e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor=-1.918928064e-6
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-6.393105e-11
+  cdsc=2.8125e-7
+  cdscb=1.0e-4
+  cdscd=1.0e-10
+  eta0=0.2
+  etab=-0.00025
+  dsub=1.0
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.030097
+  pdiblc1=0.0
+  pdiblc2=-2.337670872e-02 lpdiblc2=3.398304665e-08 wpdiblc2=6.924997802e-09 ppdiblc2=5.680267317e-16
+  pdiblcb=-0.025
+  drout=0.43496
+  pscbe1=800000000.0
+  pscbe2=8.6797e-9
+  pvag=0.0
+  delta=5.085761501e-02 ldelta=9.336769589e-09 wdelta=-1.846135063e-08 pdelta=6.516203563e-15
+  alpha0=5.0449517e-13
+  alpha1=-4.0583656e-18
+  beta0=6.2016506
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=2300000000.0
+  cgidl=0.5
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-5.763980341e-01 lkt1=-4.819060682e-08 wkt1=-1.716299371e-08 pkt1=2.330666383e-14
+  kt2=-1.970117050e-02 lkt2=-1.654489045e-8
+  at=3.358858563e+05 lat=-1.438921577e-01 wat=-5.685099496e-02 pat=2.851991948e-8
+  ute=-4.220852255e-01 lute=-5.514420659e-08 wute=3.160966287e-07 pute=-2.510736713e-14
+  ua1=3.717403100e-10 lua1=2.775447565e-16
+  ub1=6.495577630e-19 lub1=-6.796852230e-25 pub1=7.115968764e-47
+  uc1=-2.375269864e-11 luc1=1.419234749e-17 wuc1=3.081487911e-33
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+41
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=1.4472e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=1.0e-11
+  cgso=1.0e-11
+  cgbo=1.0e-13
+  capmod=2.0
+  xpart=0.0
+  cgsl=0.0
+  cgdl=0.0
+  cf=0.0
+  clc=7.0e-8
+  cle=0.492
+  dlc=-5.9781e-8
+  dwc=3.2175e-8
+  vfbcv=-1.0
+  acde=0.44
+  moin=8.7
+  noff=2.6123
+  voffcv=0.112
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000838062107
+  mjs=0.3362
+  pbs=0.6587
+  cjsws=9.9839168e-11
+  mjsws=0.2659
+  pbsws=0.7418
+  cjswgs=2.60659646e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.74e-6
+  sbref=1.74e-6
+  wlod={0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.31 pmos
* DC IV MOS Parameters
+  lmin=3.5e-07 lmax=5e-07 wmin=1e-06 wmax=3.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.4525e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=3.9651e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-7.916e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.44996e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.44996e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope3/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-5.855674667e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0=2.630111726e-08 wvth0=5.933286044e-08 pvth0=-3.952765473e-14
+  k1=0.64774
+  k2=-8.047438114e-02 lk2=3.219316063e-09 wk2=-8.081048162e-09 pk2=-3.444064869e-15
+  k3=3.39
+  dvt0=2.4422
+  dvt1=0.16136
+  dvt2=0.026237
+  dvt0w=0.5
+  dvt1w=1928100.0
+  dvt2w=-0.032
+  w0=1.0e-8
+  k3b=1.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=5.931577528e+04 lvsat=3.983146883e-02 wvsat=-6.644049483e-02 pvsat=2.247396129e-8
+  ua=-2.289271917e-09 lua=-2.487117972e-16 wua=-4.934463281e-16 pua=1.797528637e-22
+  ub=1.942141365e-18 lub=4.965409176e-25 wub=4.951959785e-25 pub=-1.831681681e-31
+  uc=1.209930687e-10 luc=-2.781714310e-17 wuc=-5.906928481e-17 puc=2.561118802e-23
+  rdsw=484.7
+  prwb=0.1
+  prwg=0.052
+  wr=1.0
+  u0=3.090874518e-03 lu0=2.802487812e-10 wu0=-4.952321830e-10 pu0=-6.093442327e-17
+  a0=1.951184927e+00 la0=-1.154856576e-07 wa0=-7.259564954e-07 pa0=1.063274139e-13
+  keta=-1.170170705e-02 lketa=-4.646608862e-10 wketa=-2.565228468e-09 pketa=1.357134121e-15
+  a1=0.0
+  a2=0.46703705
+  ags=3.284294801e-01 wags=-6.580180735e-8
+  b0=-9.554429628e-06 lb0=3.692374859e-12 wb0=7.299909422e-12 pb0=-2.973723525e-18
+  b1=-5.981628469e-07 lb1=1.981547888e-13 wb1=1.747053031e-12 pb1=-5.787502953e-19
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={4.621510093e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor=-1.918928064e-6
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-6.393105e-11
+  cdsc=2.8125e-7
+  cdscb=1.0e-4
+  cdscd=1.0e-10
+  eta0=0.2
+  etab=-0.00025
+  dsub=1.0
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.030097
+  pdiblc1=0.0
+  pdiblc2=-1.093536695e-01 lpdiblc2=7.946915773e-08 wpdiblc2=4.716342391e-08 ppdiblc2=-2.072011260e-14
+  pdiblcb=-0.025
+  drout=0.43496
+  pscbe1=800000000.0
+  pscbe2=8.6797e-9
+  pvag=0.0
+  delta=-2.141797656e-02 ldelta=4.757417130e-08 wdelta=9.966517876e-08 pdelta=-5.597863681e-14
+  alpha0=5.0449517e-13
+  alpha1=-4.0583656e-18
+  beta0=6.2016506
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=2300000000.0
+  cgidl=0.5
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-6.783390915e-01 lkt1=5.741309610e-09 wkt1=1.194113223e-08 pkt1=7.909126003e-15
+  kt2=-7.234805859e-02 lkt2=1.130794570e-08 wkt2=9.963279416e-08 pkt2=-5.271072975e-14
+  at=1.597401410e+05 lat=-5.070226701e-02 wat=-4.743955351e-03 pat=9.526901776e-10
+  ute=-6.328382875e-01 lute=5.635470083e-08 wute=3.150850974e-07 pute=-2.457221647e-14
+  ua1=6.948893730e-10 lua1=1.065827447e-16 wua1=5.884056504e-16 pua1=-3.112960094e-22
+  ub1=-2.993746697e-19 lub1=-1.776525195e-25 wub1=-1.246089458e-24 pub1=6.592436276e-31
+  uc1=3.439716556e-11 luc1=-1.657183817e-17 wuc1=-9.148725942e-17 puc1=4.840133460e-23
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+41
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=1.4472e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=1.0e-11
+  cgso=1.0e-11
+  cgbo=1.0e-13
+  capmod=2.0
+  xpart=0.0
+  cgsl=0.0
+  cgdl=0.0
+  cf=0.0
+  clc=7.0e-8
+  cle=0.492
+  dlc=-5.9781e-8
+  dwc=3.2175e-8
+  vfbcv=-1.0
+  acde=0.44
+  moin=8.7
+  noff=2.6123
+  voffcv=0.112
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000838062107
+  mjs=0.3362
+  pbs=0.6587
+  cjsws=9.9839168e-11
+  mjsws=0.2659
+  pbsws=0.7418
+  cjswgs=2.60659646e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.44e-6
+  sbref=1.44e-6
+  wlod={0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.32 pmos
* DC IV MOS Parameters
+  lmin=2.0e-05 lmax=1.0e-04 wmin=5.5e-07 wmax=1.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.4525e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=3.9651e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-7.916e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.44996e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.44996e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-5.663176092e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0=3.700985840e-8
+  k1=0.64774
+  k2=-1.059354191e-01 wk2=2.056969986e-8
+  k3=3.39
+  dvt0=2.4422
+  dvt1=0.16136
+  dvt2=0.026237
+  dvt0w=0.5
+  dvt1w=1928100.0
+  dvt2w=-0.032
+  w0=1.0e-8
+  k3b=1.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=123760.0
+  ua=-2.735362841e-09 wua=-1.389675401e-16
+  ub=2.796698609e-18 wub=1.319373042e-25
+  uc=6.931494591e-11 wuc=-4.353931038e-18
+  rdsw=484.7
+  prwb=0.1
+  prwg=0.052
+  wr=1.0
+  u0=2.678126491e-03 wu0=-8.518527230e-11
+  a0=1.052930080e+00 wa0=3.158241996e-7
+  keta=-0.01258
+  a1=0.0
+  a2=0.46703705
+  ags=7.975100024e-01 wags=-2.508349653e-7
+  b0=2.867073818e-07 wb0=-2.639709130e-13
+  b1=-2.047222501e-07 wb1=1.884873663e-13
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-6.393105e-11
+  cdsc=2.8125e-7
+  cdscb=1.0e-4
+  cdscd=1.0e-10
+  eta0=0.2
+  etab=-0.00025
+  dsub=1.0
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.030097
+  pdiblc1=0.0
+  pdiblc2=2.395602617e-03 wpdiblc2=-9.238307822e-10
+  pdiblcb=-0.025
+  drout=0.43496
+  pscbe1=800000000.0
+  pscbe2=8.6797e-9
+  pvag=0.0
+  delta=1.220932096e-02 wdelta=6.423516927e-10
+  alpha0=5.0449517e-13
+  alpha1=-4.0583656e-18
+  beta0=6.2016506
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=2300000000.0
+  cgidl=0.5
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-5.657030364e-01 wkt1=-5.123404805e-8
+  kt2=-0.055045
+  at=2.659443353e+05 wat=7.656215827e-3
+  ute=-2.978481541e-01 wute=5.614558273e-9
+  ua1=6.8217e-10
+  ub1=-1.5013e-19
+  uc1=-9.961e-12
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+41
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=1.4472e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=1.0e-11
+  cgso=1.0e-11
+  cgbo=1.0e-13
+  capmod=2.0
+  xpart=0.0
+  cgsl=0.0
+  cgdl=0.0
+  cf=0.0
+  clc=7.0e-8
+  cle=0.492
+  dlc=-5.9781e-8
+  dwc=3.2175e-8
+  vfbcv=-1.0
+  acde=0.44
+  moin=8.7
+  noff=2.6123
+  voffcv=0.112
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000838062107
+  mjs=0.3362
+  pbs=0.6587
+  cjsws=9.9839168e-11
+  mjsws=0.2659
+  pbsws=0.7418
+  cjswgs=2.60659646e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.33 pmos
* DC IV MOS Parameters
+  lmin=8e-06 lmax=2.0e-05 wmin=5.5e-07 wmax=1.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.4525e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=3.9651e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-7.916e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.44996e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.44996e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-5.663176092e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} wvth0=3.700985840e-8
+  k1=0.64774
+  k2=-1.059354191e-01 wk2=2.056969986e-8
+  k3=3.39
+  dvt0=2.4422
+  dvt1=0.16136
+  dvt2=0.026237
+  dvt0w=0.5
+  dvt1w=1928100.0
+  dvt2w=-0.032
+  w0=1.0e-8
+  k3b=1.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=123760.0
+  ua=-2.735362841e-09 wua=-1.389675401e-16
+  ub=2.796698609e-18 wub=1.319373042e-25
+  uc=6.931494591e-11 wuc=-4.353931038e-18
+  rdsw=484.7
+  prwb=0.1
+  prwg=0.052
+  wr=1.0
+  u0=2.678126491e-03 wu0=-8.518527230e-11
+  a0=1.052930080e+00 wa0=3.158241996e-7
+  keta=-0.01258
+  a1=0.0
+  a2=0.46703705
+  ags=7.975100024e-01 wags=-2.508349653e-7
+  b0=2.867073818e-07 wb0=-2.639709130e-13
+  b1=-2.047222501e-07 wb1=1.884873663e-13
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-6.393105e-11
+  cdsc=2.8125e-7
+  cdscb=1.0e-4
+  cdscd=1.0e-10
+  eta0=0.2
+  etab=-0.00025
+  dsub=1.0
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.030097
+  pdiblc1=0.0
+  pdiblc2=2.395602617e-03 wpdiblc2=-9.238307822e-10
+  pdiblcb=-0.025
+  drout=0.43496
+  pscbe1=800000000.0
+  pscbe2=8.6797e-9
+  pvag=0.0
+  delta=1.220932096e-02 wdelta=6.423516927e-10
+  alpha0=5.0449517e-13
+  alpha1=-4.0583656e-18
+  beta0=6.2016506
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=2300000000.0
+  cgidl=0.5
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-5.657030364e-01 wkt1=-5.123404805e-8
+  kt2=-0.055045
+  at=2.659443353e+05 wat=7.656215827e-3
+  ute=-2.978481541e-01 wute=5.614558273e-9
+  ua1=6.8217e-10
+  ub1=-1.5013e-19
+  uc1=-9.961e-12
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+41
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=1.4472e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=1.0e-11
+  cgso=1.0e-11
+  cgbo=1.0e-13
+  capmod=2.0
+  xpart=0.0
+  cgsl=0.0
+  cgdl=0.0
+  cf=0.0
+  clc=7.0e-8
+  cle=0.492
+  dlc=-5.9781e-8
+  dwc=3.2175e-8
+  vfbcv=-1.0
+  acde=0.44
+  moin=8.7
+  noff=2.6123
+  voffcv=0.112
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000838062107
+  mjs=0.3362
+  pbs=0.6587
+  cjsws=9.9839168e-11
+  mjsws=0.2659
+  pbsws=0.7418
+  cjswgs=2.60659646e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.34 pmos
* DC IV MOS Parameters
+  lmin=4e-06 lmax=8e-06 wmin=5.5e-07 wmax=1.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.4525e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=3.9651e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-7.916e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.44996e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.44996e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-6.262261829e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0=4.810089340e-07 wvth0=7.089336041e-08 pvth0=-2.720523318e-13
+  k1=0.64774
+  k2=-1.327743302e-01 lk2=2.154909594e-07 wk2=3.782962403e-08 pk2=-1.385807942e-13
+  k3=3.39
+  dvt0=2.4422
+  dvt1=0.16136
+  dvt2=0.026237
+  dvt0w=0.5
+  dvt1w=1928100.0
+  dvt2w=-0.032
+  w0=1.0e-8
+  k3b=1.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=123760.0
+  ua=-2.674779873e-09 lua=-4.864236821e-16 wua=-1.483769294e-16 pua=7.554845745e-23
+  ub=2.658098314e-18 lub=1.112828699e-24 wub=1.825733994e-25 pub=-4.065597401e-31
+  uc=6.361922702e-11 luc=4.573121170e-17 wuc=8.901059460e-19 puc=-4.210463515e-23
+  rdsw=484.7
+  prwb=0.1
+  prwg=0.052
+  wr=1.0
+  u0=2.523360383e-03 lu0=1.242624817e-09 wu0=6.476838239e-11 pu0=-1.203985391e-15
+  a0=7.932422176e-01 la0=2.085046828e-06 wa0=4.544157742e-07 pa0=-1.112758682e-12
+  keta=-0.01258
+  a1=0.0
+  a2=0.46703705
+  ags=7.404502544e-01 lags=4.581355699e-07 wags=-2.114319349e-07 pags=-3.163689012e-13
+  b0=7.213281504e-08 lb0=1.722829925e-12 wb0=-6.641253854e-14 pb0=-1.586206066e-18
+  b1=-2.258573076e-07 lb1=1.696944334e-13 wb1=2.079463714e-13 pb1=-1.562373254e-19
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-6.393105e-11
+  cdsc=2.8125e-7
+  cdscb=1.0e-4
+  cdscd=1.0e-10
+  eta0=0.2
+  etab=-0.00025
+  dsub=1.0
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.030097
+  pdiblc1=0.0
+  pdiblc2=-1.386866005e-03 lpdiblc2=3.036962968e-08 wpdiblc2=-3.970795867e-10 ppdiblc2=-4.229311687e-15
+  pdiblcb=-0.025
+  drout=0.43496
+  pscbe1=800000000.0
+  pscbe2=8.6797e-9
+  pvag=0.0
+  delta=-3.154668088e-03 ldelta=1.233582363e-07 wdelta=5.750583058e-09 pdelta=-4.101424504e-14
+  alpha0=5.0449517e-13
+  alpha1=-4.0583656e-18
+  beta0=6.2016506
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=2300000000.0
+  cgidl=0.5
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-5.959419833e-01 lkt1=2.427900161e-07 wkt1=-5.121464725e-08 pkt1=-1.557700154e-16
+  kt2=-0.055045
+  at=2.569372405e+05 lat=7.231841472e-02 wat=1.803564530e-02 pat=-8.333695821e-8
+  ute=-4.246842150e-01 lute=1.018373075e-06 wute=-2.484858221e-08 pute=2.445900781e-13
+  ua1=6.681489060e-10 lua1=1.125760648e-16
+  ub1=-2.815681308e-19 lub1=1.055323324e-24 wub1=4.847387572e-26 pub1=-3.891991719e-31
+  uc1=-9.961e-12
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+41
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=1.4472e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=1.0e-11
+  cgso=1.0e-11
+  cgbo=1.0e-13
+  capmod=2.0
+  xpart=0.0
+  cgsl=0.0
+  cgdl=0.0
+  cf=0.0
+  clc=7.0e-8
+  cle=0.492
+  dlc=-5.9781e-8
+  dwc=3.2175e-8
+  vfbcv=-1.0
+  acde=0.44
+  moin=8.7
+  noff=2.6123
+  voffcv=0.112
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000838062107
+  mjs=0.3362
+  pbs=0.6587
+  cjsws=9.9839168e-11
+  mjsws=0.2659
+  pbsws=0.7418
+  cjswgs=2.60659646e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.35 pmos
* DC IV MOS Parameters
+  lmin=2e-06 lmax=4e-06 wmin=5.5e-07 wmax=1.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.4525e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=3.9651e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-7.916e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.44996e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.44996e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-4.866832918e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0=-8.121635169e-08 wvth0=-1.551541118e-08 pvth0=7.609292933e-14
+  k1=0.64774
+  k2=-6.101840430e-02 lk2=-7.361725383e-08 wk2=-7.930640412e-09 pk2=4.578959928e-14
+  k3=3.39
+  dvt0=2.4422
+  dvt1=0.16136
+  dvt2=0.026237
+  dvt0w=0.5
+  dvt1w=1928100.0
+  dvt2w=-0.032
+  w0=1.0e-8
+  k3b=1.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=123760.0
+  ua=-2.909906567e-09 lua=4.609135232e-16 wua=-7.100393819e-17 pua=-2.361911930e-22
+  ub=3.081104025e-18 lub=-5.914824616e-25 wub=3.015044277e-27 pub=3.168898506e-31
+  uc=7.496959788e-11 wuc=-9.560157801e-18
+  rdsw=484.7
+  prwb=0.1
+  prwg=0.052
+  wr=1.0
+  u0=2.610662560e-03 lu0=8.908799796e-10 wu0=-1.399888822e-10 pu0=-3.790081343e-16
+  a0=1.517494938e+00 la0=-8.330035955e-07 wa0=8.091536886e-08 pa0=3.920931264e-13
+  keta=-0.01258
+  a1=0.0
+  a2=0.46703705
+  ags=9.754529466e-01 lags=-4.887020271e-07 wags=-3.857130223e-07 pags=3.858183137e-13
+  b0=6.714457706e-07 lb0=-6.918319386e-13 wb0=-6.181987781e-13 pb0=6.369682822e-19
+  b1=-1.773936712e-07 lb1=-2.556798092e-14 wb1=1.633259983e-13 pb1=2.354038890e-20
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-6.393105e-11
+  cdsc=2.8125e-7
+  cdscb=1.0e-4
+  cdscd=1.0e-10
+  eta0=0.2
+  etab=-0.00025
+  dsub=1.0
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.030097
+  pdiblc1=0.0
+  pdiblc2=9.799133174e-04 lpdiblc2=2.083375746e-08 wpdiblc2=-9.634451817e-10 ppdiblc2=-1.947396386e-15
+  pdiblcb=-0.025
+  drout=0.43496
+  pscbe1=800000000.0
+  pscbe2=8.6797e-9
+  pvag=0.0
+  delta=3.144489659e-02 ldelta=-1.604513975e-08 wdelta=-9.407038179e-09 pdelta=2.005656880e-14
+  alpha0=5.0449517e-13
+  alpha1=-4.0583656e-18
+  beta0=6.2016506
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=2300000000.0
+  cgidl=0.5
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-5.356821165e-01 wkt1=-5.125330897e-8
+  kt2=-0.055045
+  at=3.017099639e+05 lat=-1.080731266e-01 wat=2.461512633e-03 pat=-2.058799899e-8
+  ute=-1.277554122e-01 lute=-1.779679181e-07 wute=1.506676632e-08 pute=8.376914311e-14
+  ua1=6.9609e-10
+  ub1=8.408593026e-20 lub1=-4.179151708e-25 wub1=-9.694775144e-26 pub1=1.967118351e-31
+  uc1=-9.961e-12
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+41
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=1.4472e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=1.0e-11
+  cgso=1.0e-11
+  cgbo=1.0e-13
+  capmod=2.0
+  xpart=0.0
+  cgsl=0.0
+  cgdl=0.0
+  cf=0.0
+  clc=7.0e-8
+  cle=0.492
+  dlc=-5.9781e-8
+  dwc=3.2175e-8
+  vfbcv=-1.0
+  acde=0.44
+  moin=8.7
+  noff=2.6123
+  voffcv=0.112
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000838062107
+  mjs=0.3362
+  pbs=0.6587
+  cjsws=9.9839168e-11
+  mjsws=0.2659
+  pbsws=0.7418
+  cjswgs=2.60659646e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.36 pmos
* DC IV MOS Parameters
+  lmin=1.5e-06 lmax=2e-06 wmin=5.5e-07 wmax=1.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.4525e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=3.9651e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-7.916e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.44996e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.44996e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-5.267100785e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} wvth0=2.198634055e-8
+  k1=0.64774
+  k2=-9.730004045e-02 wk2=1.463637335e-8
+  k3=3.39
+  dvt0=2.4422
+  dvt1=0.16136
+  dvt2=0.026237
+  dvt0w=0.5
+  dvt1w=1928100.0
+  dvt2w=-0.032
+  w0=1.0e-8
+  k3b=1.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=123760.0
+  ua=-2.682749265e-09 wua=-1.874087547e-16
+  ub=2.789596935e-18 wub=1.591915064e-25
+  uc=7.496959788e-11 wuc=-9.560157801e-18
+  rdsw=484.7
+  prwb=0.1
+  prwg=0.052
+  wr=1.0
+  u0=3.049725166e-03 wu0=-3.267798111e-10
+  a0=1.106956215e+00 wa0=2.741551246e-7
+  keta=-0.01258
+  a1=0.0
+  a2=0.46703705
+  ags=7.346003175e-01 wags=-1.955657545e-7
+  b0=3.304822958e-07 wb0=-3.042743888e-13
+  b1=-1.899946327e-07 wb1=1.749276783e-13
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-6.393105e-11
+  cdsc=2.8125e-7
+  cdscb=1.0e-4
+  cdscd=1.0e-10
+  eta0=0.2
+  etab=-0.00025
+  dsub=1.0
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.030097
+  pdiblc1=0.0
+  pdiblc2=1.124765312e-02 wpdiblc2=-1.923202894e-9
+  pdiblcb=-0.025
+  drout=0.43496
+  pscbe1=800000000.0
+  pscbe2=8.6797e-9
+  pvag=0.0
+  delta=2.353718620e-02 wdelta=4.776708239e-10
+  alpha0=5.0449517e-13
+  alpha1=-4.0583656e-18
+  beta0=6.2016506
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=2300000000.0
+  cgidl=0.5
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-5.356821165e-01 wkt1=-5.125330897e-8
+  kt2=-0.055045
+  at=2.484470445e+05 wat=-7.685107208e-3
+  ute=-2.154653839e-01 wute=5.635167458e-8
+  ua1=6.9609e-10
+  ub1=-1.2188e-19
+  uc1=-9.961e-12
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+41
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=1.4472e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=1.0e-11
+  cgso=1.0e-11
+  cgbo=1.0e-13
+  capmod=2.0
+  xpart=0.0
+  cgsl=0.0
+  cgdl=0.0
+  cf=0.0
+  clc=7.0e-8
+  cle=0.492
+  dlc=-5.9781e-8
+  dwc=3.2175e-8
+  vfbcv=-1.0
+  acde=0.44
+  moin=8.7
+  noff=2.6123
+  voffcv=0.112
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000838062107
+  mjs=0.3362
+  pbs=0.6587
+  cjsws=9.9839168e-11
+  mjsws=0.2659
+  pbsws=0.7418
+  cjswgs=2.60659646e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.37 pmos
* DC IV MOS Parameters
+  lmin=1e-06 lmax=1.5e-06 wmin=5.5e-07 wmax=1.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.4525e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=3.9651e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-7.916e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.44996e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.44996e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-6.001423886e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0=1.122816737e-07 wvth0=8.402434922e-08 pvth0=-9.485921716e-14
+  k1=0.64774
+  k2=-1.172475432e-01 lk2=3.050072901e-08 wk2=5.247955864e-08 pk2=-5.786412247e-14
+  k3=3.39
+  dvt0=2.4422
+  dvt1=0.16136
+  dvt2=0.026237
+  dvt0w=0.5
+  dvt1w=1928100.0
+  dvt2w=-0.032
+  w0=1.0e-8
+  k3b=1.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=5.855710054e+04 lvsat=9.969849342e-02 wvsat=6.003217913e-02 pvsat=-9.179220350e-8
+  ua=-2.009580133e-09 lua=-1.029309261e-15 wua=-8.071942280e-16 pua=9.476829778e-22
+  ub=2.065192033e-18 lub=1.107651315e-24 wub=8.261496508e-25 pub=-1.019812351e-30
+  uc=1.145481540e-10 luc=-6.051759118e-17 wuc=-4.600005523e-17 puc=5.571842516e-23
+  rdsw=484.7
+  prwb=0.1
+  prwg=0.052
+  wr=1.0
+  u0=4.361108121e-03 lu0=-2.005170107e-09 wu0=-1.698115127e-09 pu0=2.096840266e-15
+  a0=9.817333103e-01 la0=1.914720828e-07 wa0=6.924042796e-07 pa0=-6.395238705e-13
+  keta=-1.095466359e-02 lketa=-2.485220633e-09 wketa=-1.496443979e-09 pketa=2.288137666e-15
+  a1=0.0
+  a2=0.46703705
+  ags=3.980510533e-01 lags=5.146006523e-07 wags=-1.833167163e-07 pags=-1.872939176e-14
+  b0=1.999494838e-07 lb0=1.995911961e-13 wb0=-1.840930898e-13 pb0=-1.837632151e-19
+  b1=4.953591402e-07 lb1=-1.047940186e-12 wb1=-4.560761696e-13 pb1=9.648364337e-19
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-6.393105e-11
+  cdsc=2.8125e-7
+  cdscb=1.0e-4
+  cdscd=1.0e-10
+  eta0=0.2
+  etab=-0.00025
+  dsub=1.0
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.030097
+  pdiblc1=0.0
+  pdiblc2=3.039967539e-03 lpdiblc2=1.254996164e-08 wpdiblc2=-1.067987773e-08 ppdiblc2=1.338939366e-14
+  pdiblcb=-0.025
+  drout=0.43496
+  pscbe1=800000000.0
+  pscbe2=8.6797e-9
+  pvag=0.0
+  delta=-5.738684764e-02 ldelta=1.237368939e-07 wdelta=3.196840187e-08 pdelta=-4.815090231e-14
+  alpha0=5.0449517e-13
+  alpha1=-4.0583656e-18
+  beta0=6.2016506
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=2300000000.0
+  cgidl=0.5
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-2.836360978e-01 lkt1=-3.853909649e-07 wkt1=-2.341960630e-07 pkt1=2.797286180e-13
+  kt2=-2.013873113e-01 lkt2=2.237647111e-07 wkt2=9.823015047e-08 pkt2=-1.501988116e-13
+  at=3.056280674e+05 lat=-8.743264300e-02 wat=8.309255405e-02 pat=-1.388035829e-7
+  ute=-2.052953764e-01 lute=-1.555045000e-08 wute=5.568570746e-08 pute=1.018297028e-15
+  ua1=9.844684134e-10 lua1=-4.409450130e-16 wua1=-1.619727179e-16 pua1=2.476643842e-22
+  ub1=-5.289022027e-19 lub1=6.223572990e-25 wub1=1.645255918e-25 pub1=-2.515678562e-31
+  uc1=7.606558034e-11 luc1=-1.315389427e-16 wuc1=-7.920450047e-17 puc1=1.211076414e-22
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+41
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=1.4472e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=1.0e-11
+  cgso=1.0e-11
+  cgbo=1.0e-13
+  capmod=2.0
+  xpart=0.0
+  cgsl=0.0
+  cgdl=0.0
+  cf=0.0
+  clc=7.0e-8
+  cle=0.492
+  dlc=-5.9781e-8
+  dwc=3.2175e-8
+  vfbcv=-1.0
+  acde=0.44
+  moin=8.7
+  noff=2.6123
+  voffcv=0.112
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000838062107
+  mjs=0.3362
+  pbs=0.6587
+  cjsws=9.9839168e-11
+  mjsws=0.2659
+  pbsws=0.7418
+  cjswgs=2.60659646e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=2.74e-6
+  sbref=2.74e-6
+  wlod={0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.38 pmos
* DC IV MOS Parameters
+  lmin=5e-07 lmax=1e-06 wmin=5.5e-07 wmax=1.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.4525e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=3.9651e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-7.916e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.44996e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.44996e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-4.402475431e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0=-5.225811700e-08 wvth0=-3.602074272e-09 pvth0=-4.687246069e-15
+  k1=0.64774
+  k2=-8.147022059e-02 lk2=-6.315924781e-09 wk2=-1.080967023e-08 pk2=7.263658505e-15
+  k3=3.39
+  dvt0=2.4422
+  dvt1=0.16136
+  dvt2=0.026237
+  dvt0w=0.5
+  dvt1w=1928100.0
+  dvt2w=-0.032
+  w0=1.0e-8
+  k3b=1.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=2.081935340e+05 lvsat=-5.428487838e-02 wvsat=-6.294957324e-02 pvsat=3.476216877e-8
+  ua=-3.075528622e-09 lua=6.760503146e-17 wua=2.131900359e-16 pua=-1.023434488e-22
+  ub=3.287355515e-18 lub=-1.500160165e-25 wub=-3.770290676e-25 pub=2.183187095e-31
+  uc=6.652797470e-11 luc=-1.110242571e-17 wuc=5.762004567e-18 puc=2.452677529e-24
+  rdsw=484.7
+  prwb=0.1
+  prwg=0.052
+  wr=1.0
+  u0=2.312748758e-03 lu0=1.026940951e-10 wu0=2.596725526e-10 pu0=8.217885333e-17
+  a0=1.173196622e+00 la0=-5.553237612e-09 wa0=1.459895069e-07 pa0=-7.723574864e-14
+  keta=-1.336972664e-02 wketa=7.270997421e-10
+  a1=0.0
+  a2=0.46703705
+  ags=1.845529671e+00 lags=-9.749272195e-07 wags=-6.624004318e-07 pags=4.742717057e-13
+  b0=2.106052285e-06 lb0=-1.761883891e-12 wb0=-1.206914442e-12 pb0=8.687710971e-19
+  b1=-2.022240091e-06 lb1=1.542795302e-12 wb1=1.388659345e-12 pb1=-9.334886481e-19
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-6.393105e-11
+  cdsc=2.8125e-7
+  cdscb=1.0e-4
+  cdscd=1.0e-10
+  eta0=0.2
+  etab=-0.00025
+  dsub=1.0
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.030097
+  pdiblc1=0.0
+  pdiblc2=9.416624177e-03 lpdiblc2=5.988063131e-09 wpdiblc2=-2.326775821e-08 ppdiblc2=2.634295207e-14
+  pdiblcb=-0.025
+  drout=0.43496
+  pscbe1=800000000.0
+  pscbe2=8.6797e-9
+  pvag=0.0
+  delta=3.367580265e-02 ldelta=3.002887367e-08 wdelta=-2.642090357e-09 pdelta=-1.253497528e-14
+  alpha0=5.0449517e-13
+  alpha1=-4.0583656e-18
+  beta0=6.2016506
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=2300000000.0
+  cgidl=0.5
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-6.502937403e-01 lkt1=-8.081917916e-09 wkt1=5.087263518e-08 pkt1=-1.362132582e-14
+  kt2=4.895570743e-02 lkt2=-3.385077232e-08 wkt2=-6.321225020e-08 pkt2=1.593349083e-14
+  at=4.336676181e+05 lat=-2.191917426e-01 wat=-1.468784675e-01 pat=9.784809673e-8
+  ute=-5.654798730e-02 lute=-1.686189508e-07 wute=-2.045277548e-08 pute=7.936860289e-14
+  ua1=4.146416170e-12 lua1=5.678553383e-16 wua1=3.384429629e-16 pua1=-2.672883720e-22
+  ub1=1.222496144e-18 lub1=-1.179919170e-24 wub1=-5.275032219e-25 pub1=4.605643946e-31
+  uc1=-7.997778252e-11 luc1=2.903747988e-17 wuc1=5.176632227e-17 puc1=-1.366788370e-23
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+41
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=1.4472e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=1.0e-11
+  cgso=1.0e-11
+  cgbo=1.0e-13
+  capmod=2.0
+  xpart=0.0
+  cgsl=0.0
+  cgdl=0.0
+  cf=0.0
+  clc=7.0e-8
+  cle=0.492
+  dlc=-5.9781e-8
+  dwc=3.2175e-8
+  vfbcv=-1.0
+  acde=0.44
+  moin=8.7
+  noff=2.6123
+  voffcv=0.112
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000838062107
+  mjs=0.3362
+  pbs=0.6587
+  cjsws=9.9839168e-11
+  mjsws=0.2659
+  pbsws=0.7418
+  cjswgs=2.60659646e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.74e-6
+  sbref=1.74e-6
+  wlod={0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.39 pmos
* DC IV MOS Parameters
+  lmin=3.5e-07 lmax=5e-07 wmin=5.5e-07 wmax=1.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.4525e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=3.9651e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-7.916e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.44996e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.44996e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope3/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-3.367833652e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0=-1.069958403e-07 wvth0=-1.697221642e-07 pvth0=8.319858753e-14
+  k1=0.64774
+  k2=-4.911887884e-02 lk2=-2.343140213e-08 wk2=-3.694999642e-08 pk2=2.109319807e-14
+  k3=3.39
+  dvt0=2.4422
+  dvt1=0.16136
+  dvt2=0.026237
+  dvt0w=0.5
+  dvt1w=1928100.0
+  dvt2w=-0.032
+  w0=1.0e-8
+  k3b=1.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=-2.864325589e+04 lvsat=7.101362528e-02 wvsat=1.454320924e-02 pvsat=-6.235387796e-9
+  ua=-3.057592724e-09 lua=5.811604481e-17 wua=2.139451025e-16 pua=-1.027429168e-22
+  ub=2.562876580e-18 lub=2.332695643e-25 wub=-7.631369240e-26 pub=5.922524027e-32
+  uc=1.850477845e-11 luc=1.430424627e-17 wuc=3.529147902e-17 puc=-1.316989093e-23
+  rdsw=484.7
+  prwb=0.1
+  prwg=0.052
+  wr=1.0
+  u0=7.031209847e-04 lu0=9.542676686e-10 wu0=1.703167720e-09 pu0=-6.815022648e-16
+  a0=1.1627
+  keta=-1.727325087e-02 lketa=2.065159494e-09 wketa=2.564480790e-09 pketa=-9.720664436e-16
+  a1=0.0
+  a2=0.46703705
+  ags=-6.872212874e-01 lags=3.650246752e-07 wags=8.693058230e-07 pags=-3.360774884e-13
+  b0=-2.221007410e-06 lb0=5.273470401e-13 wb0=5.480422528e-13 pb0=-5.968874215e-20
+  b1=2.306080819e-06 lb1=-7.471028750e-13 wb1=-9.268783038e-13 pb1=2.915465453e-19
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-6.393105e-11
+  cdsc=2.8125e-7
+  cdscb=1.0e-4
+  cdscd=1.0e-10
+  eta0=0.2
+  etab=-0.00025
+  dsub=1.0
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=0.030097
+  pdiblc1=0.0
+  pdiblc2=-1.109557813e-02 lpdiblc2=1.684004376e-08 wpdiblc2=-4.330260427e-08 ppdiblc2=3.694238737e-14
+  pdiblcb=-0.025
+  drout=0.43496
+  pscbe1=800000000.0
+  pscbe2=8.6797e-9
+  pvag=0.0
+  delta=1.482881207e-01 ldelta=-3.060677319e-08 wdelta=-5.658288556e-08 pdelta=1.600240242e-14
+  alpha0=5.0449517e-13
+  alpha1=-4.0583656e-18
+  beta0=6.2016506
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=2300000000.0
+  cgidl=0.5
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-7.880536625e-01 lkt1=6.479996892e-08 wkt1=1.129551183e-07 pkt1=-4.646606351e-14
+  kt2=1.626466176e-01 lkt2=-9.399894837e-08 wkt2=-1.167263343e-07 pkt2=4.424511700e-14
+  at=-2.555188328e+04 lat=2.375833456e-02 wat=1.658540408e-01 pat=-6.760303676e-8
+  ute=-7.869626397e-01 lute=2.178069211e-07 wute=4.569870802e-07 pute=-1.732209527e-13
+  ua1=1.972876075e-09 lua1=-4.737010877e-16 wua1=-5.882341500e-16 pua1=2.229701546e-22
+  ub1=-2.966932209e-18 lub1=1.036497900e-24 wub1=1.209925434e-24 pub1=-4.586222356e-31
+  uc1=-1.643084397e-10 luc1=7.365261409e-17 wuc1=9.146059397e-17 puc1=-3.466813815e-23
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+41
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=1.4472e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=1.0e-11
+  cgso=1.0e-11
+  cgbo=1.0e-13
+  capmod=2.0
+  xpart=0.0
+  cgsl=0.0
+  cgdl=0.0
+  cf=0.0
+  clc=7.0e-8
+  cle=0.492
+  dlc=-5.9781e-8
+  dwc=3.2175e-8
+  vfbcv=-1.0
+  acde=0.44
+  moin=8.7
+  noff=2.6123
+  voffcv=0.112
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000838062107
+  mjs=0.3362
+  pbs=0.6587
+  cjsws=9.9839168e-11
+  mjsws=0.2659
+  pbsws=0.7418
+  cjswgs=2.60659646e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.44e-6
+  sbref=1.44e-6
+  wlod={0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.40 pmos
* DC IV MOS Parameters
+  lmin=2.0e-05 lmax=1.0e-04 wmin=4.2e-07 wmax=5.5e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.4525e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=3.9651e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-7.916e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.44996e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.44996e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-5.583193162e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} wvth0=3.324507785e-8
+  k1=0.64774
+  k2=-7.830546258e-02 wk2=7.564334598e-9
+  k3=3.39
+  dvt0=2.4422
+  dvt1=0.16136
+  dvt2=0.026237
+  dvt0w=0.5
+  dvt1w=1928100.0
+  dvt2w=-0.032
+  w0=1.0e-8
+  k3b=1.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=123760.0
+  ua=-3.303158400e-09 wua=1.282926938e-16
+  ub=3.584115869e-18 wub=-2.386984254e-25
+  uc=5.990775477e-11 wuc=7.401501563e-20
+  rdsw=484.7
+  prwb=0.1
+  prwg=0.052
+  wr=1.0
+  u0=2.531468772e-03 wu0=-1.615377716e-11
+  a0=1.991478968e+00 wa0=-1.259488849e-7
+  keta=-0.01258
+  a1=0.0
+  a2=0.46703705
+  ags=5.586323740e-01 wags=-1.383957434e-7
+  b0=-4.838127228e-07 wb0=9.871135918e-14
+  b1=1.841100605e-07 wb1=5.464775321e-15
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-6.393105e-11
+  cdsc=2.8125e-7
+  cdscb=1.0e-4
+  cdscd=1.0e-10
+  eta0=0.2
+  etab=-0.00025
+  dsub=1.0
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-3.757870104e-01 wpclm=1.910487919e-7
+  pdiblc1=0.0
+  pdiblc2=1.219119946e-03 wpdiblc2=-3.700627423e-10
+  pdiblcb=-0.025
+  drout=4.577605585e-01 wdrout=-1.073217727e-8
+  pscbe1=800000000.0
+  pscbe2=8.6797e-9
+  pvag=0.0
+  delta=1.083269148e-02 wdelta=1.290328439e-9
+  alpha0=5.0449517e-13
+  alpha1=-4.0583656e-18
+  beta0=6.2016506
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=2300000000.0
+  cgidl=0.5
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-8.317952308e-01 wkt1=7.401501563e-8
+  kt2=-0.055045
+  at=2.613750069e+05 wat=9.806989571e-3
+  ute=-5.706649054e-01 wute=1.340288575e-7
+  ua1=6.8217e-10
+  ub1=-8.324836185e-20 wub1=-3.148105332e-26
+  uc1=-9.961e-12
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+41
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=1.4472e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=1.0e-11
+  cgso=1.0e-11
+  cgbo=1.0e-13
+  capmod=2.0
+  xpart=0.0
+  cgsl=0.0
+  cgdl=0.0
+  cf=0.0
+  clc=7.0e-8
+  cle=0.492
+  dlc=-5.9781e-8
+  dwc=3.2175e-8
+  vfbcv=-1.0
+  acde=0.44
+  moin=8.7
+  noff=2.6123
+  voffcv=0.112
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000838062107
+  mjs=0.3362
+  pbs=0.6587
+  cjsws=9.9839168e-11
+  mjsws=0.2659
+  pbsws=0.7418
+  cjswgs=2.60659646e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.41 pmos
* DC IV MOS Parameters
+  lmin=8e-06 lmax=2.0e-05 wmin=4.2e-07 wmax=5.5e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.4525e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=3.9651e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-7.916e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.44996e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.44996e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-6.345620892e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0=1.527070313e-06 wvth0=6.913239863e-08 pvth0=-7.187889422e-13
+  k1=0.64774
+  k2=-1.039190363e-01 lk2=5.130155488e-07 wk2=1.962059252e-08 pk2=-2.414753928e-13
+  k3=3.39
+  dvt0=2.4422
+  dvt1=0.16136
+  dvt2=0.026237
+  dvt0w=0.5
+  dvt1w=1928100.0
+  dvt2w=-0.032
+  w0=1.0e-8
+  k3b=1.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=123760.0
+  ua=-3.303158400e-09 wua=1.282926938e-16
+  ub=3.584115869e-18 wub=-2.386984254e-25
+  uc=5.990775477e-11 wuc=7.401501563e-20
+  rdsw=484.7
+  prwb=0.1
+  prwg=0.052
+  wr=1.0
+  u0=2.809795224e-03 lu0=-5.574614431e-09 wu0=-1.471614816e-10 pu0=2.623959863e-15
+  a0=1.695310514e+00 la0=5.931972766e-06 wa0=1.345701385e-08 pa0=-2.792167717e-12
+  keta=-0.01258
+  a1=0.0
+  a2=0.46703705
+  ags=5.586323740e-01 wags=-1.383957434e-7
+  b0=-4.901078367e-07 lb0=1.260851523e-13 wb0=1.016744567e-13 pb0=-5.934802904e-20
+  b1=1.973666236e-07 lb1=-2.655163654e-13 wb1=-7.750624224e-16 pb1=1.249780222e-19
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-6.393105e-11
+  cdsc=2.8125e-7
+  cdscb=1.0e-4
+  cdscd=1.0e-10
+  eta0=0.2
+  etab=-0.00025
+  dsub=1.0
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-3.757870104e-01 wpclm=1.910487919e-7
+  pdiblc1=0.0
+  pdiblc2=3.130572559e-03 lpdiblc2=-3.828457995e-08 wpdiblc2=-1.269779664e-09 ppdiblc2=1.802047521e-14
+  pdiblcb=-0.025
+  drout=4.577605585e-01 wdrout=-1.073217727e-8
+  pscbe1=800000000.0
+  pscbe2=8.6797e-9
+  pvag=0.0
+  delta=2.061905110e-02 ldelta=-1.960114861e-07 wdelta=-3.316091461e-09 pdelta=9.226221450e-14
+  alpha0=5.0449517e-13
+  alpha1=-4.0583656e-18
+  beta0=6.2016506
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=2300000000.0
+  cgidl=0.5
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-8.317952308e-01 wkt1=7.401501563e-8
+  kt2=-0.055045
+  at=2.325823130e+05 lat=5.766903068e-01 wat=2.335965303e-02 pat=-2.714469740e-7
+  ute=-5.706649054e-01 wute=1.340288575e-7
+  ua1=6.8217e-10
+  ub1=-3.849869378e-20 lub1=-8.962933392e-25 wub1=-5.254463258e-26 pub1=4.218834822e-31
+  uc1=-9.961e-12
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+41
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=1.4472e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=1.0e-11
+  cgso=1.0e-11
+  cgbo=1.0e-13
+  capmod=2.0
+  xpart=0.0
+  cgsl=0.0
+  cgdl=0.0
+  cf=0.0
+  clc=7.0e-8
+  cle=0.492
+  dlc=-5.9781e-8
+  dwc=3.2175e-8
+  vfbcv=-1.0
+  acde=0.44
+  moin=8.7
+  noff=2.6123
+  voffcv=0.112
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000838062107
+  mjs=0.3362
+  pbs=0.6587
+  cjsws=9.9839168e-11
+  mjsws=0.2659
+  pbsws=0.7418
+  cjswgs=2.60659646e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.42 pmos
* DC IV MOS Parameters
+  lmin=4e-06 lmax=8e-06 wmin=4.2e-07 wmax=5.5e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.4525e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=3.9651e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-7.916e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.44996e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.44996e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-3.847228985e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0=-4.789010406e-07 wvth0=-4.278175256e-08 pvth0=1.797753734e-13
+  k1=0.64774
+  k2=-5.815802816e-03 lk2=-2.746602181e-07 wk2=-2.192950090e-08 pk2=9.213238477e-14
+  k3=3.39
+  dvt0=2.4422
+  dvt1=0.16136
+  dvt2=0.026237
+  dvt0w=0.5
+  dvt1w=1928100.0
+  dvt2w=-0.032
+  w0=1.0e-8
+  k3b=1.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=123760.0
+  ua=-3.340967397e-09 lua=3.035703294e-16 wua=1.651962059e-16 pua=-2.963001438e-22
+  ub=3.871714484e-18 lub=-2.309143655e-24 wub=-3.886733045e-25 pub=1.204155803e-30
+  uc=9.549674441e-11 luc=-2.857457773e-16 wuc=-1.411457773e-17 puc=1.139209206e-22
+  rdsw=484.7
+  prwb=0.1
+  prwg=0.052
+  wr=1.0
+  u0=3.046000475e-03 lu0=-7.471118199e-09 wu0=-1.812372634e-10 pu0=2.897556019e-15
+  a0=2.738397109e+00 la0=-2.443021655e-06 wa0=-4.611647427e-07 pa0=1.018594097e-12
+  keta=-0.01258
+  a1=0.0
+  a2=0.46703705
+  ags=6.551333056e-01 lags=-7.748108052e-07 wags=-1.712734178e-07 pags=2.639764917e-13
+  b0=1.950206143e-07 lb0=-5.374845438e-12 wb0=-1.242555799e-13 pb0=1.754655532e-18
+  b1=1.769266582e-07 lb1=-1.014028617e-13 wb1=1.835676425e-14 pb1=-2.863237080e-20
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-6.393105e-11
+  cdsc=2.8125e-7
+  cdscb=1.0e-4
+  cdscd=1.0e-10
+  eta0=0.2
+  etab=-0.00025
+  dsub=1.0
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-3.757870104e-01 wpclm=1.910487919e-7
+  pdiblc1=0.0
+  pdiblc2=9.870057003e-04 lpdiblc2=-2.107377446e-08 wpdiblc2=-1.514456250e-09 ppdiblc2=1.998499576e-14
+  pdiblcb=-0.025
+  drout=4.577605585e-01 wdrout=-1.073217727e-8
+  pscbe1=800000000.0
+  pscbe2=8.6797e-9
+  pvag=0.0
+  delta=-1.998813163e-03 ldelta=-1.441152310e-08 wdelta=5.206524457e-09 pdelta=2.383370517e-14
+  alpha0=5.0449517e-13
+  alpha1=-4.0583656e-18
+  beta0=6.2016506
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=2300000000.0
+  cgidl=0.5
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-9.411865726e-01 lkt1=8.783085535e-07 wkt1=1.112912905e-07 pkt1=-2.992930745e-13
+  kt2=-0.055045
+  at=3.398108309e+05 lat=-2.842528254e-01 wat=-2.097278797e-02 pat=8.450041137e-8
+  ute=-1.049032909e+00 lute=3.840840622e-06 wute=2.690310995e-07 pute=-1.083939752e-12
+  ua1=6.681489060e-10 lua1=1.125760648e-16
+  ub1=-1.785851656e-19 lub1=2.284679476e-25
+  uc1=-9.961e-12
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+41
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=1.4472e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=1.0e-11
+  cgso=1.0e-11
+  cgbo=1.0e-13
+  capmod=2.0
+  xpart=0.0
+  cgsl=0.0
+  cgdl=0.0
+  cf=0.0
+  clc=7.0e-8
+  cle=0.492
+  dlc=-5.9781e-8
+  dwc=3.2175e-8
+  vfbcv=-1.0
+  acde=0.44
+  moin=8.7
+  noff=2.6123
+  voffcv=0.112
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000838062107
+  mjs=0.3362
+  pbs=0.6587
+  cjsws=9.9839168e-11
+  mjsws=0.2659
+  pbsws=0.7418
+  cjswgs=2.60659646e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.43 pmos
* DC IV MOS Parameters
+  lmin=2e-06 lmax=4e-06 wmin=4.2e-07 wmax=5.5e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.4525e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=3.9651e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-7.916e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.44996e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.44996e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-5.867775219e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0=3.351871395e-07 wvth0=3.159874274e-08 pvth0=-1.199073612e-13
+  k1=0.64774
+  k2=-9.497691035e-02 lk2=8.457434225e-08 wk2=8.053560467e-09 pk2=-2.867086861e-14
+  k3=3.39
+  dvt0=2.4422
+  dvt1=0.16136
+  dvt2=0.026237
+  dvt0w=0.5
+  dvt1w=1928100.0
+  dvt2w=-0.032
+  w0=1.0e-8
+  k3b=1.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=123760.0
+  ua=-3.228888558e-09 lua=-1.480009186e-16 wua=7.914024707e-17 pua=5.042361698e-23
+  ub=3.225123974e-18 lub=2.960018373e-25 wub=-6.477485772e-26 pub=-1.008472340e-31
+  uc=2.457536660e-11 wuc=1.416030607e-17
+  rdsw=484.7
+  prwb=0.1
+  prwg=0.052
+  wr=1.0
+  u0=9.411001758e-04 lu0=1.009630351e-09 wu0=6.458707932e-10 pu0=-4.349036964e-16
+  a0=1.952309073e+00 la0=7.241663461e-07 wa0=-1.237507747e-07 pa0=-3.408636508e-13
+  keta=-0.01258
+  a1=0.0
+  a2=0.46703705
+  ags=3.112859283e-01 lags=6.105674706e-07 wags=-7.309093508e-08 pags=-1.316056403e-13
+  b0=-1.782920227e-06 lb0=2.594377110e-12 wb0=5.370663884e-13 pb0=-9.098437448e-19
+  b1=1.625221979e-07 lb1=-4.336657078e-14 wb1=3.328278542e-15 pb1=3.191814955e-20
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-6.393105e-11
+  cdsc=2.8125e-7
+  cdscb=1.0e-4
+  cdscd=1.0e-10
+  eta0=0.2
+  etab=-0.00025
+  dsub=1.0
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-3.757870104e-01 wpclm=1.910487919e-7
+  pdiblc1=0.0
+  pdiblc2=-1.456551683e-02 lpdiblc2=4.158811642e-08 wpdiblc2=6.353757696e-09 ppdiblc2=-1.171643164e-14
+  pdiblcb=-0.025
+  drout=4.577605585e-01 wdrout=-1.073217727e-8
+  pscbe1=800000000.0
+  pscbe2=8.6797e-9
+  pvag=0.0
+  delta=-3.952571668e-02 ldelta=1.367862475e-07 wdelta=2.399868754e-08 pdelta=-5.188085951e-14
+  alpha0=5.0449517e-13
+  alpha1=-4.0583656e-18
+  beta0=6.2016506
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=2300000000.0
+  cgidl=0.5
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-6.844536037e-01 lkt1=-1.560814151e-07 wkt1=1.877313248e-08 pkt1=7.346720994e-14
+  kt2=-0.055045
+  at=3.069394585e+05 lat=-1.518124223e-1
+  ute=-1.364897622e-01 lute=1.641586551e-07 wute=1.917800739e-08 pute=-7.726915066e-14
+  ua1=6.9609e-10
+  ub1=-1.2188e-19
+  uc1=-9.961e-12
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+41
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=1.4472e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=1.0e-11
+  cgso=1.0e-11
+  cgbo=1.0e-13
+  capmod=2.0
+  xpart=0.0
+  cgsl=0.0
+  cgdl=0.0
+  cf=0.0
+  clc=7.0e-8
+  cle=0.492
+  dlc=-5.9781e-8
+  dwc=3.2175e-8
+  vfbcv=-1.0
+  acde=0.44
+  moin=8.7
+  noff=2.6123
+  voffcv=0.112
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000838062107
+  mjs=0.3362
+  pbs=0.6587
+  cjsws=9.9839168e-11
+  mjsws=0.2659
+  pbsws=0.7418
+  cjswgs=2.60659646e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.44 pmos
* DC IV MOS Parameters
+  lmin=1.5e-06 lmax=2e-06 wmin=4.2e-07 wmax=5.5e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.4525e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=3.9651e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-7.916e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.44996e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.44996e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-4.215833968e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} wvth0=-2.749657831e-8
+  k1=0.64774
+  k2=-5.329516655e-02 wk2=-6.076632783e-9
+  k3=3.39
+  dvt0=2.4422
+  dvt1=0.16136
+  dvt2=0.026237
+  dvt0w=0.5
+  dvt1w=1928100.0
+  dvt2w=-0.032
+  w0=1.0e-8
+  k3b=1.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=123760.0
+  ua=-3.301829549e-09 wua=1.039910970e-16
+  ub=3.371005957e-18 wub=-1.144765575e-25
+  uc=2.457536660e-11 wuc=1.416030607e-17
+  rdsw=484.7
+  prwb=0.1
+  prwg=0.052
+  wr=1.0
+  u0=1.438687890e-03 wu0=4.315322128e-10
+  a0=2.309208285e+00 wa0=-2.917425200e-7
+  keta=-0.01258
+  a1=0.0
+  a2=0.46703705
+  ags=6.121989026e-01 wags=-1.379516533e-7
+  b0=-5.043035789e-07 wb0=8.865765289e-14
+  b1=1.411493531e-07 wb1=1.905886653e-14
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-6.393105e-11
+  cdsc=2.8125e-7
+  cdscb=1.0e-4
+  cdscd=1.0e-10
+  eta0=0.2
+  etab=-0.00025
+  dsub=1.0
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-3.757870104e-01 wpclm=1.910487919e-7
+  pdiblc1=0.0
+  pdiblc2=5.930831918e-03 wpdiblc2=5.794142140e-10
+  pdiblcb=-0.025
+  drout=4.577605585e-01 wdrout=-1.073217727e-8
+  pscbe1=800000000.0
+  pscbe2=8.6797e-9
+  pvag=0.0
+  delta=2.788821965e-02 wdelta=-1.570351915e-9
+  alpha0=5.0449517e-13
+  alpha1=-4.0583656e-18
+  beta0=6.2016506
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=2300000000.0
+  cgidl=0.5
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-7.613769989e-01 wkt1=5.498082078e-8
+  kt2=-0.055045
+  at=232120.0
+  ute=-5.558556806e-02 wute=-1.890343499e-8
+  ua1=6.9609e-10
+  ub1=-1.2188e-19
+  uc1=-9.961e-12
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+41
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=1.4472e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=1.0e-11
+  cgso=1.0e-11
+  cgbo=1.0e-13
+  capmod=2.0
+  xpart=0.0
+  cgsl=0.0
+  cgdl=0.0
+  cf=0.0
+  clc=7.0e-8
+  cle=0.492
+  dlc=-5.9781e-8
+  dwc=3.2175e-8
+  vfbcv=-1.0
+  acde=0.44
+  moin=8.7
+  noff=2.6123
+  voffcv=0.112
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000838062107
+  mjs=0.3362
+  pbs=0.6587
+  cjsws=9.9839168e-11
+  mjsws=0.2659
+  pbsws=0.7418
+  cjswgs=2.60659646e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.45 pmos
* DC IV MOS Parameters
+  lmin=1e-06 lmax=1.5e-06 wmin=4.2e-07 wmax=5.5e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.4525e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=3.9651e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-7.916e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.44996e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.44996e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-4.108427007e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0=-1.642306134e-08 wvth0=-5.078635284e-09 pvth0=-3.427815578e-14
+  k1=0.64774
+  k2=-2.865391556e-02 lk2=-3.767770483e-08 wk2=1.077871532e-08 pk2=-2.577267001e-14
+  k3=3.39
+  dvt0=2.4422
+  dvt1=0.16136
+  dvt2=0.026237
+  dvt0w=0.5
+  dvt1w=1928100.0
+  dvt2w=-0.032
+  w0=1.0e-8
+  k3b=1.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=3.494623443e+05 lvsat=-3.451101695e-01 wvsat=-7.689633729e-02 pvsat=1.175783445e-7
+  ua=-4.405486298e-09 lua=1.687546352e-15 wua=3.205540120e-16 pua=-3.311355253e-22
+  ub=5.026345175e-18 lub=-2.531096431e-24 wub=-5.676592109e-25 pub=6.929389362e-31
+  uc=-6.585748721e-11 luc=1.382763551e-16 wuc=3.891651926e-17 puc=-3.785348777e-23
+  rdsw=484.7
+  prwb=0.1
+  prwg=0.052
+  wr=1.0
+  u0=5.546819766e-04 lu0=1.351689241e-09 wu0=9.356204573e-11 pu0=5.167732840e-16
+  a0=4.186371800e+00 la0=-2.870276874e-06 wa0=-8.160126484e-07 pa0=8.016352399e-13
+  keta=-1.820616449e-02 lketa=8.602686807e-09 wketa=1.916822988e-09 pketa=-2.930918190e-15
+  a1=0.0
+  a2=0.46703705
+  ags=-8.080961211e-01 lags=2.171702106e-06 wags=3.844143464e-07 pags=-7.987237318e-13
+  b0=-1.776643651e-06 lb0=1.945471588e-12 wb0=7.462853457e-13 pb0=-1.005545624e-18
+  b1=-5.982641671e-07 lb1=1.130600243e-12 wb1=5.869013386e-14 pb1=-6.059818932e-20
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-6.393105e-11
+  cdsc=2.8125e-7
+  cdscb=1.0e-4
+  cdscd=1.0e-10
+  eta0=0.2
+  etab=-0.00025
+  dsub=1.0
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-3.757870104e-01 wpclm=1.910487919e-7
+  pdiblc1=0.0
+  pdiblc2=-4.237301763e-02 lpdiblc2=7.385900115e-08 wpdiblc2=1.069592356e-08 ppdiblc2=-1.546864862e-14
+  pdiblcb=-0.025
+  drout=4.577605585e-01 wdrout=-1.073217727e-8
+  pscbe1=800000000.0
+  pscbe2=8.6797e-9
+  pvag=0.0
+  delta=1.769596352e-02 ldelta=1.558446922e-08 wdelta=-3.372927175e-09 pdelta=2.756227702e-15
+  alpha0=5.0449517e-13
+  alpha1=-4.0583656e-18
+  beta0=6.2016506
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=2300000000.0
+  cgidl=0.5
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-1.121349837e+00 lkt1=5.504164683e-07 wkt1=1.601141187e-07 pkt1=-1.607540692e-13
+  kt2=7.303081400e-03 lkt2=-9.533333386e-8
+  at=9.199711632e+05 lat=-1.051758821e+00 wat=-2.060775125e-01 pat=3.151028205e-7
+  ute=-1.691396183e-01 lute=1.736298206e-07 wute=3.866726444e-08 pute=-8.802847797e-14
+  ua1=4.063208202e-10 lua1=4.430715643e-16 wua1=1.101601979e-16 pua1=-1.684404507e-22
+  ub1=-4.225828834e-19 lub1=4.597897439e-25 wub1=1.144813009e-25 pub1=-1.750476331e-31
+  uc1=-9.220473410e-11 luc1=1.257547816e-16 puc1=5.877471754e-39
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+41
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=1.4472e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=1.0e-11
+  cgso=1.0e-11
+  cgbo=1.0e-13
+  capmod=2.0
+  xpart=0.0
+  cgsl=0.0
+  cgdl=0.0
+  cf=0.0
+  clc=7.0e-8
+  cle=0.492
+  dlc=-5.9781e-8
+  dwc=3.2175e-8
+  vfbcv=-1.0
+  acde=0.44
+  moin=8.7
+  noff=2.6123
+  voffcv=0.112
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000838062107
+  mjs=0.3362
+  pbs=0.6587
+  cjsws=9.9839168e-11
+  mjsws=0.2659
+  pbsws=0.7418
+  cjswgs=2.60659646e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=2.74e-6
+  sbref=2.74e-6
+  wlod={0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.46 pmos
* DC IV MOS Parameters
+  lmin=5e-07 lmax=1e-06 wmin=4.2e-07 wmax=5.5e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.4525e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=3.9651e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-7.916e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.44996e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.44996e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-1.881480639e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope2/sqrt(l*w*mult))} lvth0=-2.455869773e-07 wvth0=-1.222647949e-07 pvth0=8.631226181e-14
+  k1=0.64774
+  k2=-1.916237259e-02 lk2=-4.744497712e-08 wk2=-4.013784967e-08 pk2=2.662302118e-14
+  k3=3.39
+  dvt0=2.4422
+  dvt1=0.16136
+  dvt2=0.026237
+  dvt0w=0.5
+  dvt1w=1928100.0
+  dvt2w=-0.032
+  w0=1.0e-8
+  k3b=1.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=2.432375758e+04 lvsat=-1.052630688e-02 wvsat=2.359756276e-02 pvsat=1.416509669e-8
+  ua=-2.737560719e-09 lua=-2.883246528e-17 wua=5.410921996e-17 pua=-5.695051199e-23
+  ub=2.158046041e-18 lub=4.205267928e-25 wub=1.545346435e-25 pub=-5.023464973e-32
+  uc=8.789783820e-11 luc=-1.994556250e-17 wuc=-4.296747443e-18 puc=6.615124329e-24
+  rdsw=484.7
+  prwb=0.1
+  prwg=0.052
+  wr=1.0
+  u0=1.774797136e-05 lu0=1.904221179e-09 wu0=1.339924833e-09 pu0=-7.657963421e-16
+  a0=3.105714632e+00 la0=-1.758226614e-06 wa0=-7.636428554e-07 pa0=7.477441044e-13
+  keta=-9.846330846e-03 wketa=-9.313556134e-10
+  a1=0.0
+  a2=0.46703705
+  ags=1.187365417e+00 lags=1.182724101e-07 wags=-3.526038337e-07 pags=-4.029517358e-14
+  b0=1.085606693e-07 lb0=5.502081643e-15 wb0=-2.666991332e-13 pb0=3.686605431e-20
+  b1=1.255505918e-06 lb1=-7.770218633e-13 wb1=-1.541691454e-13 pb1=1.584446520e-19
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-6.393105e-11
+  cdsc=2.8125e-7
+  cdscb=1.0e-4
+  cdscd=1.0e-10
+  eta0=0.2
+  etab=-0.00025
+  dsub=1.0
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-7.143172486e-01 lpclm=3.483645416e-07 wpclm=3.503942980e-07 ppclm=-1.639744930e-13
+  pdiblc1=0.0
+  pdiblc2=-1.209408857e-01 lpdiblc2=1.547092658e-07 wpdiblc2=3.809126096e-08 ppdiblc2=-4.365982057e-14
+  pdiblcb=-0.025
+  drout=4.577605585e-01 wdrout=-1.073217727e-8
+  pscbe1=800000000.0
+  pscbe2=8.6797e-9
+  pvag=0.0
+  delta=8.733065673e-02 ldelta=-5.607311182e-08 wdelta=-2.789732286e-08 pdelta=2.799305709e-14
+  alpha0=5.0449517e-13
+  alpha1=-4.0583656e-18
+  beta0=6.2016506
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=2300000000.0
+  cgidl=0.5
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-4.653090187e-01 lkt1=-1.246823360e-07 wkt1=-3.619930332e-08 pkt1=4.126225775e-14
+  kt2=-0.085339
+  at=-2.433971696e+05 lat=1.454053617e-01 wat=1.718145740e-01 pat=-7.376703110e-8
+  ute=1.049633926e-01 lute=-1.084358829e-07 wute=-9.647585899e-08 pute=5.104055320e-14
+  ua1=8.769823734e-10 lua1=-4.126270701e-17 wua1=-7.239917656e-17 pua1=1.942227367e-23
+  ub1=8.150006008e-19 lub1=-8.137455405e-25 wub1=-3.356958845e-25 pub1=2.882071995e-31
+  uc1=3.0e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+41
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=1.4472e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=1.0e-11
+  cgso=1.0e-11
+  cgbo=1.0e-13
+  capmod=2.0
+  xpart=0.0
+  cgsl=0.0
+  cgdl=0.0
+  cf=0.0
+  clc=7.0e-8
+  cle=0.492
+  dlc=-5.9781e-8
+  dwc=3.2175e-8
+  vfbcv=-1.0
+  acde=0.44
+  moin=8.7
+  noff=2.6123
+  voffcv=0.112
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000838062107
+  mjs=0.3362
+  pbs=0.6587
+  cjsws=9.9839168e-11
+  mjsws=0.2659
+  pbsws=0.7418
+  cjswgs=2.60659646e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.74e-6
+  sbref=1.74e-6
+  wlod={0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.47 pmos
* DC IV MOS Parameters
+  lmin=3.5e-07 lmax=5e-07 wmin=4.2e-07 wmax=5.5e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=4.23e-9
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=-1.4525e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=3.9651e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-7.916e-9
+  dwb=0.0
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.69
+  rnoib=0.34
+  tnoia=25000000.0
+  tnoib=0.0
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={4.44996e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.44996e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope3/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={-5.587360718e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0=-4.952739170e-08 wvth0=-6.524946914e-08 pvth0=5.614830370e-14
+  k1=0.64774
+  k2=-1.045534012e-01 lk2=-2.268853432e-09 wk2=-1.085707761e-08 pk2=1.113202872e-14
+  k3=3.39
+  dvt0=2.4422
+  dvt1=0.16136
+  dvt2=0.026237
+  dvt0w=0.5
+  dvt1w=1928100.0
+  dvt2w=-0.032
+  w0=1.0e-8
+  k3b=1.0
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=-2.148436102e+05 lvsat=1.160051891e-01 wvsat=1.021873436e-01 pvsat=-2.741282688e-8
+  ua=-2.098588630e-09 lua=-3.668806491e-16 wua=-2.374562067e-16 pua=9.730217700e-23
+  ub=1.356266796e-18 lub=8.447081019e-25 wub=4.916351194e-25 pub=-2.285776565e-31
+  uc=8.475458580e-11 luc=-1.828262481e-17 wuc=4.107827200e-18 puc=2.168684114e-24
+  rdsw=484.7
+  prwb=0.1
+  prwg=0.052
+  wr=1.0
+  u0=4.628781384e-03 lu0=-5.352460477e-10 wu0=-1.446327791e-10 pu0=1.960886245e-17
+  a0=-2.176510508e-01 wa0=6.497284789e-7
+  keta=-9.846330846e-03 wketa=-9.313556134e-10
+  a1=0.0
+  a2=0.46703705
+  ags=3.799253448e+00 lags=-1.263546953e-06 wags=-1.242468862e-06 pags=4.304879197e-13
+  b0=4.195740248e-07 lb0=-1.590395341e-13 wb0=-6.948741474e-13 pb0=2.633920456e-19
+  b1=-7.519763816e-07 lb1=2.850366475e-13 wb1=5.125431043e-13 pb1=-1.942794637e-19
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-6.393105e-11
+  cdsc=2.8125e-7
+  cdscb=1.0e-4
+  cdscd=1.0e-10
+  eta0=0.2
+  etab=-0.00025
+  dsub=1.0
* BSIM4 - Sub-threshold parameters
+  voffl=0.0
+  minv=0.0
* Rout Parameters
+  pclm=-5.584538088e-02 wpclm=4.045290679e-8
+  pdiblc1=0.0
+  pdiblc2=-1.024427626e-01 lpdiblc2=1.449228338e-07 wpdiblc2=-3.056672116e-10 ppdiblc2=-2.334592572e-14
+  pdiblcb=-0.025
+  drout=4.577605585e-01 wdrout=-1.073217727e-8
+  pscbe1=800000000.0
+  pscbe2=8.6797e-9
+  pvag=0.0
+  delta=1.249699033e-01 ldelta=-7.598615521e-08 wdelta=-4.560704726e-08 pdelta=3.736238678e-14
+  alpha0=5.0449517e-13
+  alpha1=-4.0583656e-18
+  beta0=6.2016506
* BSIM4 - Rout Parameters
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=2300000000.0
+  cgidl=0.5
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=4.23e-9
* Temperature Effects Parameters
+  kt1=-8.612463619e-01 lkt1=8.478831547e-08 wkt1=1.474067755e-07 pkt1=-5.587453825e-14
+  kt2=-0.085339
+  at=8.416654710e+04 lat=-2.789222258e-02 wat=1.142097951e-01 pat=-4.329122282e-8
+  ute=1.839084500e-01 lute=-1.502017655e-7
+  ua1=9.905815277e-10 lua1=-1.013623396e-16 wua1=-1.258700713e-16 pua1=4.771105052e-23
+  ub1=-1.963011461e-18 lub1=6.559617409e-25 wub1=7.373819454e-25 pub1=-2.795046264e-31
+  uc1=3.0e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=3.0e+41
+  noib=0.0
+  noic=0.0
+  em=41000000.0
+  af=1.0
+  ef=0.88
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.3632
+  jss=2.1483e-5
+  jsws=1.4472e-10
+  xtis=5.2
+  bvs=12.69
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001671
+  tpbsw=0.001246
+  tpbswg=0.0
+  tcj=0.0012407
+  tcjsw=0.00037357
+  tcjswg=2.0e-12
+  cgdo=1.0e-11
+  cgso=1.0e-11
+  cgbo=1.0e-13
+  capmod=2.0
+  xpart=0.0
+  cgsl=0.0
+  cgdl=0.0
+  cf=0.0
+  clc=7.0e-8
+  cle=0.492
+  dlc=-5.9781e-8
+  dwc=3.2175e-8
+  vfbcv=-1.0
+  acde=0.44
+  moin=8.7
+  noff=2.6123
+  voffcv=0.112
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000838062107
+  mjs=0.3362
+  pbs=0.6587
+  cjsws=9.9839168e-11
+  mjsws=0.2659
+  pbsws=0.7418
+  cjswgs=2.60659646e-10
+  mjswgs=0.9274
+  pbswgs=1.4338
* Stress Parameters
+  saref=1.44e-6
+  sbref=1.44e-6
+  wlod={0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+  kvth0={0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+  lku0={0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+  wku0={0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.ends sky130_fd_pr__pfet_01v8_lvt
