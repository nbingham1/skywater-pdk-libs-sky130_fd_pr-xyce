* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param sky130_fd_pr__rf_nfet_g5v0d10v5__b_toxe_slope_spectre=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5__b_voff_slope_spectre=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5__b_nfactor_slope_spectre=0.0
* statistics {
*   process {
*   }
*   mismatch {
*     vary sky130_fd_pr__rf_nfet_g5v0d10v5__b_toxe_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__rf_nfet_g5v0d10v5__b_voff_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__rf_nfet_g5v0d10v5__b_nfactor_slope_spectre dist=gauss std = 1.0
*   }
* }
.subckt sky130_fd_pr__rf_nfet_g5v0d10v5_bM02 d g s b
.param l=1 w=1 ad=0 as=0 pd=0 ps=0 nrd=0 nrs=0 sa=0 sb=0 sd=0 mult=1 nf=1.0
msky130_fd_pr__rf_nfet_g5v0d10v5_bM02 d g s b sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__model l={l} w={w} ad={ad} as={as} pd={pd} ps={ps} nrd={nrd} nrs={nrs} sa={sa} sb={sb} sd={sd} nf={nf}
.model sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__model.0 nmos
* DC IV MOS Parameters
+  lmin=4.95E-07 lmax=5.05E-07 wmin=3.005E-06 wmax=3.015e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint={7.345E-08+sky130_fd_pr__rf_nfet_g5v0d10v5_b__lint_diff}
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint={2.135E-08+sky130_fd_pr__rf_nfet_g5v0d10v5_b__wint_diff}
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.129e-9
+  dwb=-1.694e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=3.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=1.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.5e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.16E-08*sky130_fd_pr__rf_nfet_g5v0d10v5_b__toxe_mult+sky130_fd_pr__rf_nfet_g5v0d10v5__b_toxe_slope_spectre*(1.16e-08*sky130_fd_pr__rf_nfet_g5v0d10v5_b__toxe_mult*(sky130_fd_pr__rf_nfet_g5v0d10v5__b_toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=6.0e+17
+  nsd=1.0e+20
+  rshg={49.2+sky130_fd_pr__rf_nfet_g5v0d10v5_b__rshg_diff}
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.8292+sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__vth0_diff_0}
+  k1=0.8833
+  k2={-0.03308+sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__k2_diff_0}
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.1925
+  dvt0w=0.16
+  dvt1w=6.909e+6
+  dvt2w=-0.03602
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat={1.0868E+05+sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__vsat_diff_0}
+  ua={1.663E-09+sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__ua_diff_0}
+  ub={1.238E-18+sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__ub_diff_0}
+  uc=6.62e-11
+  rdsw={724.6+sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__rdsw_diff_0}
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0={0.0636+sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__u0_diff_0}
+  a0={0.1745+sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__a0_diff_0}
+  keta=-0.01066
+  a1=0.0
+  a2=0.6597
+  ags={0+sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__ags_diff_0}
+  b0={3.293E-08+sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__b0_diff_0}
+  b1={0+sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__b1_diff_0}
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=370.0
+  rdwmin=0.0
+  rsw=370.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.2309+sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__voff_diff_0+sky130_fd_pr__rf_nfet_g5v0d10v5__b_voff_slope_spectre*(sky130_fd_pr__rf_nfet_g5v0d10v5__b_voff_slope/sqrt(l*w*mult))}
+  nfactor={0.627+sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__nfactor_diff_0+sky130_fd_pr__rf_nfet_g5v0d10v5__b_nfactor_slope_spectre*(sky130_fd_pr__rf_nfet_g5v0d10v5__b_nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-0.0008
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.05
+  etab=-0.01932
+  dsub=0.2822
* BSIM4 - Sub-threshold parameters
+  voffl=-4.258e-7
+  minv=0.0
* Rout Parameters
+  pclm={0.5653+sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__pclm_diff_0}
+  pdiblc1=0.211
+  pdiblc2=0.015
+  pdiblcb=-0.2683
+  drout=0.3896
+  pscbe1=9.373e+8
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.03542
+  alpha0=1.447e-5
+  alpha1=0.0
+  beta0=36.96
* BSIM4 - Rout Parameters
+  fprout=10.13
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1.058e+9
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1={-0.3307+sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__kt1_diff_0}
+  kt2=-0.01915
+  at=4.0e+4
+  ute=-1.299
+  ua1=3.604e-9
+  ub1=-3.553e-18
+  uc1=-5.982e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=10.0
+  xrcrg2=2.0
+  rbpb={200*sky130_fd_pr__rf_nfet_g5v0d10v5_b__rbpb_mult}
+  rbpd=200.0
+  rbps=200.0
+  rbdb=1.0e+5
+  rbsb=1.0e+5
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw={9E-07+sky130_fd_pr__rf_nfet_g5v0d10v5_b__xgw_diff}
+  xgl=0.0
+  ngcon=2.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.077
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.64
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.0009901
+  tpbswg=0.0
+  tcj=0.0006743
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo={2.7E-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult}
+  cgso={4.1E-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult}
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl={8E-11*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult}
+  cgdl={2.2E-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult}
+  cf=0.0
+  clc=1.0e-11
+  cle=0.6
+  dlc={1E-07+sky130_fd_pr__rf_nfet_g5v0d10v5_b__dlc_diff+sky130_fd_pr__rf_nfet_g5v0d10v5__base__dlc_rotweak}
+  dwc={0+sky130_fd_pr__rf_nfet_g5v0d10v5_b__dwc_diff}
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=2.0
+  voffcv=-0.1204
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs={0.001*sky130_fd_pr__rf_nfet_g5v0d10v5_b__ajunction_mult}
+  mjs=0.295
+  pbs=0.985
+  cjsws={4.864E-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__pjunction_mult}
+  mjsws=0.03759
+  pbsws=0.8907
+  cjswgs={3.948E-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__pjunction_mult}
+  mjswgs=0.1869
+  pbswgs=0.99
.ends sky130_fd_pr__rf_nfet_g5v0d10v5_bM02
.subckt sky130_fd_pr__rf_nfet_g5v0d10v5_bM02W5p00 d g s b
.param l=1 w=5.05 ad=0 as=0 pd=0 ps=0 nrd=0 nrs=0 sa=0 sb=0 sd=0 mult=1 nf=1.0
msky130_fd_pr__rf_nfet_g5v0d10v5_bM02W5p00 d g s b sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__model l={l} w=5.05 ad={ad} as={as} pd={pd} ps={ps} nrd={nrd} nrs={nrs} sa={sa} sb={sb} sd={sd} nf={nf}
.model sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__model.1 nmos
* DC IV MOS Parameters
+  lmin=4.95e-07 lmax=5.05E-07 wmin=4.995E-06 wmax=5.095e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint={7.345e-08+sky130_fd_pr__rf_nfet_g5v0d10v5_b__lint_diff}
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint={2.135e-08+sky130_fd_pr__rf_nfet_g5v0d10v5_b__wint_diff}
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.129e-9
+  dwb=-1.694e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=3.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=1.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.16e-08*sky130_fd_pr__rf_nfet_g5v0d10v5_b__toxe_mult+sky130_fd_pr__rf_nfet_g5v0d10v5__b_toxe_slope_spectre*(1.16e-08*sky130_fd_pr__rf_nfet_g5v0d10v5_b__toxe_mult*(sky130_fd_pr__rf_nfet_g5v0d10v5__b_toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=6.0e+17
+  nsd=1.0e+20
+  rshg={49.2+sky130_fd_pr__rf_nfet_g5v0d10v5_b__rshg_diff}
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.815+sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__vth0_diff_1}
+  k1=0.8833
+  k2={-0.03308+sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__k2_diff_1}
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.1925
+  dvt0w=0.16
+  dvt1w=6.909e+6
+  dvt2w=-0.03602
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat={1.035e+05+sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__vsat_diff_1}
+  ua={1.512e-09+sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__ua_diff_1}
+  ub={8.845e-19+sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__ub_diff_1}
+  uc=6.62e-11
+  rdsw={724.6+sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__rdsw_diff_1}
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0={0.0626+sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__u0_diff_1}
+  a0={0.1745+sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__a0_diff_1}
+  keta=-0.01066
+  a1=0.0
+  a2=0.6597
+  ags={0+sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__ags_diff_1}
+  b0={3.293e-08+sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__b0_diff_1}
+  b1={0+sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__b1_diff_1}
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=370.0
+  rdwmin=0.0
+  rsw=370.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.2309+sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__voff_diff_1+sky130_fd_pr__rf_nfet_g5v0d10v5__b_voff_slope_spectre*(sky130_fd_pr__rf_nfet_g5v0d10v5__b_voff_slope/sqrt(l*w*mult))}
+  nfactor={0.7788+sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__nfactor_diff_1+sky130_fd_pr__rf_nfet_g5v0d10v5__b_nfactor_slope_spectre*(sky130_fd_pr__rf_nfet_g5v0d10v5__b_nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-0.0008
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.05
+  etab=-0.01932
+  dsub=0.2822
* BSIM4 - Sub-threshold parameters
+  voffl=-4.258e-7
+  minv=0.0
* Rout Parameters
+  pclm={0.5653+sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__pclm_diff_1}
+  pdiblc1=0.211
+  pdiblc2=0.015
+  pdiblcb=-0.2683
+  drout=0.3896
+  pscbe1=9.373e+8
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.03542
+  alpha0=1.447e-5
+  alpha1=0.0
+  beta0=36.96
* BSIM4 - Rout Parameters
+  fprout=10.13
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1.058e+9
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1={-0.3507+sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__kt1_diff_1}
+  kt2=-0.01915
+  at=4.0e+4
+  ute=-1.299
+  ua1=3.004e-9
+  ub1=-3.553e-18
+  uc1=-5.982e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=10.0
+  xrcrg2=2.0
+  rbpb={140*sky130_fd_pr__rf_nfet_g5v0d10v5_b__rbpb_mult}
+  rbpd=140.0
+  rbps=140.0
+  rbdb=1.0e+5
+  rbsb=1.0e+5
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw={1.21e-06+sky130_fd_pr__rf_nfet_g5v0d10v5_b__xgw_diff}
+  xgl=0.0
+  ngcon=2.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.077
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.64
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.0009901
+  tpbswg=0.0
+  tcj=0.0006743
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo={2.2e-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult}
+  cgso={2.755e-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult}
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl={5e-11*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult}
+  cgdl={2e-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult}
+  cf=0.0
+  clc=1.0e-11
+  cle=0.6
+  dlc={5e-08+sky130_fd_pr__rf_nfet_g5v0d10v5_b__dlc_diff+sky130_fd_pr__rf_nfet_g5v0d10v5__base__dlc_rotweak}
+  dwc={0+sky130_fd_pr__rf_nfet_g5v0d10v5_b__dwc_diff}
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=2.0
+  voffcv=-0.1204
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs={0.001*sky130_fd_pr__rf_nfet_g5v0d10v5_b__ajunction_mult}
+  mjs=0.295
+  pbs=0.985
+  cjsws={4.864e-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__pjunction_mult}
+  mjsws=0.03759
+  pbsws=0.8907
+  cjswgs={3.748e-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__pjunction_mult}
+  mjswgs=0.1569
+  pbswgs=0.99
.ends sky130_fd_pr__rf_nfet_g5v0d10v5_bM02W5p00
.subckt sky130_fd_pr__rf_nfet_g5v0d10v5_bM04 d g s b
.param l=1 w=1 ad=0 as=0 pd=0 ps=0 nrd=0 nrs=0 sa=0 sb=0 sd=0 mult=1 nf=1.0
msky130_fd_pr__rf_nfet_g5v0d10v5_bM04 d g s b sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__model l={l} w={w} ad={ad} as={as} pd={pd} ps={ps} nrd={nrd} nrs={nrs} sa={sa} sb={sb} sd={sd} nf={nf}
.model sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__model.0 nmos
* DC IV MOS Parameters
+  lmin=4.95E-07 lmax=5.05E-07 wmin=3.005E-06 wmax=3.015e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint={7.345E-08+sky130_fd_pr__rf_nfet_g5v0d10v5_b__lint_diff}
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint={2.135E-08+sky130_fd_pr__rf_nfet_g5v0d10v5_b__wint_diff}
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.129e-9
+  dwb=-1.694e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=3.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=1.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.5e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.16E-08*sky130_fd_pr__rf_nfet_g5v0d10v5_b__toxe_mult+sky130_fd_pr__rf_nfet_g5v0d10v5__b_toxe_slope_spectre*(1.16e-08*sky130_fd_pr__rf_nfet_g5v0d10v5_b__toxe_mult*(sky130_fd_pr__rf_nfet_g5v0d10v5__b_toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=6.0e+17
+  nsd=1.0e+20
+  rshg={49.2+sky130_fd_pr__rf_nfet_g5v0d10v5_b__rshg_diff}
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.8372+sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__vth0_diff_0}
+  k1=0.8833
+  k2={-0.03308+sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__k2_diff_0}
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.1925
+  dvt0w=0.16
+  dvt1w=6.909e+6
+  dvt2w=-0.03602
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat={1.0868E+05+sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__vsat_diff_0}
+  ua={1.663E-09+sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__ua_diff_0}
+  ub={1.238E-18+sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__ub_diff_0}
+  uc=6.62e-11
+  rdsw={724.6+sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__rdsw_diff_0}
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0={0.0636+sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__u0_diff_0}
+  a0={0.1745+sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__a0_diff_0}
+  keta=-0.01066
+  a1=0.0
+  a2=0.6597
+  ags={0+sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__ags_diff_0}
+  b0={3.293E-08+sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__b0_diff_0}
+  b1={0+sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__b1_diff_0}
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=370.0
+  rdwmin=0.0
+  rsw=370.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.2309+sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__voff_diff_0+sky130_fd_pr__rf_nfet_g5v0d10v5__b_voff_slope_spectre*(sky130_fd_pr__rf_nfet_g5v0d10v5__b_voff_slope/sqrt(l*w*mult))}
+  nfactor={0.627+sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__nfactor_diff_0+sky130_fd_pr__rf_nfet_g5v0d10v5__b_nfactor_slope_spectre*(sky130_fd_pr__rf_nfet_g5v0d10v5__b_nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-0.0008
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.05
+  etab=-0.01932
+  dsub=0.2822
* BSIM4 - Sub-threshold parameters
+  voffl=-4.258e-7
+  minv=0.0
* Rout Parameters
+  pclm={0.5653+sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__pclm_diff_0}
+  pdiblc1=0.211
+  pdiblc2=0.015
+  pdiblcb=-0.2683
+  drout=0.3896
+  pscbe1=9.373e+8
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.03542
+  alpha0=1.447e-5
+  alpha1=0.0
+  beta0=36.96
* BSIM4 - Rout Parameters
+  fprout=10.13
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1.058e+9
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1={-0.3307+sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__kt1_diff_0}
+  kt2=-0.01915
+  at=4.0e+4
+  ute=-1.299
+  ua1=3.604e-9
+  ub1=-3.553e-18
+  uc1=-5.982e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=10.0
+  xrcrg2=2.0
+  rbpb={400*sky130_fd_pr__rf_nfet_g5v0d10v5_b__rbpb_mult}
+  rbpd=400.0
+  rbps=400.0
+  rbdb=1.0e+5
+  rbsb=1.0e+5
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw={1.25E-06+sky130_fd_pr__rf_nfet_g5v0d10v5_b__xgw_diff}
+  xgl=0.0
+  ngcon=2.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.077
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.64
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.0009901
+  tpbswg=0.0
+  tcj=0.0006743
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo={2.6E-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult}
+  cgso={3.7E-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult}
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl={5E-11*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult}
+  cgdl={2.1E-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult}
+  cf=0.0
+  clc=1.0e-11
+  cle=0.6
+  dlc={1E-07+sky130_fd_pr__rf_nfet_g5v0d10v5_b__dlc_diff+sky130_fd_pr__rf_nfet_g5v0d10v5__base__dlc_rotweak}
+  dwc={0+sky130_fd_pr__rf_nfet_g5v0d10v5_b__dwc_diff}
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=2.0
+  voffcv=-0.1204
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs={0.001*sky130_fd_pr__rf_nfet_g5v0d10v5_b__ajunction_mult}
+  mjs=0.295
+  pbs=0.985
+  cjsws={4.864E-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__pjunction_mult}
+  mjsws=0.03759
+  pbsws=0.8907
+  cjswgs={3.348E-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__pjunction_mult}
+  mjswgs=0.3069
+  pbswgs=0.99
.ends sky130_fd_pr__rf_nfet_g5v0d10v5_bM04
.subckt sky130_fd_pr__rf_nfet_g5v0d10v5_bM04W5p00 d g s b
.param l=1 w=5.05 ad=0 as=0 pd=0 ps=0 nrd=0 nrs=0 sa=0 sb=0 sd=0 mult=1 nf=1.0
msky130_fd_pr__rf_nfet_g5v0d10v5_bM04W5p00 d g s b sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__model l={l} w=5.05 ad={ad} as={as} pd={pd} ps={ps} nrd={nrd} nrs={nrs} sa={sa} sb={sb} sd={sd} nf={nf}
.model sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__model.1 nmos
* DC IV MOS Parameters
+  lmin=4.95e-07 lmax=5.05E-07 wmin=4.995E-06 wmax=5.095e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint={7.345e-08+sky130_fd_pr__rf_nfet_g5v0d10v5_b__lint_diff}
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint={2.135e-08+sky130_fd_pr__rf_nfet_g5v0d10v5_b__wint_diff}
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.129e-9
+  dwb=-1.694e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=3.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=1.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.16e-08*sky130_fd_pr__rf_nfet_g5v0d10v5_b__toxe_mult+sky130_fd_pr__rf_nfet_g5v0d10v5__b_toxe_slope_spectre*(1.16e-08*sky130_fd_pr__rf_nfet_g5v0d10v5_b__toxe_mult*(sky130_fd_pr__rf_nfet_g5v0d10v5__b_toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=6.0e+17
+  nsd=1.0e+20
+  rshg={49.2+sky130_fd_pr__rf_nfet_g5v0d10v5_b__rshg_diff}
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.815+sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__vth0_diff_1}
+  k1=0.8833
+  k2={-0.03308+sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__k2_diff_1}
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.1925
+  dvt0w=0.16
+  dvt1w=6.909e+6
+  dvt2w=-0.03602
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat={1.035e+05+sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__vsat_diff_1}
+  ua={1.512e-09+sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__ua_diff_1}
+  ub={8.845e-19+sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__ub_diff_1}
+  uc=6.62e-11
+  rdsw={724.6+sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__rdsw_diff_1}
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0={0.06175+sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__u0_diff_1}
+  a0={0.1745+sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__a0_diff_1}
+  keta=-0.01066
+  a1=0.0
+  a2=0.6597
+  ags={0+sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__ags_diff_1}
+  b0={3.293e-08+sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__b0_diff_1}
+  b1={0+sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__b1_diff_1}
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=370.0
+  rdwmin=0.0
+  rsw=370.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.2309+sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__voff_diff_1+sky130_fd_pr__rf_nfet_g5v0d10v5__b_voff_slope_spectre*(sky130_fd_pr__rf_nfet_g5v0d10v5__b_voff_slope/sqrt(l*w*mult))}
+  nfactor={0.6181+sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__nfactor_diff_1+sky130_fd_pr__rf_nfet_g5v0d10v5__b_nfactor_slope_spectre*(sky130_fd_pr__rf_nfet_g5v0d10v5__b_nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-0.0008
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.05
+  etab=-0.01932
+  dsub=0.2822
* BSIM4 - Sub-threshold parameters
+  voffl=-4.258e-7
+  minv=0.0
* Rout Parameters
+  pclm={0.5653+sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__pclm_diff_1}
+  pdiblc1=0.211
+  pdiblc2=0.015
+  pdiblcb=-0.2683
+  drout=0.3896
+  pscbe1=9.373e+8
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.03542
+  alpha0=1.447e-5
+  alpha1=0.0
+  beta0=36.96
* BSIM4 - Rout Parameters
+  fprout=10.13
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1.058e+9
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1={-0.3507+sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__kt1_diff_1}
+  kt2=-0.01915
+  at=4.0e+4
+  ute=-1.299
+  ua1=3.004e-9
+  ub1=-3.553e-18
+  uc1=-5.982e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=10.0
+  xrcrg2=2.0
+  rbpb={280*sky130_fd_pr__rf_nfet_g5v0d10v5_b__rbpb_mult}
+  rbpd=280.0
+  rbps=280.0
+  rbdb=1.0e+5
+  rbsb=1.0e+5
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw={9e-7+sky130_fd_pr__rf_nfet_g5v0d10v5_b__xgw_diff}
+  xgl=0.0
+  ngcon=2.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.077
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.64
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.0009901
+  tpbswg=0.0
+  tcj=0.0006743
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo={2.3e-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult}
+  cgso={3.755e-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult}
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl={5e-11*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult}
+  cgdl={2.2e-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult}
+  cf=0.0
+  clc=1.0e-11
+  cle=0.6
+  dlc={1.00e-07+sky130_fd_pr__rf_nfet_g5v0d10v5_b__dlc_diff+sky130_fd_pr__rf_nfet_g5v0d10v5__base__dlc_rotweak}
+  dwc={0+sky130_fd_pr__rf_nfet_g5v0d10v5_b__dwc_diff}
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=2.0
+  voffcv=-0.1204
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs={0.001*sky130_fd_pr__rf_nfet_g5v0d10v5_b__ajunction_mult}
+  mjs=0.295
+  pbs=0.985
+  cjsws={4.864e-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__pjunction_mult}
+  mjsws=0.03759
+  pbsws=0.8907
+  cjswgs={3.348e-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__pjunction_mult}
+  mjswgs=0.3069
+  pbswgs=0.99
.ends sky130_fd_pr__rf_nfet_g5v0d10v5_bM04W5p00
.subckt sky130_fd_pr__rf_nfet_g5v0d10v5_bM04W7p00 d g s b
.param l=1 w=7.09 ad=0 as=0 pd=0 ps=0 nrd=0 nrs=0 sa=0 sb=0 sd=0 mult=1 nf=1.0
msky130_fd_pr__rf_nfet_g5v0d10v5_bM04W7p00 d g s b sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__model l={l} w=7.09 ad={ad} as={as} pd={pd} ps={ps} nrd={nrd} nrs={nrs} sa={sa} sb={sb} sd={sd} nf={nf}
.model sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__model.2 nmos
* DC IV MOS Parameters
+  lmin=4.95E-07 lmax=5.05E-07 wmin=7.085E-06 wmax=7.095e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint={7.345E-08+sky130_fd_pr__rf_nfet_g5v0d10v5_b__lint_diff}
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint={2.135E-08+sky130_fd_pr__rf_nfet_g5v0d10v5_b__wint_diff}
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.129e-9
+  dwb=-1.694e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=3.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=1.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.5e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.16E-08*sky130_fd_pr__rf_nfet_g5v0d10v5_b__toxe_mult+sky130_fd_pr__rf_nfet_g5v0d10v5__b_toxe_slope_spectre*(1.16e-08*sky130_fd_pr__rf_nfet_g5v0d10v5_b__toxe_mult*(sky130_fd_pr__rf_nfet_g5v0d10v5__b_toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=6.0e+17
+  nsd=1.0e+20
+  rshg={49.2+sky130_fd_pr__rf_nfet_g5v0d10v5_b__rshg_diff}
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.811+sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__vth0_diff_2}
+  k1=0.8833
+  k2={-0.03308+sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__k2_diff_2}
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.1925
+  dvt0w=0.16
+  dvt1w=6.909e+6
+  dvt2w=-0.03602
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat={1.056E+05+sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__vsat_diff_2}
+  ua={1.588E-09+sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__ua_diff_2}
+  ub={8.757E-19+sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__ub_diff_2}
+  uc=6.62e-11
+  rdsw={724.6+sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__rdsw_diff_2}
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0={0.06298+sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__u0_diff_2}
+  a0={0.1745+sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__a0_diff_2}
+  keta=-0.01066
+  a1=0.0
+  a2=0.6597
+  ags={0+sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__ags_diff_2}
+  b0={3.293E-08+sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__b0_diff_2}
+  b1={0+sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__b1_diff_2}
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=370.0
+  rdwmin=0.0
+  rsw=370.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.2309+sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__voff_diff_2+sky130_fd_pr__rf_nfet_g5v0d10v5__b_voff_slope_spectre*(sky130_fd_pr__rf_nfet_g5v0d10v5__b_voff_slope/sqrt(l*w*mult))}
+  nfactor={0.7232+sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__nfactor_diff_2+sky130_fd_pr__rf_nfet_g5v0d10v5__b_nfactor_slope_spectre*(sky130_fd_pr__rf_nfet_g5v0d10v5__b_nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-0.0008
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.05
+  etab=-0.01932
+  dsub=0.2822
* BSIM4 - Sub-threshold parameters
+  voffl=-4.258e-7
+  minv=0.0
* Rout Parameters
+  pclm={0.5653+sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__pclm_diff_2}
+  pdiblc1=0.211
+  pdiblc2=0.015
+  pdiblcb=-0.2683
+  drout=0.3896
+  pscbe1=9.373e+8
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.03542
+  alpha0=1.447e-5
+  alpha1=0.0
+  beta0=36.96
* BSIM4 - Rout Parameters
+  fprout=10.13
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1.058e+9
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1={-0.3507+sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__kt1_diff_2}
+  kt2=-0.01915
+  at=4.0e+4
+  ute=-1.299
+  ua1=3.004e-9
+  ub1=-3.553e-18
+  uc1=-5.982e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=10.0
+  xrcrg2=2.0
+  rbpb={220*sky130_fd_pr__rf_nfet_g5v0d10v5_b__rbpb_mult}
+  rbpd=220.0
+  rbps=220.0
+  rbdb=1.0e+5
+  rbsb=1.0e+5
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw={1.5E-06+sky130_fd_pr__rf_nfet_g5v0d10v5_b__xgw_diff}
+  xgl=0.0
+  ngcon=2.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.077
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.64
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.0009901
+  tpbswg=0.0
+  tcj=0.0006743
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo={2.3E-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult}
+  cgso={3.2E-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult}
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl={5E-11*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult}
+  cgdl={2E-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult}
+  cf=0.0
+  clc=1.0e-11
+  cle=0.6
+  dlc={1E-07+sky130_fd_pr__rf_nfet_g5v0d10v5_b__dlc_diff+sky130_fd_pr__rf_nfet_g5v0d10v5__base__dlc_rotweak}
+  dwc={0+sky130_fd_pr__rf_nfet_g5v0d10v5_b__dwc_diff}
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=2.0
+  voffcv=-0.1204
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs={0.001*sky130_fd_pr__rf_nfet_g5v0d10v5_b__ajunction_mult}
+  mjs=0.295
+  pbs=0.985
+  cjsws={4.864E-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__pjunction_mult}
+  mjsws=0.03759
+  pbsws=0.8907
+  cjswgs={3.348E-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__pjunction_mult}
+  mjswgs=0.3069
+  pbswgs=0.99
.ends sky130_fd_pr__rf_nfet_g5v0d10v5_bM04W7p00
.subckt sky130_fd_pr__rf_nfet_g5v0d10v5_bM10 d g s b
.param l=1 w=1 ad=0 as=0 pd=0 ps=0 nrd=0 nrs=0 sa=0 sb=0 sd=0 mult=1 nf=1.0
msky130_fd_pr__rf_nfet_g5v0d10v5_bM10 d g s b sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__model l={l} w={w} ad={ad} as={as} pd={pd} ps={ps} nrd={nrd} nrs={nrs} sa={sa} sb={sb} sd={sd} nf={nf}
.model sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__model.0 nmos
* DC IV MOS Parameters
+  lmin=4.95E-07 lmax=5.05E-07 wmin=3.005E-06 wmax=3.015e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint={7.345E-08+sky130_fd_pr__rf_nfet_g5v0d10v5_b__lint_diff}
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint={2.135E-08+sky130_fd_pr__rf_nfet_g5v0d10v5_b__wint_diff}
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.129e-9
+  dwb=-1.694e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=3.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=1.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.5e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.16E-08*sky130_fd_pr__rf_nfet_g5v0d10v5_b__toxe_mult+sky130_fd_pr__rf_nfet_g5v0d10v5__b_toxe_slope_spectre*(1.16e-08*sky130_fd_pr__rf_nfet_g5v0d10v5_b__toxe_mult*(sky130_fd_pr__rf_nfet_g5v0d10v5__b_toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=6.0e+17
+  nsd=1.0e+20
+  rshg={49.2+sky130_fd_pr__rf_nfet_g5v0d10v5_b__rshg_diff}
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.8292+sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__vth0_diff_0}
+  k1=0.8833
+  k2={-0.03308+sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__k2_diff_0}
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.1925
+  dvt0w=0.16
+  dvt1w=6.909e+6
+  dvt2w=-0.03602
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat={1.0868E+05+sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__vsat_diff_0}
+  ua={1.663E-09+sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__ua_diff_0}
+  ub={1.238E-18+sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__ub_diff_0}
+  uc=6.62e-11
+  rdsw={724.6+sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__rdsw_diff_0}
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0={0.06175+sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__u0_diff_0}
+  a0={0.1745+sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__a0_diff_0}
+  keta=-0.01066
+  a1=0.0
+  a2=0.6597
+  ags={0+sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__ags_diff_0}
+  b0={3.293E-08+sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__b0_diff_0}
+  b1={0+sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__b1_diff_0}
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=370.0
+  rdwmin=0.0
+  rsw=370.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.2309+sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__voff_diff_0+sky130_fd_pr__rf_nfet_g5v0d10v5__b_voff_slope_spectre*(sky130_fd_pr__rf_nfet_g5v0d10v5__b_voff_slope/sqrt(l*w*mult))}
+  nfactor={0.7376+sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__nfactor_diff_0+sky130_fd_pr__rf_nfet_g5v0d10v5__b_nfactor_slope_spectre*(sky130_fd_pr__rf_nfet_g5v0d10v5__b_nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-0.0008
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.05
+  etab=-0.01932
+  dsub=0.2822
* BSIM4 - Sub-threshold parameters
+  voffl=-4.258e-7
+  minv=0.0
* Rout Parameters
+  pclm={0.5653+sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__pclm_diff_0}
+  pdiblc1=0.211
+  pdiblc2=0.015
+  pdiblcb=-0.2683
+  drout=0.3896
+  pscbe1=9.373e+8
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.03542
+  alpha0=1.447e-5
+  alpha1=0.0
+  beta0=36.96
* BSIM4 - Rout Parameters
+  fprout=10.13
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1.058e+9
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1={-0.3307+sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__kt1_diff_0}
+  kt2=-0.01915
+  at=4.0e+4
+  ute=-1.299
+  ua1=3.604e-9
+  ub1=-3.553e-18
+  uc1=-5.982e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=10.0
+  xrcrg2=2.0
+  rbpb={1000*sky130_fd_pr__rf_nfet_g5v0d10v5_b__rbpb_mult}
+  rbpd=1000.0
+  rbps=1000.0
+  rbdb=1.0e+5
+  rbsb=1.0e+5
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw={1.25E-06+sky130_fd_pr__rf_nfet_g5v0d10v5_b__xgw_diff}
+  xgl=0.0
+  ngcon=2.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.077
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.64
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.0009901
+  tpbswg=0.0
+  tcj=0.0006743
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo={2.7E-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult}
+  cgso={3.7E-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult}
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl={5E-11*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult}
+  cgdl={2.2E-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult}
+  cf=0.0
+  clc=1.0e-11
+  cle=0.6
+  dlc={1E-07+sky130_fd_pr__rf_nfet_g5v0d10v5_b__dlc_diff+sky130_fd_pr__rf_nfet_g5v0d10v5__base__dlc_rotweak}
+  dwc={0+sky130_fd_pr__rf_nfet_g5v0d10v5_b__dwc_diff}
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=2.0
+  voffcv=-0.1204
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs={0.001*sky130_fd_pr__rf_nfet_g5v0d10v5_b__ajunction_mult}
+  mjs=0.295
+  pbs=0.985
+  cjsws={4.864E-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__pjunction_mult}
+  mjsws=0.03759
+  pbsws=0.8907
+  cjswgs={3.048E-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__pjunction_mult}
+  mjswgs=0.2969
+  pbswgs=0.99
.ends sky130_fd_pr__rf_nfet_g5v0d10v5_bM10
.subckt sky130_fd_pr__rf_nfet_g5v0d10v5_bM10W5p00 d g s b
.param l=1 w=5.05 ad=0 as=0 pd=0 ps=0 nrd=0 nrs=0 sa=0 sb=0 sd=0 mult=1 nf=1.0
msky130_fd_pr__rf_nfet_g5v0d10v5_bM10W5p00 d g s b sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__model l={l} w=5.05 ad={ad} as={as} pd={pd} ps={ps} nrd={nrd} nrs={nrs} sa={sa} sb={sb} sd={sd} nf={nf}
.model sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__model.1 nmos
* DC IV MOS Parameters
+  lmin=4.95E-07 lmax=5.05E-07 wmin=5.045E-06 wmax=5.055e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint={7.345E-08+sky130_fd_pr__rf_nfet_g5v0d10v5_b__lint_diff}
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint={2.135E-08+sky130_fd_pr__rf_nfet_g5v0d10v5_b__wint_diff}
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.129e-9
+  dwb=-1.694e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=3.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=1.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.5e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.16E-08*sky130_fd_pr__rf_nfet_g5v0d10v5_b__toxe_mult+sky130_fd_pr__rf_nfet_g5v0d10v5__b_toxe_slope_spectre*(1.16e-08*sky130_fd_pr__rf_nfet_g5v0d10v5_b__toxe_mult*(sky130_fd_pr__rf_nfet_g5v0d10v5__b_toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=6.0e+17
+  nsd=1.0e+20
+  rshg={49.2+sky130_fd_pr__rf_nfet_g5v0d10v5_b__rshg_diff}
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.815+sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__vth0_diff_1}
+  k1=0.8833
+  k2={-0.03308+sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__k2_diff_1}
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.1925
+  dvt0w=0.16
+  dvt1w=6.909e+6
+  dvt2w=-0.03602
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat={1.056E+05+sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__vsat_diff_1}
+  ua={1.724E-09+sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__ua_diff_1}
+  ub={1.624E-18+sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__ub_diff_1}
+  uc=6.62e-11
+  rdsw={724.6+sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__rdsw_diff_1}
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0={0.06545+sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__u0_diff_1}
+  a0={0.1745+sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__a0_diff_1}
+  keta=-0.01066
+  a1=0.0
+  a2=0.6597
+  ags={0+sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__ags_diff_1}
+  b0={3.293E-08+sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__b0_diff_1}
+  b1={0+sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__b1_diff_1}
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=370.0
+  rdwmin=0.0
+  rsw=370.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.2309+sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__voff_diff_1+sky130_fd_pr__rf_nfet_g5v0d10v5__b_voff_slope_spectre*(sky130_fd_pr__rf_nfet_g5v0d10v5__b_voff_slope/sqrt(l*w*mult))}
+  nfactor={0.7664+sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__nfactor_diff_1+sky130_fd_pr__rf_nfet_g5v0d10v5__b_nfactor_slope_spectre*(sky130_fd_pr__rf_nfet_g5v0d10v5__b_nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-0.0008
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.05
+  etab=-0.01932
+  dsub=0.2822
* BSIM4 - Sub-threshold parameters
+  voffl=-4.258e-7
+  minv=0.0
* Rout Parameters
+  pclm={0.5653+sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__pclm_diff_1}
+  pdiblc1=0.211
+  pdiblc2=0.015
+  pdiblcb=-0.2683
+  drout=0.3896
+  pscbe1=9.373e+8
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.03542
+  alpha0=1.447e-5
+  alpha1=0.0
+  beta0=36.96
* BSIM4 - Rout Parameters
+  fprout=10.13
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1.058e+9
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1={-0.3207+sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__kt1_diff_1}
+  kt2=-0.01915
+  at=4.0e+4
+  ute=-1.377
+  ua1=3.094e-9
+  ub1=-1.812e-18
+  uc1=-5.982e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=10.0
+  xrcrg2=2.0
+  rbpb={700*sky130_fd_pr__rf_nfet_g5v0d10v5_b__rbpb_mult}
+  rbpd=700.0
+  rbps=700.0
+  rbdb=1.0e+5
+  rbsb=1.0e+5
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw={1.25E-06+sky130_fd_pr__rf_nfet_g5v0d10v5_b__xgw_diff}
+  xgl=0.0
+  ngcon=2.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.077
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.64
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.0009901
+  tpbswg=0.0
+  tcj=0.0006743
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo={2.3E-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult}
+  cgso={3.6E-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult}
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl={5E-11*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult}
+  cgdl={2E-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult}
+  cf=0.0
+  clc=1.0e-11
+  cle=0.6
+  dlc={1E-07+sky130_fd_pr__rf_nfet_g5v0d10v5_b__dlc_diff+sky130_fd_pr__rf_nfet_g5v0d10v5__base__dlc_rotweak}
+  dwc={0+sky130_fd_pr__rf_nfet_g5v0d10v5_b__dwc_diff}
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=2.0
+  voffcv=-0.1204
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs={0.001*sky130_fd_pr__rf_nfet_g5v0d10v5_b__ajunction_mult}
+  mjs=0.295
+  pbs=0.985
+  cjsws={4.864E-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__pjunction_mult}
+  mjsws=0.03759
+  pbsws=0.8907
+  cjswgs={2.848E-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__pjunction_mult}
+  mjswgs=0.3069
+  pbswgs=0.99
.ends sky130_fd_pr__rf_nfet_g5v0d10v5_bM10W5p00
.subckt sky130_fd_pr__rf_nfet_g5v0d10v5_bM10W7p00 d g s b
.param l=1 w=7.09 ad=0 as=0 pd=0 ps=0 nrd=0 nrs=0 sa=0 sb=0 sd=0 mult=1 nf=1.0
msky130_fd_pr__rf_nfet_g5v0d10v5_bM10W7p00 d g s b sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__model l={l} w=7.09 ad={ad} as={as} pd={pd} ps={ps} nrd={nrd} nrs={nrs} sa={sa} sb={sb} sd={sd} nf={nf}
.model sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__model.2 nmos
* DC IV MOS Parameters
+  lmin=4.95E-07 lmax=5.05E-07 wmin=7.085E-06 wmax=7.095e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint={7.345E-08+sky130_fd_pr__rf_nfet_g5v0d10v5_b__lint_diff}
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint={2.135E-08+sky130_fd_pr__rf_nfet_g5v0d10v5_b__wint_diff}
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.129e-9
+  dwb=-1.694e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=3.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=1.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.5e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.16E-08*sky130_fd_pr__rf_nfet_g5v0d10v5_b__toxe_mult+sky130_fd_pr__rf_nfet_g5v0d10v5__b_toxe_slope_spectre*(1.16e-08*sky130_fd_pr__rf_nfet_g5v0d10v5_b__toxe_mult*(sky130_fd_pr__rf_nfet_g5v0d10v5__b_toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=6.0e+17
+  nsd=1.0e+20
+  rshg={49.2+sky130_fd_pr__rf_nfet_g5v0d10v5_b__rshg_diff}
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.811+sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__vth0_diff_2}
+  k1=0.8833
+  k2={-0.03308+sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__k2_diff_2}
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.1925
+  dvt0w=0.16
+  dvt1w=6.909e+6
+  dvt2w=-0.03602
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat={1.056E+05+sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__vsat_diff_2}
+  ua={1.89E-09+sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__ua_diff_2}
+  ub={1.437E-18+sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__ub_diff_2}
+  uc=6.62e-11
+  rdsw={724.6+sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__rdsw_diff_2}
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0={0.0655+sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__u0_diff_2}
+  a0={0.1745+sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__a0_diff_2}
+  keta=-0.01066
+  a1=0.0
+  a2=0.6597
+  ags={0+sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__ags_diff_2}
+  b0={3.293E-08+sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__b0_diff_2}
+  b1={0+sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__b1_diff_2}
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=370.0
+  rdwmin=0.0
+  rsw=370.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.2309+sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__voff_diff_2+sky130_fd_pr__rf_nfet_g5v0d10v5__b_voff_slope_spectre*(sky130_fd_pr__rf_nfet_g5v0d10v5__b_voff_slope/sqrt(l*w*mult))}
+  nfactor={0.687+sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__nfactor_diff_2+sky130_fd_pr__rf_nfet_g5v0d10v5__b_nfactor_slope_spectre*(sky130_fd_pr__rf_nfet_g5v0d10v5__b_nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-0.0008
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.05
+  etab=-0.01932
+  dsub=0.2822
* BSIM4 - Sub-threshold parameters
+  voffl=-4.258e-7
+  minv=0.0
* Rout Parameters
+  pclm={0.5653+sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__pclm_diff_2}
+  pdiblc1=0.211
+  pdiblc2=0.015
+  pdiblcb=-0.2683
+  drout=0.3896
+  pscbe1=9.373e+8
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.03542
+  alpha0=1.447e-5
+  alpha1=0.0
+  beta0=36.96
* BSIM4 - Rout Parameters
+  fprout=10.13
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1.058e+9
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1={-0.3507+sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__kt1_diff_2}
+  kt2=-0.01915
+  at=4.0e+4
+  ute=-1.299
+  ua1=3.004e-9
+  ub1=-3.553e-18
+  uc1=-5.982e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=10.0
+  xrcrg2=2.0
+  rbpb={550*sky130_fd_pr__rf_nfet_g5v0d10v5_b__rbpb_mult}
+  rbpd=550.0
+  rbps=550.0
+  rbdb=1.0e+5
+  rbsb=1.0e+5
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw={1.5E-06+sky130_fd_pr__rf_nfet_g5v0d10v5_b__xgw_diff}
+  xgl=0.0
+  ngcon=2.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.077
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.64
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.0009901
+  tpbswg=0.0
+  tcj=0.0006743
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo={2.3E-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult}
+  cgso={3.4E-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult}
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl={5E-11*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult}
+  cgdl={1.8E-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult}
+  cf=0.0
+  clc=1.0e-11
+  cle=0.6
+  dlc={1E-07+sky130_fd_pr__rf_nfet_g5v0d10v5_b__dlc_diff+sky130_fd_pr__rf_nfet_g5v0d10v5__base__dlc_rotweak}
+  dwc={0+sky130_fd_pr__rf_nfet_g5v0d10v5_b__dwc_diff}
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=2.0
+  voffcv=-0.1204
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs={0.001*sky130_fd_pr__rf_nfet_g5v0d10v5_b__ajunction_mult}
+  mjs=0.295
+  pbs=0.985
+  cjsws={4.864E-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__pjunction_mult}
+  mjsws=0.03759
+  pbsws=0.8907
+  cjswgs={2.748E-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__pjunction_mult}
+  mjswgs=0.3069
+  pbswgs=0.99
.ends sky130_fd_pr__rf_nfet_g5v0d10v5_bM10W7p00
