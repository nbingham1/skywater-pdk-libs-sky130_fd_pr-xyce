* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param
+  sky130_fd_pr__nfet_01v8_lvt__ajunction_mult=8.7784e-1
+  sky130_fd_pr__nfet_01v8_lvt__pjunction_mult=7.8244e-1
.include "sky130_fd_pr__nfet_01v8_lvt__ff.pm3.spice"
