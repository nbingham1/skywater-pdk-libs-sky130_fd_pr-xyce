* SKY130 Spice File.
*  P+ Poly Preres Corner Parameters
.param
+  sky130_fd_pr__res_high_po__var_mult=-5.0
+  sky130_fd_pr__res_high_po__var=-0.125
+  sky130_fd_pr__res_xhigh_po__var_mult=-0.15
+  camimc=2.231e-15 ; Units: farad/micrometer^2
+  cpmimc=0.35e-15 ; Units: farad/micrometer
+  cvpp_cor=1.136
+  cvpp3_cor=1.3
+  cvpp4_cor=1.3
+  cvpp5_cor=1.3
+  cm3m2_vpp=1.620
+  c0m5m4_vpp=1.487
+  c1m5m4_vpp=1.419
+  c0m5m4_vpp0p4shield=3.04132
+  c1m5m4_vpp0p4shield=1.50414
+  c0m4m3_vpp=1.487
+  c1m4m3_vpp=1.419
+  c0m5m3_vpp=1.366
+  c1m5m3_vpp=1.496
+  cpl2s_vpp=1.460
+  cpl2s_vpp0p4shield=1.5250
+  cli2s_vpp=1.347
+  sky130_fd_pr__cap_vpp_08p6x07p8_m1m2m3_shieldl1__cor=1.190
+  sky130_fd_pr__cap_vpp_04p4x04p6_m1m2m3_shieldl1__cor=1.225
+  sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3_shieldl1__cor=1.145
+  sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_noshield__cor=1.173
+  sky130_fd_pr__cap_vpp_04p4x04p6_l1m1m2_noshield__cor=1.204
+  sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2_noshield__cor=1.132
+  sky130_fd_pr__cap_vpp_01p8x01p8_m1m2_noshield__cor=1.214
+  sky130_fd_pr__cap_vpp_08p6x07p8_m1m2_shieldl1__cor=1.173
+  sky130_fd_pr__cap_vpp_04p4x04p6_m1m2_shieldl1__cor=1.204
+  sky130_fd_pr__cap_vpp_11p5x11p7_m1m2_shieldl1__cor=1.132
+  sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_shieldpo_floatm3__cor=1.154
+  sky130_fd_pr__cap_vpp_04p4x04p6_l1m1m2_shieldpo_floatm3__cor=1.184
+  sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2_shieldpom3__cor=1.115
+  sky130_fd_pr__cap_vpp_03p9x03p9_m1m2_shieldl1_floatm3__cor=1.123
+  sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3m4_shieldm5__cor=1.144
+  sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3m4_shieldpom5__cor=1.144
+  sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3m4_shieldl1m5__cor=1.144
+  sky130_fd_pr__cap_vpp_08p6x07p8_m1m2m3_shieldl1m5_floatm4__cor=1.208
+  sky130_fd_pr__cap_vpp_06p8x06p1_l1m1m2_noshield__cor=1.2
+  sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3_shieldm4__cor=1.2
+  sky130_fd_pr__model__cap_vpp_finger__cor=1.2
+  sky130_fd_pr__cap_vpp_11p5x11p7_pol1m1m2m3m4m5_noshield_base__cor=1.2
*.param cm3m2_vpp = 1.362
