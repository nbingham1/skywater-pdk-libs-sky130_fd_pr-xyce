* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 68
.param
+  sky130_fd_pr__pfet_01v8_hvt__toxe_mult=1.0
+  sky130_fd_pr__pfet_01v8_hvt__rshp_mult=1.0
+  sky130_fd_pr__pfet_01v8_hvt__overlap_mult=0.98867
+  sky130_fd_pr__pfet_01v8_hvt__lint_diff=0.0
+  sky130_fd_pr__pfet_01v8_hvt__wint_diff=0.0
+  sky130_fd_pr__pfet_01v8_hvt__dlc_diff=0.0
+  sky130_fd_pr__pfet_01v8_hvt__dwc_diff=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 000, W = 1.26, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_0=0.33969
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_0=-0.026922
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_0=-0.00842
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_0=9.171e-20
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_0=0.0003608
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_0=-7416.8
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_0=0.027253
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_0=3.7374e-11
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_0=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 001, W = 1.68, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_1=0.60857
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_1=-0.032244
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_1=-2.2902e-19
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_1=-0.016292
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_1=0.0010674
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_1=-7426.8
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_1=0.011921
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_1=3.4586e-10
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_1=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 002, W = 1.0, L = 1.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_2=0.20802
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_2=0.013132
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_2=-0.017437
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_2=-0.038521
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_2=3.8706e-19
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_2=-0.0057008
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_2=0.0015329
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_2=-0.011623
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_2=-4.6376e-11
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 003, W = 1.0, L = 2.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_3=-1.9658e-11
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_3=0.28726
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_3=0.003295
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_3=-0.0028993
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_3=-0.026013
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_3=3.2924e-19
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_3=-0.0085614
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_3=0.0014549
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_3=0.0035651
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_3=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 004, W = 1.0, L = 4.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_4=-7.2896e-11
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_4=0.21396
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_4=-0.017589
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_4=0.041416
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_4=-0.040491
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_4=3.5687e-19
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_4=-0.0098132
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_4=0.0012235
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_4=-0.00088957
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_4=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 005, W = 1.0, L = 8.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_5=-3.4893e-11
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_5=0.26111
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_5=0.039675
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_5=-0.037542
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_5=-0.042255
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_5=3.6307e-19
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_5=-0.010815
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_5=0.001553
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_5=-0.0012827
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_5=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 006, W = 1.0, L = 0.15
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_6=3.469e-10
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_6=1.1311
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_6=-0.080838
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_6=-2.4224e-19
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_6=-0.025463
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_6=0.0012082
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_6=-1060.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_6=-0.00020238
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 007, W = 1.0, L = 0.18
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_7=-0.00072149
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_7=5.0661e-19
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_7=53782.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_7=-0.017309
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_7=-4.5014e-10
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_7=-0.13209
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_7=-0.037453
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_7=-0.0029197
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 008, W = 1.0, L = 0.25
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_8=-0.0052868
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_8=-0.00018539
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_8=-7.4084e-20
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_8=-2120.9
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_8=-0.0048221
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_8=1.6004e-10
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_8=0.56524
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_8=-0.027699
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 009, W = 1.0, L = 0.5
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_9=-0.042856
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_9=-0.009604
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_9=0.0014206
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_9=2.5647e-19
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_9=43209.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_9=0.0008166
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_9=5.7833e-11
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_9=0.11217
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 010, W = 3.0, L = 1.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_10=2.4575e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_10=-0.038563
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_10=-0.00053177
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_10=0.0019237
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_10=0.14974
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_10=0.00087842
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_10=0.0015678
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_10=-0.013242
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_10=-5.8082e-11
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 011, W = 3.0, L = 2.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_11=-3.411e-11
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_11=6.2077e-20
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_11=-0.047257
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_11=-0.0012709
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_11=0.0036608
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_11=0.21755
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_11=0.00029904
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_11=-0.00092696
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_11=-0.014467
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 012, W = 3.0, L = 4.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_12=-0.003503
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_12=-1.1408e-11
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_12=1.847e-20
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_12=0.00017941
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_12=-0.006186
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_12=0.0046314
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_12=1.1994
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_12=0.00025452
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_12=-0.00089931
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 013, W = 3.0, L = 8.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_13=1.2343
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_13=0.00012243
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_13=0.010767
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_13=-0.005387
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_13=-1.1232e-11
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_13=-2.0802e-21
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_13=-0.0079777
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_13=-0.0029371
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_13=0.0015899
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_13=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 014, W = 3.0, L = 0.15
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_14=-10254.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_14=0.28742
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_14=0.0003873
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_14=0.025528
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_14=-0.01124
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_14=3.7828e-11
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_14=7.0659e-20
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_14=-0.041324
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_14=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 015, W = 3.0, L = 0.18
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_15=32924.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_15=0.12614
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_15=0.00053254
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_15=-0.0089102
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_15=-0.013393
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_15=-1.4565e-11
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_15=2.0802e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_15=-0.05768
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_15=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 016, W = 3.0, L = 0.25
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_16=-1972.5
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_16=0.12457
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_16=0.00034854
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_16=-0.014326
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_16=0.0064619
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_16=5.6362e-12
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_16=1.7598e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_16=-0.029991
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_16=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 017, W = 3.0, L = 0.5
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_17=1.2823
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_17=0.00015563
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_17=165.11
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_17=0.0040546
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_17=-0.0031058
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_17=-1.1089e-11
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_17=4.2583e-20
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_17=-0.021129
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_17=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 018, W = 5.0, L = 1.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_18=0.048434
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_18=-0.065263
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_18=0.066563
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_18=0.0013661
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_18=-0.00096728
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_18=-0.011723
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_18=-9.6778e-11
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_18=4.4102e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_18=-0.040201
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 019, W = 5.0, L = 2.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_19=-0.044717
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_19=0.081124
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_19=-0.089078
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_19=0.16473
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_19=0.0012189
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_19=-0.0065271
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_19=-0.0077911
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_19=-2.0191e-10
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_19=5.2225e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_19=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 020, W = 5.0, L = 4.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_20=-0.037085
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_20=0.050634
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_20=-0.055889
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_20=0.2151
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_20=0.0019142
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_20=-0.0070601
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_20=-0.0071071
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_20=-1.9209e-10
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_20=6.3617e-19
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 021, W = 5.0, L = 8.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_21=6.067e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_21=-0.04099
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_21=0.019994
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_21=0.029645
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_21=-0.36321
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_21=-0.0010838
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_21=0.012193
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_21=-0.0044603
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_21=-6.1271e-10
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 022, W = 5.0, L = 0.15
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_22=4.0977e-11
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_22=2.7114e-20
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_22=-0.020779
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_22=-13087.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_22=0.23398
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_22=0.0003458
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_22=0.0095259
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_22=-0.011624
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 023, W = 5.0, L = 0.18
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_23=-0.0073835
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_23=1.6227e-10
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_23=7.6056e-20
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_23=-0.010974
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_23=18753.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_23=0.58698
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_23=0.0010731
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_23=0.0075373
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 024, W = 5.0, L = 0.25
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_24=0.077678
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_24=0.00033325
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_24=-0.014274
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_24=-0.0045308
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_24=-5.212e-11
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_24=2.6633e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_24=-0.030909
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_24=9905.6
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 025, W = 5.0, L = 0.5
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_25=44080.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_25=-0.33053
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_25=-1.5876e-5
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_25=0.0066358
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_25=-0.0099005
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_25=-1.5878e-10
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_25=2.6336e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_25=-0.03415
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_25=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 026, W = 7.0, L = 1.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_26=-0.00032957
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_26=0.0018471
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_26=-0.0071289
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_26=-0.0095046
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_26=-1.4936e-10
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_26=5.6221e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_26=-0.044741
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_26=0.075088
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_26=-0.099607
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_26=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 027, W = 7.0, L = 2.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_27=0.089097
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_27=0.0018216
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_27=-0.003648
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_27=-0.007636
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_27=-1.7667e-10
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_27=5.8807e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_27=-0.030487
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_27=0.0713
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_27=-0.080217
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_27=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 028, W = 7.0, L = 4.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_28=1.2166
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_28=0.0014352
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_28=0.0091366
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_28=-0.0053636
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_28=-1.3672e-11
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_28=2.9847e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_28=-0.0059034
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_28=0.016269
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_28=-0.0091092
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 029, W = 7.0, L = 8.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_29=0.0032924
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_29=-0.0026106
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_29=1.2187
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_29=0.0017419
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_29=0.0035905
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_29=-0.0088595
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_29=-1.4852e-11
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_29=3.3671e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_29=-0.0078252
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 030, W = 7.0, L = 0.15
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_30=-0.028843
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_30=-6543.4
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_30=0.61482
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_30=0.0012299
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_30=0.0025174
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_30=-0.029749
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_30=3.1813e-10
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_30=-1.8716e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_30=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 031, W = 7.0, L = 0.18
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_31=-0.047465
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_31=23924.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_31=0.10005
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_31=0.00013514
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_31=-0.019852
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_31=-0.011281
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_31=-1.4225e-10
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_31=3.0833e-19
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 032, W = 7.0, L = 0.25
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_32=1.6451e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_32=-0.032636
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_32=1010.5
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_32=0.12366
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_32=0.00016779
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_32=-0.0046762
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_32=-0.0028117
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_32=-1.7243e-11
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 033, W = 7.0, L = 0.5
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_33=-2.4885e-11
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_33=2.5424e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_33=-0.01298
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_33=31235.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_33=1.2891
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_33=0.0010899
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_33=-0.0053108
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_33=-0.010171
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 034, W = 0.42, L = 1.0
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_34=-0.0031312
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_34=-2.371e-11
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_34=3.4376e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_34=-0.054193
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_34=-6.4067e-8
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_34=1.7873e-10
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_34=1.387
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_34=0.0014966
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_34=-0.012619
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 035, W = 0.42, L = 20.0
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_35=0.22953
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_35=0.0021307
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_35=-0.044112
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_35=-0.009361
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_35=-1.4456e-10
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_35=5.2005e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_35=-0.055437
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_35=-8.762e-8
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_35=-6.7636e-9
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_35=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 036, W = 0.42, L = 2.0
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_36=1.2381
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_36=-0.00021399
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_36=0.0051836
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_36=0.0069385
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_36=-9.0008e-12
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_36=-2.4281e-20
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_36=-0.01182
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_36=2.0301e-8
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_36=1.2557e-11
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 037, W = 0.42, L = 4.0
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_37=-2.1753e-9
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_37=0.22912
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_37=0.0020212
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_37=-0.021515
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_37=-0.0055742
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_37=-1.3629e-10
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_37=5.3159e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_37=-0.050147
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_37=-5.1402e-8
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_37=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 038, W = 0.42, L = 8.0
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_38=-2.5362e-8
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_38=-5.6582e-12
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_38=1.2423
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_38=0.00075206
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_38=-0.020202
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_38=-0.0019647
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_38=-2.527e-11
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_38=9.7792e-20
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_38=-0.015728
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_38=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 039, W = 0.42, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_39=0.86891
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_39=0.00046554
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_39=2238.5
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_39=0.040258
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_39=-0.0064094
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_39=7.7102e-11
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_39=8.1554e-20
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_39=-0.075719
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_39=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 040, W = 0.42, L = 0.18
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_40=32843.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_40=0.046556
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_40=-0.00098229
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_40=0.027158
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_40=-0.0075535
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_40=-4.8538e-10
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_40=4.9561e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_40=-0.074451
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_40=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 041, W = 0.42, L = 0.5
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_41=-0.040166
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_41=23061.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_41=1.4109
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_41=0.00077482
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_41=0.029596
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_41=-0.010991
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_41=-2.5485e-11
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_41=2.1997e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_41=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 042, W = 0.55, L = 1.0
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_42=-0.06677
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_42=-9.3827e-8
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_42=-1.2472e-10
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_42=0.29746
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_42=0.0021119
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_42=-0.019844
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_42=-0.010603
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_42=1.1179e-10
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_42=2.6904e-19
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 043, W = 0.55, L = 2.0
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_43=3.8482e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_43=-0.042159
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_43=-3.9783e-8
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_43=-1.5632e-9
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_43=0.27193
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_43=0.0013084
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_43=-0.0037886
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_43=-0.0028399
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_43=-5.5028e-11
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 044, W = 0.55, L = 4.0
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_44=-8.7318e-11
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_44=4.68e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_44=-0.046546
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_44=-6.9914e-8
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_44=2.0353e-10
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_44=0.29301
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_44=0.0018679
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_44=-0.011246
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_44=-0.0048261
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 045, W = 0.55, L = 8.0
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_45=0.00053147
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_45=-4.9698e-12
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_45=-3.4539e-20
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_45=-0.017283
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_45=2.2471e-8
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_45=2.9204e-11
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_45=0.088947
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_45=5.5852e-5
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_45=0.013275
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 046, W = 0.55, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_46=0.67021
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_46=0.00071212
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_46=-0.012126
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_46=-0.02751
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_46=1.5449e-10
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_46=-2.8376e-20
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_46=-0.047133
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_46=8984.7
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 047, W = 0.55, L = 0.5
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_47=-13168.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_47=1.3992
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_47=0.00092803
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_47=0.01785
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_47=-0.0026549
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_47=1.1727e-12
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_47=2.7682e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_47=-0.03499
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_47=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 048, W = 0.64, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_48=5421.6
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_48=0.80607
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_48=-3.1943e-5
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_48=0.018044
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_48=-0.0084157
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_48=-8.6721e-11
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_48=1.5947e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_48=-0.092261
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_48=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 049, W = 0.84, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_49=-6146.4
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_49=1.4145
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_49=0.00019282
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_49=0.048161
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_49=-0.01019
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_49=-7.9353e-12
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_49=7.604e-20
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_49=-0.049003
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_49=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 050, W = 0.64, L = 0.18
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_50=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 051, W = 2.0, L = 0.15
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_51=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 052, W = 1.12, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_52=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 053, W = 1.65, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_53=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 054, W = 0.84, L = 0.18
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_54=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 055, W = 1.68, L = 0.18
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_55=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 056, W = 0.36, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_56=-0.020934
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_56=81981.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_56=-0.00017582
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_56=0.020586
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 057, W = 0.54, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_57=-0.00017618
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_57=0.0039256
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_57=-0.014348
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_57=78372.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_57=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 058, W = 0.63, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_58=36202.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_58=-0.00020189
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_58=0.0075757
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_58=-0.015801
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_58=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 059, W = 0.7, L = 0.15
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_59=25602.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_59=-0.00016346
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_59=0.0034029
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_59=-0.014445
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_59=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 060, W = 0.75, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_60=25454.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_60=-0.0001819
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_60=0.0026511
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_60=-0.013785
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_60=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 061, W = 0.79, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_61=36053.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_61=-0.00021998
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_61=0.0019836
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_61=-0.013308
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_61=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 062, W = 0.82, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_62=37969.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_62=-0.00022145
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_62=0.0036256
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_62=-0.011949
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_62=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 063, W = 0.82, L = 0.18
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_63=27669.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_63=-0.00015603
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_63=0.0066454
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_63=-0.0098916
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_63=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 064, W = 0.82, L = 0.25
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_64=58607.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_64=-0.00011722
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_64=-0.0043943
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_64=-0.0068897
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_64=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 065, W = 0.82, L = 0.5
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_65=51004.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_65=-0.00031453
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_65=0.0021112
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_65=-0.0073046
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_65=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 066, W = 0.86, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_66=52818.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_66=-0.0002412
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_66=0.0035355
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_66=-0.012563
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 067, W = 0.94, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_67=-0.01279
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_67=64603.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_67=-0.00029595
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_67=0.0072012
.include "sky130_fd_pr__pfet_01v8_hvt__tt.pm3.spice"
