* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 52
.param
+  sky130_fd_pr__pfet_01v8__toxe_mult=1.0
+  sky130_fd_pr__pfet_01v8__rshp_mult=1.0
+  sky130_fd_pr__pfet_01v8__overlap_mult=0.95435
+  sky130_fd_pr__pfet_01v8__ajunction_mult=0.99626
+  sky130_fd_pr__pfet_01v8__pjunction_mult=1.0009
+  sky130_fd_pr__pfet_01v8__lint_diff=0.0
+  sky130_fd_pr__pfet_01v8__wint_diff=0.0
+  sky130_fd_pr__pfet_01v8__dlc_diff=0.0
+  sky130_fd_pr__pfet_01v8__dwc_diff=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 000, W = 1.26, L = 0.15
* -----------------------------------
+  sky130_fd_pr__pfet_01v8__agidl_diff_0=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_0=0.25683
+  sky130_fd_pr__pfet_01v8__vsat_diff_0=16185.0
+  sky130_fd_pr__pfet_01v8__a0_diff_0=0.0
+  sky130_fd_pr__pfet_01v8__pdits_diff_0=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_0=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_0=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_0=0.030227
+  sky130_fd_pr__pfet_01v8__eta0_diff_0=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_0=-1.0309e-11
+  sky130_fd_pr__pfet_01v8__keta_diff_0=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_0=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_0=-0.019468
+  sky130_fd_pr__pfet_01v8__vth0_diff_0=0.036794
+  sky130_fd_pr__pfet_01v8__pditsd_diff_0=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_0=0.00038711
+  sky130_fd_pr__pfet_01v8__b1_diff_0=0.0
+  sky130_fd_pr__pfet_01v8__cgidl_diff_0=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_0=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_0=-0.078458
+  sky130_fd_pr__pfet_01v8__ags_diff_0=0.0
+  sky130_fd_pr__pfet_01v8__bgidl_diff_0=0.0
+  sky130_fd_pr__pfet_01v8__ub_diff_0=2.3766e-19
*
* sky130_fd_pr__pfet_01v8, Bin 001, W = 1.68, L = 0.15
* -----------------------------------
+  sky130_fd_pr__pfet_01v8__bgidl_diff_1=0.0
+  sky130_fd_pr__pfet_01v8__ub_diff_1=1.9928e-19
+  sky130_fd_pr__pfet_01v8__agidl_diff_1=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_1=0.065612
+  sky130_fd_pr__pfet_01v8__vsat_diff_1=-522.1
+  sky130_fd_pr__pfet_01v8__a0_diff_1=0.0
+  sky130_fd_pr__pfet_01v8__pdits_diff_1=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_1=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_1=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_1=0.079136
+  sky130_fd_pr__pfet_01v8__eta0_diff_1=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_1=-2.9528e-11
+  sky130_fd_pr__pfet_01v8__keta_diff_1=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_1=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_1=-0.023277
+  sky130_fd_pr__pfet_01v8__vth0_diff_1=-0.015775
+  sky130_fd_pr__pfet_01v8__pditsd_diff_1=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_1=0.0003417
+  sky130_fd_pr__pfet_01v8__b1_diff_1=0.0
+  sky130_fd_pr__pfet_01v8__cgidl_diff_1=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_1=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_1=-0.021939
+  sky130_fd_pr__pfet_01v8__ags_diff_1=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 002, W = 1.0, L = 1.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__cgidl_diff_2=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_2=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_2=-0.065739
+  sky130_fd_pr__pfet_01v8__ags_diff_2=0.082231
+  sky130_fd_pr__pfet_01v8__bgidl_diff_2=0.0
+  sky130_fd_pr__pfet_01v8__ub_diff_2=3.0975e-19
+  sky130_fd_pr__pfet_01v8__agidl_diff_2=-2.7915e-12
+  sky130_fd_pr__pfet_01v8__nfactor_diff_2=-0.079944
+  sky130_fd_pr__pfet_01v8__vsat_diff_2=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_2=-0.079498
+  sky130_fd_pr__pfet_01v8__pdits_diff_2=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_2=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_2=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_2=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_2=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_2=-1.8999e-11
+  sky130_fd_pr__pfet_01v8__keta_diff_2=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_2=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_2=-0.010076
+  sky130_fd_pr__pfet_01v8__vth0_diff_2=-0.0057939
+  sky130_fd_pr__pfet_01v8__pditsd_diff_2=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_2=0.0014217
+  sky130_fd_pr__pfet_01v8__b1_diff_2=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 003, W = 1.0, L = 2.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__b1_diff_3=0.0
+  sky130_fd_pr__pfet_01v8__cgidl_diff_3=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_3=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_3=-0.068427
+  sky130_fd_pr__pfet_01v8__ags_diff_3=0.061811
+  sky130_fd_pr__pfet_01v8__bgidl_diff_3=0.0
+  sky130_fd_pr__pfet_01v8__ub_diff_3=3.4961e-19
+  sky130_fd_pr__pfet_01v8__nfactor_diff_3=0.074091
+  sky130_fd_pr__pfet_01v8__vsat_diff_3=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_3=-1.6202e-10
+  sky130_fd_pr__pfet_01v8__a0_diff_3=-0.070079
+  sky130_fd_pr__pfet_01v8__pdits_diff_3=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_3=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_3=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_3=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_3=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_3=-8.1128e-12
+  sky130_fd_pr__pfet_01v8__keta_diff_3=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_3=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_3=-0.013508
+  sky130_fd_pr__pfet_01v8__vth0_diff_3=-0.00071929
+  sky130_fd_pr__pfet_01v8__pditsd_diff_3=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_3=0.0015781
*
* sky130_fd_pr__pfet_01v8, Bin 004, W = 1.0, L = 4.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__pditsd_diff_4=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_4=0.0015543
+  sky130_fd_pr__pfet_01v8__vth0_diff_4=-0.013029
+  sky130_fd_pr__pfet_01v8__b1_diff_4=0.0
+  sky130_fd_pr__pfet_01v8__cgidl_diff_4=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_4=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_4=-0.066359
+  sky130_fd_pr__pfet_01v8__ags_diff_4=0.043153
+  sky130_fd_pr__pfet_01v8__ub_diff_4=3.2388e-19
+  sky130_fd_pr__pfet_01v8__bgidl_diff_4=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_4=0.065236
+  sky130_fd_pr__pfet_01v8__vsat_diff_4=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_4=3.2697e-11
+  sky130_fd_pr__pfet_01v8__a0_diff_4=-0.04408
+  sky130_fd_pr__pfet_01v8__pdits_diff_4=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_4=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_4=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_4=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_4=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_4=-7.8248e-12
+  sky130_fd_pr__pfet_01v8__keta_diff_4=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_4=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_4=-0.014149
*
* sky130_fd_pr__pfet_01v8, Bin 005, W = 1.0, L = 8.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__keta_diff_5=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_5=-0.01529
+  sky130_fd_pr__pfet_01v8__pditsd_diff_5=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_5=0.0014113
+  sky130_fd_pr__pfet_01v8__vth0_diff_5=-0.023685
+  sky130_fd_pr__pfet_01v8__b1_diff_5=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_5=-0.073497
+  sky130_fd_pr__pfet_01v8__cgidl_diff_5=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_5=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_5=0.085722
+  sky130_fd_pr__pfet_01v8__ub_diff_5=3.2181e-19
+  sky130_fd_pr__pfet_01v8__bgidl_diff_5=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_5=0.086719
+  sky130_fd_pr__pfet_01v8__vsat_diff_5=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_5=-2.7806e-11
+  sky130_fd_pr__pfet_01v8__a0_diff_5=-0.081463
+  sky130_fd_pr__pfet_01v8__pdits_diff_5=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_5=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_5=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_5=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_5=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_5=-2.3572e-11
+  sky130_fd_pr__pfet_01v8__rdsw_diff_5=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 006, W = 1.0, L = 0.15
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__rdsw_diff_6=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_6=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_6=-0.025848
+  sky130_fd_pr__pfet_01v8__pditsd_diff_6=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_6=0.00044044
+  sky130_fd_pr__pfet_01v8__vth0_diff_6=-0.050863
+  sky130_fd_pr__pfet_01v8__b1_diff_6=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_6=0.0086622
+  sky130_fd_pr__pfet_01v8__cgidl_diff_6=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_6=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_6=0.0
+  sky130_fd_pr__pfet_01v8__ub_diff_6=2.1528e-19
+  sky130_fd_pr__pfet_01v8__bgidl_diff_6=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_6=-0.2601
+  sky130_fd_pr__pfet_01v8__vsat_diff_6=-16.083
+  sky130_fd_pr__pfet_01v8__agidl_diff_6=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_6=0.0
+  sky130_fd_pr__pfet_01v8__pdits_diff_6=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_6=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_6=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_6=0.098454
+  sky130_fd_pr__pfet_01v8__eta0_diff_6=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_6=-2.6963e-11
*
* sky130_fd_pr__pfet_01v8, Bin 007, W = 1.0, L = 0.18
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__kt1_diff_7=0.031634
+  sky130_fd_pr__pfet_01v8__eta0_diff_7=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_7=-2.9267e-11
+  sky130_fd_pr__pfet_01v8__rdsw_diff_7=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_7=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_7=-0.018493
+  sky130_fd_pr__pfet_01v8__pditsd_diff_7=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_7=0.00019975
+  sky130_fd_pr__pfet_01v8__vth0_diff_7=-0.036221
+  sky130_fd_pr__pfet_01v8__b1_diff_7=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_7=-0.083056
+  sky130_fd_pr__pfet_01v8__cgidl_diff_7=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_7=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_7=0.0
+  sky130_fd_pr__pfet_01v8__ub_diff_7=1.8997e-19
+  sky130_fd_pr__pfet_01v8__bgidl_diff_7=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_7=0.26714
+  sky130_fd_pr__pfet_01v8__vsat_diff_7=20157.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_7=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_7=0.0
+  sky130_fd_pr__pfet_01v8__pdits_diff_7=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_7=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_7=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 008, W = 1.0, L = 0.25
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__pclm_diff_8=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_8=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_8=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_8=-2.1298e-11
+  sky130_fd_pr__pfet_01v8__rdsw_diff_8=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_8=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_8=-0.0092316
+  sky130_fd_pr__pfet_01v8__pditsd_diff_8=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_8=-0.00054137
+  sky130_fd_pr__pfet_01v8__vth0_diff_8=0.020531
+  sky130_fd_pr__pfet_01v8__b1_diff_8=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_8=-0.070563
+  sky130_fd_pr__pfet_01v8__cgidl_diff_8=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_8=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_8=0.0
+  sky130_fd_pr__pfet_01v8__ub_diff_8=1.5069e-19
+  sky130_fd_pr__pfet_01v8__bgidl_diff_8=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_8=-0.027492
+  sky130_fd_pr__pfet_01v8__vsat_diff_8=52493.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_8=6.0957e-10
+  sky130_fd_pr__pfet_01v8__a0_diff_8=0.0
+  sky130_fd_pr__pfet_01v8__pdits_diff_8=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_8=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 009, W = 1.0, L = 0.5
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__pdits_diff_9=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_9=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_9=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_9=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_9=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_9=-7.015e-12
+  sky130_fd_pr__pfet_01v8__rdsw_diff_9=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_9=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_9=-0.01065
+  sky130_fd_pr__pfet_01v8__pditsd_diff_9=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_9=0.00058728
+  sky130_fd_pr__pfet_01v8__vth0_diff_9=0.046674
+  sky130_fd_pr__pfet_01v8__b1_diff_9=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_9=-0.056914
+  sky130_fd_pr__pfet_01v8__cgidl_diff_9=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_9=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_9=0.0
+  sky130_fd_pr__pfet_01v8__ub_diff_9=2.4247e-19
+  sky130_fd_pr__pfet_01v8__bgidl_diff_9=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_9=-0.0015401
+  sky130_fd_pr__pfet_01v8__vsat_diff_9=-16234.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_9=-2.7085e-10
+  sky130_fd_pr__pfet_01v8__a0_diff_9=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 010, W = 2.0, L = 0.15
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__pditsd_diff_10=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_10=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_10=4327.8
+  sky130_fd_pr__pfet_01v8__u0_diff_10=0.00042484
+  sky130_fd_pr__pfet_01v8__vth0_diff_10=-0.051412
+  sky130_fd_pr__pfet_01v8__cgidl_diff_10=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_10=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_10=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_10=0.099019
+  sky130_fd_pr__pfet_01v8__pclm_diff_10=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_10=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_10=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_10=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_10=-2.6742e-11
+  sky130_fd_pr__pfet_01v8__bgidl_diff_10=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_10=0.077506
+  sky130_fd_pr__pfet_01v8__ub_diff_10=2.047e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_10=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_10=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_10=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_10=-0.018259
+  sky130_fd_pr__pfet_01v8__voff_diff_10=-0.030945
+  sky130_fd_pr__pfet_01v8__a0_diff_10=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 011, W = 3.0, L = 1.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__voff_diff_11=-0.055855
+  sky130_fd_pr__pfet_01v8__a0_diff_11=-0.086686
+  sky130_fd_pr__pfet_01v8__pditsd_diff_11=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_11=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_11=26714.0
+  sky130_fd_pr__pfet_01v8__u0_diff_11=0.0013927
+  sky130_fd_pr__pfet_01v8__vth0_diff_11=-0.014123
+  sky130_fd_pr__pfet_01v8__cgidl_diff_11=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_11=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_11=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_11=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_11=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_11=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_11=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_11=1.6673e-10
+  sky130_fd_pr__pfet_01v8__ua_diff_11=-3.8e-11
+  sky130_fd_pr__pfet_01v8__bgidl_diff_11=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_11=-0.025198
+  sky130_fd_pr__pfet_01v8__ub_diff_11=3.7335e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_11=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_11=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_11=0.067844
+  sky130_fd_pr__pfet_01v8__k2_diff_11=-0.015275
*
* sky130_fd_pr__pfet_01v8, Bin 012, W = 3.0, L = 2.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__pdits_diff_12=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_12=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_12=0.06063
+  sky130_fd_pr__pfet_01v8__k2_diff_12=-0.010456
+  sky130_fd_pr__pfet_01v8__voff_diff_12=-0.051762
+  sky130_fd_pr__pfet_01v8__a0_diff_12=-0.071465
+  sky130_fd_pr__pfet_01v8__pditsd_diff_12=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_12=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_12=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_12=0.0018111
+  sky130_fd_pr__pfet_01v8__vth0_diff_12=-0.010167
+  sky130_fd_pr__pfet_01v8__cgidl_diff_12=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_12=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_12=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_12=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_12=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_12=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_12=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_12=-1.1943e-10
+  sky130_fd_pr__pfet_01v8__ua_diff_12=-7.0667e-12
+  sky130_fd_pr__pfet_01v8__bgidl_diff_12=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_12=0.011369
+  sky130_fd_pr__pfet_01v8__ub_diff_12=3.9754e-19
*
* sky130_fd_pr__pfet_01v8, Bin 013, W = 3.0, L = 4.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__bgidl_diff_13=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_13=0.046528
+  sky130_fd_pr__pfet_01v8__ub_diff_13=3.83e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_13=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_13=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_13=0.035284
+  sky130_fd_pr__pfet_01v8__k2_diff_13=-0.0085688
+  sky130_fd_pr__pfet_01v8__voff_diff_13=-0.048343
+  sky130_fd_pr__pfet_01v8__a0_diff_13=-0.040581
+  sky130_fd_pr__pfet_01v8__eta0_diff_13=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_13=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_13=0.0017986
+  sky130_fd_pr__pfet_01v8__vsat_diff_13=0.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_13=-0.00035349
+  sky130_fd_pr__pfet_01v8__cgidl_diff_13=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_13=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_13=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_13=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_13=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_13=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_13=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_13=-8.903e-11
+  sky130_fd_pr__pfet_01v8__ua_diff_13=-2.9121e-12
*
* sky130_fd_pr__pfet_01v8, Bin 014, W = 3.0, L = 8.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__agidl_diff_14=8.2999e-10
+  sky130_fd_pr__pfet_01v8__b1_diff_14=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_14=-4.0591e-12
+  sky130_fd_pr__pfet_01v8__bgidl_diff_14=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_14=0.038794
+  sky130_fd_pr__pfet_01v8__ub_diff_14=4.1037e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_14=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_14=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_14=0.01599
+  sky130_fd_pr__pfet_01v8__k2_diff_14=-0.008116
+  sky130_fd_pr__pfet_01v8__voff_diff_14=-0.038421
+  sky130_fd_pr__pfet_01v8__eta0_diff_14=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_14=-0.020004
+  sky130_fd_pr__pfet_01v8__pditsd_diff_14=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_14=0.0019508
+  sky130_fd_pr__pfet_01v8__vsat_diff_14=0.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_14=0.0024267
+  sky130_fd_pr__pfet_01v8__cgidl_diff_14=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_14=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_14=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_14=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_14=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_14=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 015, W = 3.0, L = 0.15
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__b0_diff_15=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_15=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_15=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_15=5.2325e-13
+  sky130_fd_pr__pfet_01v8__bgidl_diff_15=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_15=-0.1522
+  sky130_fd_pr__pfet_01v8__ub_diff_15=1.6415e-19
+  sky130_fd_pr__pfet_01v8__tvoff_diff_15=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_15=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_15=-0.019065
+  sky130_fd_pr__pfet_01v8__pdits_diff_15=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_15=0.023584
+  sky130_fd_pr__pfet_01v8__eta0_diff_15=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_15=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_15=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_15=0.00043907
+  sky130_fd_pr__pfet_01v8__vsat_diff_15=-7488.9
+  sky130_fd_pr__pfet_01v8__vth0_diff_15=-0.025245
+  sky130_fd_pr__pfet_01v8__cgidl_diff_15=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_15=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_15=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_15=0.11486
+  sky130_fd_pr__pfet_01v8__pclm_diff_15=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 016, W = 3.0, L = 0.18
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__pclm_diff_16=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_16=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_16=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_16=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_16=2.0071e-12
+  sky130_fd_pr__pfet_01v8__bgidl_diff_16=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_16=0.34132
+  sky130_fd_pr__pfet_01v8__tvoff_diff_16=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_16=0.0
+  sky130_fd_pr__pfet_01v8__ub_diff_16=1.9453e-19
+  sky130_fd_pr__pfet_01v8__k2_diff_16=-0.015561
+  sky130_fd_pr__pfet_01v8__pdits_diff_16=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_16=-0.077978
+  sky130_fd_pr__pfet_01v8__eta0_diff_16=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_16=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_16=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_16=0.00055238
+  sky130_fd_pr__pfet_01v8__vsat_diff_16=8562.4
+  sky130_fd_pr__pfet_01v8__vth0_diff_16=-0.0057149
+  sky130_fd_pr__pfet_01v8__cgidl_diff_16=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_16=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_16=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_16=-0.20389
*
* sky130_fd_pr__pfet_01v8, Bin 017, W = 3.0, L = 0.25
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__kt1_diff_17=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_17=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_17=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_17=2.8433e-13
+  sky130_fd_pr__pfet_01v8__b1_diff_17=0.0
+  sky130_fd_pr__pfet_01v8__bgidl_diff_17=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_17=-0.057073
+  sky130_fd_pr__pfet_01v8__ua_diff_17=-5.0889e-11
+  sky130_fd_pr__pfet_01v8__tvoff_diff_17=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_17=0.0
+  sky130_fd_pr__pfet_01v8__ub_diff_17=2.6612e-19
+  sky130_fd_pr__pfet_01v8__k2_diff_17=-0.0073251
+  sky130_fd_pr__pfet_01v8__pdits_diff_17=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_17=-0.089917
+  sky130_fd_pr__pfet_01v8__eta0_diff_17=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_17=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_17=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_17=-0.0007821
+  sky130_fd_pr__pfet_01v8__vsat_diff_17=-20000.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_17=0.16959
+  sky130_fd_pr__pfet_01v8__cgidl_diff_17=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_17=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_17=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 018, W = 3.0, L = 0.5
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__rdsw_diff_18=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_18=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_18=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_18=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_18=-1.6447e-10
+  sky130_fd_pr__pfet_01v8__b1_diff_18=0.0
+  sky130_fd_pr__pfet_01v8__bgidl_diff_18=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_18=0.13485
+  sky130_fd_pr__pfet_01v8__ua_diff_18=9.2994e-13
+  sky130_fd_pr__pfet_01v8__tvoff_diff_18=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_18=0.0
+  sky130_fd_pr__pfet_01v8__ub_diff_18=2.2388e-19
+  sky130_fd_pr__pfet_01v8__k2_diff_18=-0.015495
+  sky130_fd_pr__pfet_01v8__pdits_diff_18=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_18=-0.058923
+  sky130_fd_pr__pfet_01v8__eta0_diff_18=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_18=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_18=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_18=0.00093447
+  sky130_fd_pr__pfet_01v8__vsat_diff_18=15814.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_18=0.0018962
+  sky130_fd_pr__pfet_01v8__cgidl_diff_18=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_18=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 019, W = 5.0, L = 1.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__cgidl_diff_19=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_19=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_19=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_19=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_19=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_19=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_19=1.357e-11
+  sky130_fd_pr__pfet_01v8__b1_diff_19=0.0
+  sky130_fd_pr__pfet_01v8__bgidl_diff_19=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_19=-0.039041
+  sky130_fd_pr__pfet_01v8__ua_diff_19=-9.3266e-12
+  sky130_fd_pr__pfet_01v8__tvoff_diff_19=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_19=0.040613
+  sky130_fd_pr__pfet_01v8__ub_diff_19=2.6349e-19
+  sky130_fd_pr__pfet_01v8__k2_diff_19=-0.009616
+  sky130_fd_pr__pfet_01v8__pdits_diff_19=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_19=-0.038421
+  sky130_fd_pr__pfet_01v8__eta0_diff_19=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_19=-0.044426
+  sky130_fd_pr__pfet_01v8__pditsd_diff_19=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_19=0.0010966
+  sky130_fd_pr__pfet_01v8__vsat_diff_19=0.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_19=0.0069077
*
* sky130_fd_pr__pfet_01v8, Bin 020, W = 5.0, L = 2.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__u0_diff_20=0.0012594
+  sky130_fd_pr__pfet_01v8__vth0_diff_20=0.0013804
+  sky130_fd_pr__pfet_01v8__cgidl_diff_20=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_20=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_20=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_20=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_20=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_20=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_20=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_20=1.1728e-10
+  sky130_fd_pr__pfet_01v8__ua_diff_20=-3.626e-12
+  sky130_fd_pr__pfet_01v8__bgidl_diff_20=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_20=0.048112
+  sky130_fd_pr__pfet_01v8__ub_diff_20=2.7353e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_20=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_20=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_20=0.034607
+  sky130_fd_pr__pfet_01v8__k2_diff_20=-0.011931
+  sky130_fd_pr__pfet_01v8__voff_diff_20=-0.043221
+  sky130_fd_pr__pfet_01v8__a0_diff_20=-0.039408
+  sky130_fd_pr__pfet_01v8__pditsd_diff_20=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_20=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_20=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 021, W = 5.0, L = 4.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__pditsd_diff_21=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_21=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_21=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_21=0.0016296
+  sky130_fd_pr__pfet_01v8__vth0_diff_21=0.0048253
+  sky130_fd_pr__pfet_01v8__cgidl_diff_21=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_21=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_21=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_21=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_21=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_21=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_21=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_21=7.7837e-10
+  sky130_fd_pr__pfet_01v8__ua_diff_21=-2.4508e-12
+  sky130_fd_pr__pfet_01v8__bgidl_diff_21=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_21=0.056607
+  sky130_fd_pr__pfet_01v8__ub_diff_21=3.1849e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_21=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_21=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_21=0.011085
+  sky130_fd_pr__pfet_01v8__k2_diff_21=-0.011887
+  sky130_fd_pr__pfet_01v8__voff_diff_21=-0.043022
+  sky130_fd_pr__pfet_01v8__a0_diff_21=-0.012572
*
* sky130_fd_pr__pfet_01v8, Bin 022, W = 5.0, L = 8.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__voff_diff_22=-0.041062
+  sky130_fd_pr__pfet_01v8__a0_diff_22=-0.011407
+  sky130_fd_pr__pfet_01v8__pditsd_diff_22=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_22=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_22=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_22=0.001794
+  sky130_fd_pr__pfet_01v8__vth0_diff_22=0.00087396
+  sky130_fd_pr__pfet_01v8__cgidl_diff_22=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_22=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_22=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_22=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_22=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_22=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_22=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_22=1.2773e-9
+  sky130_fd_pr__pfet_01v8__ua_diff_22=-2.9796e-12
+  sky130_fd_pr__pfet_01v8__bgidl_diff_22=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_22=0.060845
+  sky130_fd_pr__pfet_01v8__ub_diff_22=3.5456e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_22=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_22=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_22=0.0099914
+  sky130_fd_pr__pfet_01v8__k2_diff_22=-0.012109
*
* sky130_fd_pr__pfet_01v8, Bin 023, W = 5.0, L = 0.15
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__pdits_diff_23=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_23=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_23=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_23=-0.014758
+  sky130_fd_pr__pfet_01v8__voff_diff_23=-0.030087
+  sky130_fd_pr__pfet_01v8__a0_diff_23=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_23=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_23=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_23=-3146.0
+  sky130_fd_pr__pfet_01v8__u0_diff_23=0.00043545
+  sky130_fd_pr__pfet_01v8__vth0_diff_23=-0.024632
+  sky130_fd_pr__pfet_01v8__cgidl_diff_23=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_23=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_23=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_23=0.10927
+  sky130_fd_pr__pfet_01v8__pclm_diff_23=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_23=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_23=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_23=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_23=-1.5205e-12
+  sky130_fd_pr__pfet_01v8__bgidl_diff_23=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_23=0.092629
+  sky130_fd_pr__pfet_01v8__ub_diff_23=1.6711e-19
*
* sky130_fd_pr__pfet_01v8, Bin 024, W = 5.0, L = 0.18
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__bgidl_diff_24=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_24=0.42606
+  sky130_fd_pr__pfet_01v8__ub_diff_24=1.6768e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_24=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_24=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_24=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_24=-0.011236
+  sky130_fd_pr__pfet_01v8__voff_diff_24=-0.10182
+  sky130_fd_pr__pfet_01v8__a0_diff_24=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_24=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_24=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_24=0.0003261
+  sky130_fd_pr__pfet_01v8__vsat_diff_24=15348.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_24=-0.016664
+  sky130_fd_pr__pfet_01v8__cgidl_diff_24=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_24=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_24=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_24=-0.10745
+  sky130_fd_pr__pfet_01v8__pclm_diff_24=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_24=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_24=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_24=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_24=-8.5792e-12
*
* sky130_fd_pr__pfet_01v8, Bin 025, W = 5.0, L = 0.25
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__agidl_diff_25=6.3147e-10
+  sky130_fd_pr__pfet_01v8__b1_diff_25=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_25=-5.3917e-13
+  sky130_fd_pr__pfet_01v8__bgidl_diff_25=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_25=0.11082
+  sky130_fd_pr__pfet_01v8__ub_diff_25=2.4381e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_25=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_25=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_25=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_25=-0.0081573
+  sky130_fd_pr__pfet_01v8__voff_diff_25=-0.067969
+  sky130_fd_pr__pfet_01v8__eta0_diff_25=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_25=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_25=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_25=0.00060874
+  sky130_fd_pr__pfet_01v8__vsat_diff_25=7603.4
+  sky130_fd_pr__pfet_01v8__vth0_diff_25=-0.02575
+  sky130_fd_pr__pfet_01v8__cgidl_diff_25=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_25=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_25=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_25=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_25=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_25=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 026, W = 5.0, L = 0.5
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__b0_diff_26=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_26=4.045e-11
+  sky130_fd_pr__pfet_01v8__b1_diff_26=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_26=5.7453e-12
+  sky130_fd_pr__pfet_01v8__bgidl_diff_26=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_26=0.17526
+  sky130_fd_pr__pfet_01v8__ub_diff_26=2.8055e-19
+  sky130_fd_pr__pfet_01v8__tvoff_diff_26=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_26=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_26=-0.015244
+  sky130_fd_pr__pfet_01v8__pdits_diff_26=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_26=-0.041918
+  sky130_fd_pr__pfet_01v8__eta0_diff_26=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_26=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_26=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_26=0.0012472
+  sky130_fd_pr__pfet_01v8__vsat_diff_26=7609.4
+  sky130_fd_pr__pfet_01v8__vth0_diff_26=-0.0033953
+  sky130_fd_pr__pfet_01v8__cgidl_diff_26=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_26=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_26=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_26=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_26=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 027, W = 7.0, L = 1.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__pclm_diff_27=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_27=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_27=6.8302e-11
+  sky130_fd_pr__pfet_01v8__b1_diff_27=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_27=-1.0829e-11
+  sky130_fd_pr__pfet_01v8__bgidl_diff_27=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_27=-0.077875
+  sky130_fd_pr__pfet_01v8__tvoff_diff_27=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_27=0.091645
+  sky130_fd_pr__pfet_01v8__ub_diff_27=2.9028e-19
+  sky130_fd_pr__pfet_01v8__k2_diff_27=-0.01015
+  sky130_fd_pr__pfet_01v8__pdits_diff_27=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_27=-0.031586
+  sky130_fd_pr__pfet_01v8__eta0_diff_27=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_27=-0.13367
+  sky130_fd_pr__pfet_01v8__pditsd_diff_27=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_27=0.0012177
+  sky130_fd_pr__pfet_01v8__vsat_diff_27=0.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_27=-0.0010852
+  sky130_fd_pr__pfet_01v8__cgidl_diff_27=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_27=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_27=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_27=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 028, W = 7.0, L = 2.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__kt1_diff_28=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_28=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_28=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_28=-5.2778e-11
+  sky130_fd_pr__pfet_01v8__b1_diff_28=0.0
+  sky130_fd_pr__pfet_01v8__bgidl_diff_28=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_28=0.0037674
+  sky130_fd_pr__pfet_01v8__ua_diff_28=-7.2465e-12
+  sky130_fd_pr__pfet_01v8__tvoff_diff_28=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_28=0.057603
+  sky130_fd_pr__pfet_01v8__ub_diff_28=2.958e-19
+  sky130_fd_pr__pfet_01v8__k2_diff_28=-0.012893
+  sky130_fd_pr__pfet_01v8__pdits_diff_28=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_28=-0.043436
+  sky130_fd_pr__pfet_01v8__eta0_diff_28=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_28=-0.066312
+  sky130_fd_pr__pfet_01v8__pditsd_diff_28=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_28=0.0014118
+  sky130_fd_pr__pfet_01v8__vsat_diff_28=0.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_28=0.0035519
+  sky130_fd_pr__pfet_01v8__cgidl_diff_28=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_28=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_28=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 029, W = 7.0, L = 4.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__rdsw_diff_29=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_29=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_29=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_29=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_29=-9.8052e-11
+  sky130_fd_pr__pfet_01v8__b1_diff_29=0.0
+  sky130_fd_pr__pfet_01v8__bgidl_diff_29=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_29=0.06067
+  sky130_fd_pr__pfet_01v8__ua_diff_29=-3.5733e-12
+  sky130_fd_pr__pfet_01v8__tvoff_diff_29=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_29=0.015944
+  sky130_fd_pr__pfet_01v8__ub_diff_29=3.6594e-19
+  sky130_fd_pr__pfet_01v8__k2_diff_29=-0.012367
+  sky130_fd_pr__pfet_01v8__pdits_diff_29=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_29=-0.045297
+  sky130_fd_pr__pfet_01v8__eta0_diff_29=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_29=-0.019005
+  sky130_fd_pr__pfet_01v8__pditsd_diff_29=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_29=0.0018876
+  sky130_fd_pr__pfet_01v8__vsat_diff_29=0.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_29=0.0008059
+  sky130_fd_pr__pfet_01v8__cgidl_diff_29=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_29=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 030, W = 7.0, L = 8.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__cgidl_diff_30=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_30=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_30=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_30=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_30=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_30=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_30=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_30=2.2358e-10
+  sky130_fd_pr__pfet_01v8__ua_diff_30=-5.0977e-12
+  sky130_fd_pr__pfet_01v8__bgidl_diff_30=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_30=0.093465
+  sky130_fd_pr__pfet_01v8__ub_diff_30=3.9461e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_30=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_30=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_30=-0.014315
+  sky130_fd_pr__pfet_01v8__k2_diff_30=-0.01321
+  sky130_fd_pr__pfet_01v8__voff_diff_30=-0.050926
+  sky130_fd_pr__pfet_01v8__a0_diff_30=0.016661
+  sky130_fd_pr__pfet_01v8__pditsd_diff_30=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_30=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_30=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_30=0.0020368
+  sky130_fd_pr__pfet_01v8__vth0_diff_30=-0.00026087
*
* sky130_fd_pr__pfet_01v8, Bin 031, W = 7.0, L = 0.15
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__u0_diff_31=0.00035699
+  sky130_fd_pr__pfet_01v8__vth0_diff_31=-0.026135
+  sky130_fd_pr__pfet_01v8__cgidl_diff_31=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_31=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_31=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_31=0.11383
+  sky130_fd_pr__pfet_01v8__pclm_diff_31=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_31=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_31=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_31=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_31=-3.5805e-12
+  sky130_fd_pr__pfet_01v8__bgidl_diff_31=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_31=0.015375
+  sky130_fd_pr__pfet_01v8__ub_diff_31=1.4685e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_31=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_31=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_31=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_31=-0.017121
+  sky130_fd_pr__pfet_01v8__voff_diff_31=-0.0079983
+  sky130_fd_pr__pfet_01v8__a0_diff_31=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_31=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_31=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_31=-4862.4
*
* sky130_fd_pr__pfet_01v8, Bin 032, W = 7.0, L = 0.18
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__pditsd_diff_32=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_32=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_32=8450.8
+  sky130_fd_pr__pfet_01v8__u0_diff_32=0.00050802
+  sky130_fd_pr__pfet_01v8__vth0_diff_32=-0.014432
+  sky130_fd_pr__pfet_01v8__cgidl_diff_32=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_32=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_32=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_32=-0.23267
+  sky130_fd_pr__pfet_01v8__pclm_diff_32=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_32=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_32=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_32=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_32=4.8344e-12
+  sky130_fd_pr__pfet_01v8__bgidl_diff_32=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_32=0.11128
+  sky130_fd_pr__pfet_01v8__ub_diff_32=1.885e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_32=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_32=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_32=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_32=-0.014444
+  sky130_fd_pr__pfet_01v8__voff_diff_32=-0.031532
+  sky130_fd_pr__pfet_01v8__a0_diff_32=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 033, W = 7.0, L = 0.25
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__voff_diff_33=-0.041527
+  sky130_fd_pr__pfet_01v8__a0_diff_33=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_33=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_33=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_33=11762.0
+  sky130_fd_pr__pfet_01v8__u0_diff_33=0.00061074
+  sky130_fd_pr__pfet_01v8__vth0_diff_33=-0.023852
+  sky130_fd_pr__pfet_01v8__cgidl_diff_33=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_33=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_33=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_33=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_33=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_33=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_33=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_33=1.8875e-10
+  sky130_fd_pr__pfet_01v8__ua_diff_33=8.1783e-12
+  sky130_fd_pr__pfet_01v8__bgidl_diff_33=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_33=0.10437
+  sky130_fd_pr__pfet_01v8__ub_diff_33=2.2026e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_33=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_33=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_33=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_33=-0.010822
*
* sky130_fd_pr__pfet_01v8, Bin 034, W = 7.0, L = 0.5
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__pdits_diff_34=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_34=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_34=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_34=-0.016
+  sky130_fd_pr__pfet_01v8__voff_diff_34=-0.057579
+  sky130_fd_pr__pfet_01v8__a0_diff_34=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_34=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_34=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_34=2997.3
+  sky130_fd_pr__pfet_01v8__u0_diff_34=0.0013699
+  sky130_fd_pr__pfet_01v8__vth0_diff_34=-0.0020141
+  sky130_fd_pr__pfet_01v8__cgidl_diff_34=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_34=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_34=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_34=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_34=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_34=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_34=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_34=-8.2093e-11
+  sky130_fd_pr__pfet_01v8__ua_diff_34=1.2152e-11
+  sky130_fd_pr__pfet_01v8__bgidl_diff_34=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_34=0.27919
+  sky130_fd_pr__pfet_01v8__ub_diff_34=2.8017e-19
*
* sky130_fd_pr__pfet_01v8, Bin 035, W = 0.42, L = 1.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__bgidl_diff_35=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_35=0.23441
+  sky130_fd_pr__pfet_01v8__ub_diff_35=3.3494e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_35=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_35=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_35=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_35=-0.0066897
+  sky130_fd_pr__pfet_01v8__voff_diff_35=-0.095705
+  sky130_fd_pr__pfet_01v8__a0_diff_35=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_35=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_35=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_35=0.0017171
+  sky130_fd_pr__pfet_01v8__vsat_diff_35=0.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_35=-0.031999
+  sky130_fd_pr__pfet_01v8__cgidl_diff_35=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_35=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_35=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_35=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_35=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_35=-4.0351e-9
+  sky130_fd_pr__pfet_01v8__b1_diff_35=-3.6399e-7
+  sky130_fd_pr__pfet_01v8__agidl_diff_35=-1.2307e-9
+  sky130_fd_pr__pfet_01v8__ua_diff_35=-8.8177e-12
*
* sky130_fd_pr__pfet_01v8, Bin 036, W = 0.42, L = 20.0
* -----------------------------------
+  sky130_fd_pr__pfet_01v8__agidl_diff_36=-2.4469e-10
+  sky130_fd_pr__pfet_01v8__b1_diff_36=1.6835e-11
+  sky130_fd_pr__pfet_01v8__ua_diff_36=-4.9955e-12
+  sky130_fd_pr__pfet_01v8__bgidl_diff_36=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_36=0.029222
+  sky130_fd_pr__pfet_01v8__ub_diff_36=7.6707e-21
+  sky130_fd_pr__pfet_01v8__pdits_diff_36=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_36=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_36=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_36=0.006486
+  sky130_fd_pr__pfet_01v8__voff_diff_36=-0.030456
+  sky130_fd_pr__pfet_01v8__eta0_diff_36=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_36=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_36=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_36=6.8715e-5
+  sky130_fd_pr__pfet_01v8__vsat_diff_36=20004.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_36=0.006343
+  sky130_fd_pr__pfet_01v8__cgidl_diff_36=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_36=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_36=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_36=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_36=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_36=-7.1468e-8
*
* sky130_fd_pr__pfet_01v8, Bin 037, W = 0.42, L = 2.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__b0_diff_37=3.6196e-9
+  sky130_fd_pr__pfet_01v8__agidl_diff_37=-2.9644e-10
+  sky130_fd_pr__pfet_01v8__b1_diff_37=2.639e-11
+  sky130_fd_pr__pfet_01v8__ua_diff_37=-4.996e-12
+  sky130_fd_pr__pfet_01v8__bgidl_diff_37=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_37=0.051268
+  sky130_fd_pr__pfet_01v8__ub_diff_37=-7.0453e-20
+  sky130_fd_pr__pfet_01v8__tvoff_diff_37=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_37=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_37=0.0031615
+  sky130_fd_pr__pfet_01v8__pdits_diff_37=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_37=-0.037179
+  sky130_fd_pr__pfet_01v8__eta0_diff_37=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_37=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_37=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_37=-0.00050532
+  sky130_fd_pr__pfet_01v8__vsat_diff_37=0.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_37=0.030585
+  sky130_fd_pr__pfet_01v8__cgidl_diff_37=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_37=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_37=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_37=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_37=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 038, W = 0.42, L = 4.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__pclm_diff_38=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_38=-3.5789e-8
+  sky130_fd_pr__pfet_01v8__agidl_diff_38=-6.3848e-10
+  sky130_fd_pr__pfet_01v8__b1_diff_38=4.0747e-7
+  sky130_fd_pr__pfet_01v8__ua_diff_38=-4.9282e-12
+  sky130_fd_pr__pfet_01v8__bgidl_diff_38=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_38=0.04431
+  sky130_fd_pr__pfet_01v8__tvoff_diff_38=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_38=0.0
+  sky130_fd_pr__pfet_01v8__ub_diff_38=1.428e-20
+  sky130_fd_pr__pfet_01v8__k2_diff_38=-0.001698
+  sky130_fd_pr__pfet_01v8__pdits_diff_38=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_38=-0.036994
+  sky130_fd_pr__pfet_01v8__eta0_diff_38=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_38=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_38=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_38=0.00036625
+  sky130_fd_pr__pfet_01v8__vsat_diff_38=0.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_38=0.0054604
+  sky130_fd_pr__pfet_01v8__cgidl_diff_38=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_38=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_38=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_38=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 039, W = 0.42, L = 8.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__kt1_diff_39=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_39=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_39=7.2037e-8
+  sky130_fd_pr__pfet_01v8__agidl_diff_39=-5.8047e-10
+  sky130_fd_pr__pfet_01v8__b1_diff_39=3.5899e-7
+  sky130_fd_pr__pfet_01v8__bgidl_diff_39=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_39=0.01066
+  sky130_fd_pr__pfet_01v8__ua_diff_39=-7.1907e-12
+  sky130_fd_pr__pfet_01v8__tvoff_diff_39=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_39=0.0
+  sky130_fd_pr__pfet_01v8__ub_diff_39=1.4267e-20
+  sky130_fd_pr__pfet_01v8__k2_diff_39=0.0016675
+  sky130_fd_pr__pfet_01v8__pdits_diff_39=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_39=-0.030352
+  sky130_fd_pr__pfet_01v8__eta0_diff_39=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_39=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_39=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_39=0.00022081
+  sky130_fd_pr__pfet_01v8__vsat_diff_39=20019.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_39=0.00966
+  sky130_fd_pr__pfet_01v8__cgidl_diff_39=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_39=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_39=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 040, W = 0.42, L = 0.15
* -----------------------------------
+  sky130_fd_pr__pfet_01v8__rdsw_diff_40=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_40=-0.26384
+  sky130_fd_pr__pfet_01v8__pclm_diff_40=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_40=-5.0608e-8
+  sky130_fd_pr__pfet_01v8__b1_diff_40=2.6414e-9
+  sky130_fd_pr__pfet_01v8__agidl_diff_40=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_40=-2.7512e-11
+  sky130_fd_pr__pfet_01v8__bgidl_diff_40=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_40=0.51388
+  sky130_fd_pr__pfet_01v8__ub_diff_40=2.1195e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_40=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_40=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_40=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_40=-0.030116
+  sky130_fd_pr__pfet_01v8__voff_diff_40=-0.1488
+  sky130_fd_pr__pfet_01v8__a0_diff_40=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_40=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_40=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_40=18914.0
+  sky130_fd_pr__pfet_01v8__u0_diff_40=0.00033774
+  sky130_fd_pr__pfet_01v8__vth0_diff_40=0.022711
+  sky130_fd_pr__pfet_01v8__cgidl_diff_40=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_40=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 041, W = 0.42, L = 0.18
* -----------------------------------
+  sky130_fd_pr__pfet_01v8__cgidl_diff_41=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_41=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_41=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_41=-0.36529
+  sky130_fd_pr__pfet_01v8__pclm_diff_41=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_41=-7.5986e-8
+  sky130_fd_pr__pfet_01v8__b1_diff_41=7.2273e-9
+  sky130_fd_pr__pfet_01v8__agidl_diff_41=-4.3892e-9
+  sky130_fd_pr__pfet_01v8__ua_diff_41=-2.732e-11
+  sky130_fd_pr__pfet_01v8__bgidl_diff_41=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_41=-0.48975
+  sky130_fd_pr__pfet_01v8__ub_diff_41=2.7027e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_41=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_41=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_41=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_41=-0.023178
+  sky130_fd_pr__pfet_01v8__voff_diff_41=-0.26953
+  sky130_fd_pr__pfet_01v8__a0_diff_41=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_41=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_41=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_41=18122.0
+  sky130_fd_pr__pfet_01v8__u0_diff_41=0.00049173
+  sky130_fd_pr__pfet_01v8__vth0_diff_41=0.040895
*
* sky130_fd_pr__pfet_01v8, Bin 042, W = 0.42, L = 0.5
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__u0_diff_42=0.0011702
+  sky130_fd_pr__pfet_01v8__vth0_diff_42=-0.017558
+  sky130_fd_pr__pfet_01v8__cgidl_diff_42=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_42=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_42=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_42=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_42=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_42=-4.3583e-8
+  sky130_fd_pr__pfet_01v8__b1_diff_42=4.4592e-9
+  sky130_fd_pr__pfet_01v8__agidl_diff_42=-4.7051e-10
+  sky130_fd_pr__pfet_01v8__ua_diff_42=-1.505e-11
+  sky130_fd_pr__pfet_01v8__bgidl_diff_42=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_42=0.14181
+  sky130_fd_pr__pfet_01v8__ub_diff_42=2.7814e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_42=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_42=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_42=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_42=-0.0065428
+  sky130_fd_pr__pfet_01v8__voff_diff_42=-0.089
+  sky130_fd_pr__pfet_01v8__a0_diff_42=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_42=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_42=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_42=20455.0
*
* sky130_fd_pr__pfet_01v8, Bin 043, W = 0.55, L = 1.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__pditsd_diff_43=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_43=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_43=20224.0
+  sky130_fd_pr__pfet_01v8__u0_diff_43=0.0011785
+  sky130_fd_pr__pfet_01v8__vth0_diff_43=-0.038892
+  sky130_fd_pr__pfet_01v8__cgidl_diff_43=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_43=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_43=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_43=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_43=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_43=-3.9601e-8
+  sky130_fd_pr__pfet_01v8__b1_diff_43=7.0785e-9
+  sky130_fd_pr__pfet_01v8__agidl_diff_43=-4.7279e-10
+  sky130_fd_pr__pfet_01v8__ua_diff_43=-3.0087e-11
+  sky130_fd_pr__pfet_01v8__bgidl_diff_43=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_43=0.14077
+  sky130_fd_pr__pfet_01v8__ub_diff_43=2.7797e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_43=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_43=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_43=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_43=-0.01132
+  sky130_fd_pr__pfet_01v8__voff_diff_43=-0.083804
+  sky130_fd_pr__pfet_01v8__a0_diff_43=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 044, W = 0.55, L = 2.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__voff_diff_44=-0.071307
+  sky130_fd_pr__pfet_01v8__a0_diff_44=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_44=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_44=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_44=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_44=0.0017219
+  sky130_fd_pr__pfet_01v8__vth0_diff_44=0.0005957
+  sky130_fd_pr__pfet_01v8__cgidl_diff_44=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_44=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_44=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_44=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_44=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_44=-7.8126e-8
+  sky130_fd_pr__pfet_01v8__b1_diff_44=2.4927e-8
+  sky130_fd_pr__pfet_01v8__agidl_diff_44=-1.7503e-10
+  sky130_fd_pr__pfet_01v8__ua_diff_44=-1.7426e-12
+  sky130_fd_pr__pfet_01v8__bgidl_diff_44=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_44=0.10072
+  sky130_fd_pr__pfet_01v8__ub_diff_44=3.4467e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_44=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_44=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_44=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_44=-0.0083627
*
* sky130_fd_pr__pfet_01v8, Bin 045, W = 0.55, L = 4.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__pdits_diff_45=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_45=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_45=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_45=0.00078773
+  sky130_fd_pr__pfet_01v8__voff_diff_45=-0.035423
+  sky130_fd_pr__pfet_01v8__a0_diff_45=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_45=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_45=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_45=20043.0
+  sky130_fd_pr__pfet_01v8__u0_diff_45=-1.4763e-5
+  sky130_fd_pr__pfet_01v8__vth0_diff_45=0.013746
+  sky130_fd_pr__pfet_01v8__cgidl_diff_45=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_45=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_45=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_45=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_45=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_45=2.3397e-8
+  sky130_fd_pr__pfet_01v8__b1_diff_45=1.2339e-8
+  sky130_fd_pr__pfet_01v8__agidl_diff_45=1.5067e-9
+  sky130_fd_pr__pfet_01v8__ua_diff_45=-4.8743e-12
+  sky130_fd_pr__pfet_01v8__bgidl_diff_45=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_45=0.029362
+  sky130_fd_pr__pfet_01v8__ub_diff_45=-1.3062e-20
*
* sky130_fd_pr__pfet_01v8, Bin 046, W = 0.55, L = 8.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__bgidl_diff_46=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_46=0.1837
+  sky130_fd_pr__pfet_01v8__ub_diff_46=3.1309e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_46=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_46=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_46=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_46=-0.011371
+  sky130_fd_pr__pfet_01v8__voff_diff_46=-0.082567
+  sky130_fd_pr__pfet_01v8__a0_diff_46=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_46=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_46=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_46=0.0016571
+  sky130_fd_pr__pfet_01v8__vsat_diff_46=0.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_46=-0.021094
+  sky130_fd_pr__pfet_01v8__cgidl_diff_46=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_46=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_46=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_46=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_46=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_46=-1.1444e-7
+  sky130_fd_pr__pfet_01v8__b1_diff_46=2.7921e-7
+  sky130_fd_pr__pfet_01v8__agidl_diff_46=-9.8638e-10
+  sky130_fd_pr__pfet_01v8__ua_diff_46=-7.5875e-12
*
* sky130_fd_pr__pfet_01v8, Bin 047, W = 0.55, L = 0.15
* -----------------------------------
+  sky130_fd_pr__pfet_01v8__agidl_diff_47=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_47=2.5223e-9
+  sky130_fd_pr__pfet_01v8__ua_diff_47=-2.3128e-11
+  sky130_fd_pr__pfet_01v8__bgidl_diff_47=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_47=0.45086
+  sky130_fd_pr__pfet_01v8__ub_diff_47=2.367e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_47=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_47=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_47=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_47=-0.024865
+  sky130_fd_pr__pfet_01v8__voff_diff_47=-0.12465
+  sky130_fd_pr__pfet_01v8__eta0_diff_47=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_47=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_47=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_47=0.00026223
+  sky130_fd_pr__pfet_01v8__vsat_diff_47=19667.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_47=0.030658
+  sky130_fd_pr__pfet_01v8__cgidl_diff_47=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_47=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_47=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_47=-0.079642
+  sky130_fd_pr__pfet_01v8__pclm_diff_47=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_47=2.6947e-8
*
* sky130_fd_pr__pfet_01v8, Bin 048, W = 0.55, L = 0.5
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__b0_diff_48=-6.8221e-8
+  sky130_fd_pr__pfet_01v8__agidl_diff_48=-1.713e-10
+  sky130_fd_pr__pfet_01v8__b1_diff_48=3.3139e-10
+  sky130_fd_pr__pfet_01v8__ua_diff_48=-1.2629e-11
+  sky130_fd_pr__pfet_01v8__bgidl_diff_48=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_48=0.10376
+  sky130_fd_pr__pfet_01v8__ub_diff_48=2.9391e-19
+  sky130_fd_pr__pfet_01v8__tvoff_diff_48=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_48=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_48=-0.018886
+  sky130_fd_pr__pfet_01v8__pdits_diff_48=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_48=-0.080025
+  sky130_fd_pr__pfet_01v8__eta0_diff_48=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_48=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_48=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_48=0.0011564
+  sky130_fd_pr__pfet_01v8__vsat_diff_48=20219.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_48=-0.0020992
+  sky130_fd_pr__pfet_01v8__cgidl_diff_48=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_48=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_48=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_48=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_48=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 049, W = 0.64, L = 0.15
* -----------------------------------
+  sky130_fd_pr__pfet_01v8__pclm_diff_49=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_49=1.3673e-7
+  sky130_fd_pr__pfet_01v8__agidl_diff_49=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_49=6.4955e-10
+  sky130_fd_pr__pfet_01v8__ua_diff_49=-1.2078e-10
+  sky130_fd_pr__pfet_01v8__bgidl_diff_49=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_49=-1.0761
+  sky130_fd_pr__pfet_01v8__tvoff_diff_49=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_49=0.0
+  sky130_fd_pr__pfet_01v8__ub_diff_49=2.2638e-19
+  sky130_fd_pr__pfet_01v8__k2_diff_49=-0.013115
+  sky130_fd_pr__pfet_01v8__pdits_diff_49=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_49=0.10157
+  sky130_fd_pr__pfet_01v8__eta0_diff_49=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_49=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_49=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_49=2.9246e-5
+  sky130_fd_pr__pfet_01v8__vsat_diff_49=21326.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_49=-0.044111
+  sky130_fd_pr__pfet_01v8__cgidl_diff_49=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_49=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_49=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_49=-0.030294
*
* sky130_fd_pr__pfet_01v8, Bin 050, W = 0.84, L = 0.15
* -----------------------------------
+  sky130_fd_pr__pfet_01v8__kt1_diff_50=0.1034
+  sky130_fd_pr__pfet_01v8__pclm_diff_50=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_50=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_50=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_50=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_50=-2.4518e-11
+  sky130_fd_pr__pfet_01v8__bgidl_diff_50=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_50=-0.61881
+  sky130_fd_pr__pfet_01v8__ub_diff_50=2.7121e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_50=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_50=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_50=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_50=-0.040295
+  sky130_fd_pr__pfet_01v8__voff_diff_50=0.094422
+  sky130_fd_pr__pfet_01v8__a0_diff_50=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_50=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_50=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_50=-198.03
+  sky130_fd_pr__pfet_01v8__u0_diff_50=0.00057136
+  sky130_fd_pr__pfet_01v8__vth0_diff_50=-0.040605
+  sky130_fd_pr__pfet_01v8__cgidl_diff_50=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_50=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_50=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 051, W = 1.65, L = 0.15
* -----------------------------------
+  sky130_fd_pr__pfet_01v8__rdsw_diff_51=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_51=0.099002
+  sky130_fd_pr__pfet_01v8__pclm_diff_51=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_51=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_51=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_51=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_51=-6.7472e-12
+  sky130_fd_pr__pfet_01v8__bgidl_diff_51=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_51=0.018346
+  sky130_fd_pr__pfet_01v8__ub_diff_51=2.3163e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_51=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_51=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_51=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_51=-0.030703
+  sky130_fd_pr__pfet_01v8__voff_diff_51=-0.0028909
+  sky130_fd_pr__pfet_01v8__a0_diff_51=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_51=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_51=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_51=2274.8
+  sky130_fd_pr__pfet_01v8__u0_diff_51=0.00055896
+  sky130_fd_pr__pfet_01v8__vth0_diff_51=0.0021626
+  sky130_fd_pr__pfet_01v8__cgidl_diff_51=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_51=0.0
.include "sky130_fd_pr__pfet_01v8.pm3.spice"
