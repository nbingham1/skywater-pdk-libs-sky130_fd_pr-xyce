* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre=0.0
* statistics {
*   process {
*   }
*   mismatch {
*     vary sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre dist=gauss std = 1.0
*   }
* }
.subckt sky130_fd_pr__nfet_g5v0d10v5 d g s b
.param l=1 w=1 ad=0 as=0 pd=0 ps=0 nrd=0 nrs=0 sa=0 sb=0 sd=0 mult=1 nf=1.0
msky130_fd_pr__nfet_g5v0d10v5 d g s b sky130_fd_pr__nfet_g5v0d10v5__model l={l} w={w} ad={ad} as={as} pd={pd} ps={ps} nrd={nrd} nrs={nrs} sa={sa} sb={sb} sd={sd} nf={nf}
.model sky130_fd_pr__nfet_g5v0d10v5__model.0 nmos
* DC IV MOS Parameters
+  lmin=2.0e-05 lmax=1.0e-04 wmin=2.0e-05 wmax=1.0e-4
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.791968+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+  k1=0.88325
+  k2=-0.0388233
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=105660.0
+  ua=-6.02229e-11
+  ub=1.73106e-18
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0426101
+  a0=0.9440931
+  keta=-0.02132
+  a1=0.0
+  a2=0.65972622
+  ags=0.1460627
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.93087+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.33405
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.4467e-5
+  alpha1=0.0
+  beta0=24.0
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.40273
+  kt2=-0.019151
+  at=160000.0
+  ute=-1.2986
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.1 nmos
* DC IV MOS Parameters
+  lmin=8e-06 lmax=2.0e-05 wmin=2.0e-05 wmax=1.0e-4
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.791968+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+  k1=0.88325
+  k2=-0.0388233
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=105660.0
+  ua=-6.02229e-11
+  ub=1.73106e-18
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0426101
+  a0=0.9440931
+  keta=-0.02132
+  a1=0.0
+  a2=0.65972622
+  ags=0.1460627
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.93087+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.33405
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.4467e-5
+  alpha1=0.0
+  beta0=24.0
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.40273
+  kt2=-0.019151
+  at=160000.0
+  ute=-1.2986
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.2 nmos
* DC IV MOS Parameters
+  lmin=4e-06 lmax=8e-06 wmin=2.0e-05 wmax=1.0e-4
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.787009917893+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=3.87857425989731e-8
+  k1=0.88325
+  k2=-0.040038259480075 lk2=9.50430118852657e-09 wk2=-2.11758236813575e-22
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=110438.41375 lvsat=-0.0373802453729513
+  ua=-1.026911477714e-10 lua=3.32217678357012e-16
+  ub=1.872940661065e-18 lub=-1.10989424561367e-24
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0426265377433 lu0=-1.28588044082879e-10
+  a0=1.03171951755192 la0=-6.85477893002309e-7
+  keta=-0.01729370857425 lketa=-3.14965947512488e-8
+  a1=0.0
+  a2=0.65972622
+  ags=0.158828805742775 lags=-9.98658111432839e-8
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.9704065953675+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-3.09284150215799e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.2603764168025 lpclm=5.76328623160162e-7
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.4467e-5
+  alpha1=0.0
+  beta0=21.51522485 lbeta0=1.94377275939346e-5
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.414198193 lkt1=8.97125888950827e-8
+  kt2=-0.019151
+  at=236454.62 lat=-0.59808392596722
+  ute=-1.33682731 lute=2.9904196298361e-7
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.3 nmos
* DC IV MOS Parameters
+  lmin=2e-06 lmax=4e-06 wmin=2.0e-05 wmax=1.0e-4
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.803592063161+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-2.46033381635131e-8
+  k1=0.88325
+  k2=-0.04195453332085 lk2=1.68297006041463e-8
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=93870.327025 lvsat=0.0259550933613947
+  ua=1.037893167889e-10 lua=-4.57101594412049e-16 wua=1.97215226305253e-31
+  ub=1.535692017715e-18 lub=1.79316598028321e-25
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.04299289831795 lu0=-1.52908596997534e-9
+  a0=0.484478507841295 la0=1.40647727928978e-6
+  keta=-0.0390877390815 lketa=5.18161212837616e-8
+  a1=0.0
+  a2=0.65972622
+  ags=0.1175536953818 lags=5.79178327620362e-8
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.93082131177+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.57960259463844e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.598489405835 lpclm=-7.16186381517036e-7
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.4467e-5
+  alpha1=0.0
+  beta0=23.895067196 lbeta0=1.03402304827677e-5
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.407134579 lkt1=6.27102926852489e-8
+  kt2=-0.019151
+  at=138327.392 lat=-0.222969929547552 pat=8.470329472543e-22
+  ute=-1.22214538 lute=-1.39356205967221e-7
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.4 nmos
* DC IV MOS Parameters
+  lmin=1e-06 lmax=2e-06 wmin=2.0e-05 wmax=1.0e-4
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.785561574921+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=8.26139169667085e-9
+  k1=0.88325
+  k2=-0.0399663514591 lk2=1.32057798910968e-8
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=119548.429093 lvsat=-0.020849179299113
+  ua=-1.434293897823e-10 lua=-6.48839416481854e-18
+  ub=1.73676328342e-18 lub=-1.8718223118142e-25
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.04062432093363 lu0=2.78819345432367e-9
+  a0=1.66774023460685 la0=-7.50290551199328e-7
+  keta=0.00292164334800001 lketa=-2.47556823613434e-8
+  a1=0.0
+  a2=0.65972622
+  ags=0.169635646542 lags=-3.70135541581461e-8
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.90016329917+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.02078949499433e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.0998655211199999 lpclm=1.92670830493421e-7
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.4467e-5
+  alpha1=0.0
+  beta0=27.155752708 lbeta0=4.39687791879445e-6
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.38095731 lkt1=1.49961729836101e-8
+  kt2=-0.019151
+  at=9418.15199999999 lat=0.011996938386888
+  ute=-1.2986
+  ua1=3.0044e-9
+  ub1=-3.9994838462e-18 lub1=4.50185112967972e-25
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.81e-6
+  sbref=2.81e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.5 nmos
* DC IV MOS Parameters
+  lmin=8.0e-07 lmax=1e-06 wmin=2.0e-05 wmax=1.0e-4
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.797997400694999+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-1.96994767819776e-9
+  k1=0.88325
+  k2=-0.035281286212 lk2=9.35123147528498e-9
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=101453.720647 lvsat=-0.00596210172462697
+  ua=-1.5625551402054e-10 lua=4.0640558558329e-18
+  ub=8.1144877795e-19 lub=5.74102697218418e-25
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.04542553049835 lu0=-1.161910492068e-9
+  a0=-0.385088442204999 la0=9.38635238902762e-7
+  keta=-0.07856821674 lketa=4.22885517187169e-8
+  a1=0.0
+  a2=0.65972622
+  ags=0.013791541035 lags=9.12042226097334e-8
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.7564739735+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.61387130983717e-8
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-1.82604815625 lpclm=1.77717971618972e-6
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=5.45919608500001e-06 lalpha0=7.41099952279187e-12
+  alpha1=0.0
+  beta0=23.21508079 lbeta0=7.63899086656252e-6
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.33782076 lkt1=-2.049360393444e-8
+  kt2=-0.019151
+  at=8431.72499999999 lat=0.012808502459025
+  ute=-1.4589532325 lute=1.31927575327957e-7
+  ua1=6.0953253185e-09 lua1=-2.54300007821482e-15
+  ub1=-9.6961123715e-18 lub1=5.13697799621657e-24
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.41e-6
+  sbref=2.41e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.6 nmos
* DC IV MOS Parameters
+  lmin=6e-07 lmax=8.0e-07 wmin=2.0e-05 wmax=1.0e-4
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.788372556665+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=4.02374106944794e-9
+  k1=0.88325
+  k2=-0.0083448426275 lk2=-7.4229269745343e-9
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=77796.1053695001 lvsat=0.00877022869474586
+  ua=-2.8572090550946e-10 lua=8.46861685631196e-17 wua=-1.57772181044202e-30
+  ub=1.0505226157e-18 lub=4.25224007162524e-25
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0362910518205 lu0=4.5264125494682e-9
+  a0=1.1222
+  keta=-0.01066
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.75091767705+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.95987911429766e-8
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=1.031604579 lpclm=-2.36922928524898e-9
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.674704005e-05 lalpha0=3.81709162623447e-13
+  alpha1=0.0
+  beta0=32.35801791 lbeta0=1.9454004908878e-6
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.37073
+  kt2=-0.019151
+  at=9131.64300000003 lat=0.012372641822967
+  ute=-1.13718994 lute=-6.84444015738598e-8
+  ua1=2.0117e-9
+  ub1=-1.6583655e-18 lub1=1.316238491805e-25
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.02e-6
+  sbref=2.01e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.7 nmos
* DC IV MOS Parameters
+  lmin=5e-07 lmax=6e-07 wmin=2.0e-05 wmax=1.0e-4
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.95843676326+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-6.78676710486631e-8
+  k1=0.88325
+  k2=0.00538350225699999 lk2=-1.32263239359039e-8
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=105285.196052 lvsat=-0.00285026209855802
+  ua=1.33486686931e-10 lua=-9.25258761968286e-17
+  ub=5.2928310142e-18 lub=-1.36813126444378e-24
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0504624395499 lu0=-1.46427235676878e-9
+  a0=1.1222
+  keta=-0.01066
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.649678730855+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-3.60335367893065e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.190772172 lpclm=3.53076694958268e-7
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=2.792252773e-05 lalpha0=-4.34251591983063e-12
+  alpha1=0.0
+  beta0=36.96
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.4352762 lkt1=2.72856796722001e-8
+  kt2=-0.019151
+  at=2254.128 lat=0.015279980616432
+  ute=-1.300713655 lute=6.82141991805027e-10
+  ua1=-1.192050637e-09 lua1=1.35432471052965e-15
+  ub1=5.286735705e-18 lub1=-2.80428572831036e-24 pub1=5.60519385729927e-45
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=1.81e-6
+  sbref=1.81e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.8 nmos
* DC IV MOS Parameters
+  lmin=2.0e-05 lmax=1.0e-04 wmin=1.5e-05 wmax=2.0e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.791968+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+  k1=0.88325
+  k2=-0.0388233
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=105660.0
+  ua=-6.02229e-11
+  ub=1.73106e-18
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0426101
+  a0=0.9440931
+  keta=-0.02132
+  a1=0.0
+  a2=0.65972622
+  ags=0.1460627
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.93087+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.33405
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.4467e-5
+  alpha1=0.0
+  beta0=24.0
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.40273
+  kt2=-0.019151
+  at=160000.0
+  ute=-1.2986
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.9 nmos
* DC IV MOS Parameters
+  lmin=8e-06 lmax=2.0e-05 wmin=1.5e-05 wmax=2.0e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.791968+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+  k1=0.88325
+  k2=-0.0388233
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=105660.0
+  ua=-6.02229e-11
+  ub=1.73106e-18
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0426101
+  a0=0.9440931
+  keta=-0.02132
+  a1=0.0
+  a2=0.65972622
+  ags=0.1460627
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.93087+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.33405
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.4467e-5
+  alpha1=0.0
+  beta0=24.0
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.40273
+  kt2=-0.019151
+  at=160000.0
+  ute=-1.2986
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.10 nmos
* DC IV MOS Parameters
+  lmin=4e-06 lmax=8e-06 wmin=1.5e-05 wmax=2.0e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.787009917893002+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=3.87857425989748e-8
+  k1=0.88325
+  k2=-0.040038259480075 lk2=9.50430118852636e-9
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=110438.41375 lvsat=-0.0373802453729506
+  ua=-1.026911477714e-10 lua=3.32217678357012e-16
+  ub=1.872940661065e-18 lub=-1.10989424561366e-24 wub=-2.35098870164458e-38
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0426265377433001 lu0=-1.28588044082931e-10
+  a0=1.03171951755192 la0=-6.85477893002309e-07 wa0=1.35525271560688e-20
+  keta=-0.01729370857425 lketa=-3.14965947512487e-8
+  a1=0.0
+  a2=0.65972622
+  ags=0.158828805742775 lags=-9.98658111432844e-8
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.970406595367501+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-3.09284150215798e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.2603764168025 lpclm=5.7632862316016e-7
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.4467e-5
+  alpha1=0.0
+  beta0=21.51522485 lbeta0=1.94377275939347e-5
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.414198193000001 lkt1=8.97125888950823e-8
+  kt2=-0.019151
+  at=236454.62 lat=-0.59808392596722
+  ute=-1.33682731 lute=2.9904196298361e-7
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.11 nmos
* DC IV MOS Parameters
+  lmin=2e-06 lmax=4e-06 wmin=1.5e-05 wmax=2.0e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.803592063160999+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-2.4603338163511e-8
+  k1=0.88325
+  k2=-0.04195453332085 lk2=1.68297006041463e-8
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=93870.3270250001 lvsat=0.0259550933613948
+  ua=1.037893167889e-10 lua=-4.57101594412049e-16 pua=3.00926553810506e-36
+  ub=1.535692017715e-18 lub=1.79316598028322e-25
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0429928983179501 lu0=-1.52908596997528e-9
+  a0=0.484478507841295 la0=1.40647727928978e-6
+  keta=-0.0390877390815 lketa=5.18161212837616e-8
+  a1=0.0
+  a2=0.65972622
+  ags=0.1175536953818 lags=5.79178327620359e-8
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.930821311770001+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.57960259463842e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.598489405835001 lpclm=-7.16186381517035e-7
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.4467e-5
+  alpha1=0.0
+  beta0=23.895067196 lbeta0=1.03402304827677e-5
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.407134579 lkt1=6.27102926852496e-8
+  kt2=-0.019151
+  at=138327.392 lat=-0.222969929547552
+  ute=-1.22214538 lute=-1.39356205967219e-7
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.12 nmos
* DC IV MOS Parameters
+  lmin=1e-06 lmax=2e-06 wmin=1.5e-05 wmax=2.0e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.785225848128792+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=8.8733313283599e-09 wvth0=6.71532413068488e-09 pvth0=-1.22402294680404e-14
+  k1=0.88325
+  k2=-0.038728112054894 lk2=1.09488025436291e-08 wk2=-2.47676954702401e-08 pk2=4.51448463321668e-14
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=126954.167156433 lvsat=-0.0343478476452119 wvsat=-0.148132149941629 pvsat=2.70005061795254e-7
+  ua=-1.54430860533465e-10 lua=1.35643276189229e-17 wua=2.20055246476621e-16 pua=-4.01101519465579e-22
+  ub=1.78692481590298e-18 lub=-2.78613211445664e-25 wub=-1.00334842893794e-24 pub=1.82883428522652e-30
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0397457041697843 lu0=4.38967546690488e-09 wu0=1.75743982690754e-08 pu0=-3.2033400531389e-14
+  a0=1.79236893189701 la0=-9.77455141239711e-07 wa0=-2.49286657398435e-06 pa0=4.54382518326508e-12
+  keta=0.00292164334800001 lketa=-2.47556823613434e-8
+  a1=0.0
+  a2=0.65972622
+  ags=-0.0474685019462415 lags=3.58708907519975e-07 wags=4.34259273030548e-06 pags=-7.91537838990244e-12
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.907149378743171+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.1481269330592e-07 wnfactor=-1.39737994778264e-07 pnfactor=2.54704774960184e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.0998655211200001 lpclm=1.92670830493421e-7
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.4467e-5
+  alpha1=0.0
+  beta0=27.2174671918619 lbeta0=4.28438901591029e-06 wbeta0=-1.23443458284684e-06 pbeta0=2.25004218162666e-12
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.38095731 lkt1=1.49961729836102e-8
+  kt2=-0.019151
+  at=9418.152 lat=0.011996938386888
+  ute=-1.2986
+  ua1=3.0044e-9
+  ub1=-3.9994838462e-18 lub1=4.50185112967973e-25
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.81e-6
+  sbref=2.81e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.13 nmos
* DC IV MOS Parameters
+  lmin=8.0e-07 lmax=1e-06 wmin=1.5e-05 wmax=2.0e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.799676034656045+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-3.01528508339302e-09 wvth0=-3.35766206534108e-08 pvth0=2.09092025561288e-14
+  k1=0.88325
+  k2=-0.0414724832330298 lk2=1.32066817873879e-08 wk2=1.23838477351202e-07 pk2=-7.7118058839391e-14
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=64425.0303298361 lvsat=0.0170968116252709 wvsat=0.740660749708145 pvsat=-4.61232409326504e-7
+  ua=-1.01248160264716e-10 lua=-3.01907285558855e-17 wua=-1.10027623238311e-15 pua=6.85176118468163e-22
+  ub=5.60641115535077e-19 lub=7.30288403641725e-25 wub=5.01674214468981e-24 pub=-3.12408085250485e-30
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0498186143175784 lu0=-3.89761997189992e-09 wu0=-8.78719913453745e-08 pu0=5.47206130424963e-14
+  a0=-1.00823192865578 la0=1.32668600536374e-06 wa0=1.24643328699218e-05 pa0=-7.76192647241927e-12
+  keta=-0.07856821674 lketa=4.22885517187169e-8
+  a1=0.0
+  a2=0.65972622
+  ags=1.09931228347621 lags=-5.84783194851422e-07 wags=-2.17129636515274e-05 pags=1.35213355676793e-11
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.721543575634142+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=3.78909546917761e-08 wnfactor=6.98689973891348e-07 pnfactor=-4.3509590613135e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-1.82604815625 lpclm=1.77717971618972e-6
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=5.45919608500002e-06 lalpha0=7.41099952279187e-12
+  alpha1=0.0
+  beta0=22.9065083706903 lbeta0=7.83114847781167e-06 wbeta0=6.17217291423375e-06 pbeta0=-3.84360341105397e-12
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.33782076 lkt1=-2.04936039344402e-8
+  kt2=-0.019151
+  at=8431.72499999998 lat=0.012808502459025
+  ute=-1.4589532325 lute=1.31927575327956e-7
+  ua1=6.0953253185e-09 lua1=-2.54300007821482e-15
+  ub1=-9.6961123715e-18 lub1=5.13697799621656e-24
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.41e-6
+  sbref=2.41e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.14 nmos
* DC IV MOS Parameters
+  lmin=6e-07 lmax=8.0e-07 wmin=1.5e-05 wmax=2.0e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.788372556664999+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=4.02374106944815e-9
+  k1=0.88325
+  k2=-0.00834484262750002 lk2=-7.4229269745343e-9
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=77796.1053695001 lvsat=0.00877022869474586
+  ua=-2.8572090550946e-10 lua=8.46861685631194e-17
+  ub=1.0505226157e-18 lub=4.25224007162523e-25
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0362910518205001 lu0=4.52641254946822e-9
+  a0=1.1222
+  keta=-0.01066
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.750917677050001+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.95987911429759e-8
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=1.031604579 lpclm=-2.36922928524962e-9
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.674704005e-05 lalpha0=3.81709162623451e-13
+  alpha1=0.0
+  beta0=32.3580179099999 lbeta0=1.94540049088779e-6
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.37073
+  kt2=-0.019151
+  at=9131.64299999998 lat=0.012372641822967
+  ute=-1.13718994 lute=-6.84444015738594e-8
+  ua1=2.0117e-9
+  ub1=-1.6583655e-18 lub1=1.316238491805e-25
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.02e-6
+  sbref=2.01e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.15 nmos
* DC IV MOS Parameters
+  lmin=5e-07 lmax=6e-07 wmin=1.5e-05 wmax=2.0e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={1.00533369003335+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-8.76924558004896e-08 wvth0=-9.38048649451055e-07 pvth0=3.96542243631109e-13
+  k1=0.88325
+  k2=0.0335303734220003 lk2=-2.51248789303556e-08 wk2=-5.63003512153503e-07 pk2=2.37999037696162e-13
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=158758.150694808 lvsat=-0.0254549376876666 wvsat=-1.06958464735365 pvsat=4.52146587560456e-7
+  ua=6.15764519709392e-11 lua=-6.21271906619271e-17 wua=1.4383735444329e-15 pua=-6.08045086811666e-22
+  ub=1.44757392587665e-17 lub=-5.25003124957763e-24 wub=-1.83679726359889e-22 pub=7.76471144038421e-29
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.070953481832745 lu0=-1.01264711520382e-08 wu0=-4.09868958624181e-07 pu0=1.73264314748159e-13
+  a0=1.1222
+  keta=-0.01066
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={2.32034932756341+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-6.4384861991021e-07 wnfactor=-1.34149866687293e-05 pnfactor=5.67093072945863e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-1.80014423200594 lpclm=1.1946987773401e-06 wpclm=3.98230027518355e-05 ppclm=-1.68344177762862e-11
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=2.792252773e-05 lalpha0=-4.34251591983064e-12
+  alpha1=0.0
+  beta0=36.96
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.435276200000001 lkt1=2.72856796722002e-8
+  kt2=-0.019151
+  at=-74593.6958433423 lat=0.0477659380375519 wat=1.53713691555723 pat=-6.49795425450424e-7
+  ute=-1.300713655 lute=6.82141991805451e-10
+  ua1=-1.192050637e-09 lua1=1.35432471052965e-15
+  ub1=1.89752976432841e-18 lub1=-1.37156331180431e-24 wub1=6.77920766689806e-23 pub1=-2.86578123623548e-29
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=1.81e-6
+  sbref=1.81e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.16 nmos
* DC IV MOS Parameters
+  lmin=2.0e-05 lmax=1.0e-04 wmin=1.0e-05 wmax=1.5e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.791968+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+  k1=0.88325
+  k2=-0.0388233
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=105660.0
+  ua=-6.02229e-11
+  ub=1.73106e-18
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0426101
+  a0=0.9440931
+  keta=-0.02132
+  a1=0.0
+  a2=0.65972622
+  ags=0.1460627
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.93087+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.33405
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.4467e-5
+  alpha1=0.0
+  beta0=24.0
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.40273
+  kt2=-0.019151
+  at=160000.0
+  ute=-1.2986
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.17 nmos
* DC IV MOS Parameters
+  lmin=8e-06 lmax=2.0e-05 wmin=1.0e-05 wmax=1.5e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.791968+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+  k1=0.88325
+  k2=-0.0388233
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=105660.0
+  ua=-6.02229e-11
+  ub=1.73106e-18
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0426101
+  a0=0.9440931
+  keta=-0.02132
+  a1=0.0
+  a2=0.65972622
+  ags=0.1460627
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.93087+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.33405
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.4467e-5
+  alpha1=0.0
+  beta0=24.0
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.40273
+  kt2=-0.019151
+  at=160000.0
+  ute=-1.2986
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.18 nmos
* DC IV MOS Parameters
+  lmin=4e-06 lmax=8e-06 wmin=1.0e-05 wmax=1.5e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.787009917893+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=3.87857425989748e-8
+  k1=0.88325
+  k2=-0.040038259480075 lk2=9.50430118852667e-9
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=110438.41375 lvsat=-0.0373802453729515
+  ua=-1.026911477714e-10 lua=3.32217678357012e-16
+  ub=1.872940661065e-18 lub=-1.10989424561367e-24
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0426265377433 lu0=-1.2858804408272e-10
+  a0=1.03171951755191 la0=-6.85477893002309e-7
+  keta=-0.01729370857425 lketa=-3.14965947512487e-8
+  a1=0.0
+  a2=0.65972622
+  ags=0.158828805742775 lags=-9.98658111432839e-8
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.9704065953675+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-3.09284150215798e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.2603764168025 lpclm=5.76328623160162e-7
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.4467e-5
+  alpha1=0.0
+  beta0=21.51522485 lbeta0=1.94377275939347e-5
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.414198193 lkt1=8.9712588895084e-8
+  kt2=-0.019151
+  at=236454.62 lat=-0.59808392596722
+  ute=-1.33682731 lute=2.99041962983613e-7
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.19 nmos
* DC IV MOS Parameters
+  lmin=2e-06 lmax=4e-06 wmin=1.0e-05 wmax=1.5e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.803592063161+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-2.4603338163511e-8
+  k1=0.88325
+  k2=-0.04195453332085 lk2=1.68297006041463e-8
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=93870.3270249999 lvsat=0.0259550933613948
+  ua=1.037893167889e-10 lua=-4.57101594412049e-16 wua=1.97215226305253e-31 pua=-9.4039548065783e-37
+  ub=1.535692017715e-18 lub=1.79316598028319e-25
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.04299289831795 lu0=-1.52908596997539e-9
+  a0=0.484478507841294 la0=1.40647727928978e-6
+  keta=-0.0390877390815 lketa=5.18161212837616e-8
+  a1=0.0
+  a2=0.65972622
+  ags=0.1175536953818 lags=5.79178327620362e-8
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.930821311769999+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.57960259463845e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.598489405835 lpclm=-7.16186381517035e-7
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.4467e-5
+  alpha1=0.0
+  beta0=23.895067196 lbeta0=1.03402304827677e-5
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.407134579 lkt1=6.27102926852487e-8
+  kt2=-0.019151
+  at=138327.392 lat=-0.222969929547552
+  ute=-1.22214538 lute=-1.3935620596722e-7
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.20 nmos
* DC IV MOS Parameters
+  lmin=1e-06 lmax=2e-06 wmin=1.0e-05 wmax=1.5e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.779911351247974+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=1.85602295424295e-08 wvth0=8.64452557816184e-08 pvth0=-1.57566447516098e-13
+  k1=0.88325
+  k2=-0.0394474831600657 lk2=1.22600225575297e-08 wk2=-1.39754398093107e-08 pk2=2.54734673790649e-14
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=124030.653693959 lvsat=-0.0290190690282435 wvsat=-0.10427258359491 pvsat=1.90060870568535e-7
+  ua=-1.27838964649181e-10 lua=-3.49055453581343e-17 wua=-1.78885629559177e-16 pua=3.26060382452032e-22
+  ub=1.90186225721914e-18 lub=-4.88113248793301e-25 wub=-2.72767992179251e-24 pub=4.97182675152879e-30
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0400913429392909 lu0=3.75966896692344e-09 wu0=1.2389005166646e-08 pu0=-2.25818237764059e-14
+  a0=2.39190022144611 la0=-2.07023940817084e-06 wa0=-1.14872436166888e-05 pa0=2.09381550446907e-11
+  keta=0.0300913079837162 lketa=-7.42786723524671e-08 wketa=-4.07608763908308e-07 pketa=7.42961129847354e-13
+  a1=0.0
+  a2=0.65972622
+  ags=0.35254400376926 lags=-3.70406287035348e-07 wags=-1.65853408479047e-06 pags=3.02306149090422e-12
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.918770161508955+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.35994254297379e-07 wnfactor=-3.14077021862959e-07 pnfactor=5.72477924137295e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.734241310869846 lpclm=-9.63625587133105e-07 wpclm=-9.51712636060203e-06 ppclm=1.73471612483865e-11
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.25627534538694e-05 lalpha0=3.47092921127515e-12 walpha0=2.85681693628491e-11 palpha0=-5.20720879109153e-17
+  alpha1=0.0
+  beta0=27.5877927304813 lbeta0=3.60938517657701e-06 wbeta0=-6.79018718650242e-06 pbeta0=1.2376684680641e-11
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.397415793544776 lkt1=4.49955611536631e-08 wkt1=2.46915897691003e-07 pkt1=-4.50061261114222e-13
+  kt2=-0.019151
+  at=9418.152 lat=0.011996938386888
+  ute=-1.2986
+  ua1=3.0044e-9
+  ub1=-4.49356752221417e-18 lub1=1.35076674583296e-24 wub1=7.41241524868391e-24 pub1=-1.35108390586489e-29
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.81e-6
+  sbref=2.81e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.21 nmos
* DC IV MOS Parameters
+  lmin=8.0e-07 lmax=1e-06 wmin=1.0e-05 wmax=1.5e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.826248519060131+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-1.95627948688349e-08 wvth0=-4.32226278908112e-07 pvth0=2.69160702890724e-13
+  k1=0.88325
+  k2=-0.0378756277071716 lk2=1.09668083489147e-08 wk2=6.98771990465537e-08 pk2=-4.35146980394595e-14
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=79042.5976422054 lvsat=0.00799399931527178 wvsat=0.521362917974553 pvsat=-3.2466885127321e-7
+  ua=-2.34207639686137e-10 lua=5.26072610236955e-17 wua=8.9442814779589e-16 pua=-5.56988134905083e-22
+  ub=-1.40460910456996e-20 lub=1.08816394248298e-24 wub=1.36383996089625e-23 pub=-8.49305422688886e-30
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0480904204700456 lu0=-2.82142008903199e-09 wu0=-6.19450258332292e-08 pu0=3.8575087882153e-14
+  a0=-4.00588837640129 la0=3.19341960272475e-06 wa0=5.74362180834438e-05 pa0=-3.5767313523321e-11
+  keta=-0.214416539918581 lketa=1.26885513860038e-07 wketa=2.03804381954154e-06 pketa=-1.26915306578692e-12
+  a1=0.0
+  a2=0.65972622
+  ags=-0.900750245101301 lags=6.60717743632178e-07 wags=8.29267042395233e-06 pags=-5.16410294577826e-12
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.663439661805224+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=7.40740630543705e-08 wnfactor=1.57038510931479e-06 pnfactor=-9.77927489508702e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-4.99792710499923 lpclm=3.75240706582327e-06 wpclm=4.758563180301e-05 ppclm=-2.96330480783202e-11
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.49804288156529e-05 lalpha0=1.48183274319966e-12 walpha0=-1.42840846814245e-10 palpha0=8.89514233774819e-17
+  alpha1=0.0
+  beta0=21.0548806775932 lbeta0=8.98421444276164e-06 wbeta0=3.39509359325125e-05 pbeta0=-2.11423002841896e-11
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.25552834227612 lkt1=-7.17396435160493e-08 wkt1=-1.23457948845501e-06 pkt1=7.68810919425079e-13
+  kt2=-0.019151
+  at=8431.72500000003 lat=0.012808502459025
+  ute=-1.4589532325 lute=1.31927575327958e-7
+  ua1=6.0953253185e-09 lua1=-2.54300007821482e-15
+  ub1=-7.22569399142912e-18 lub1=3.59857188797665e-24 wub1=-3.70620762434195e-23 pub1=2.30797038011409e-29
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.41e-6
+  sbref=2.41e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.22 nmos
* DC IV MOS Parameters
+  lmin=6e-07 lmax=8.0e-07 wmin=1.0e-05 wmax=1.5e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.788372556665+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=4.02374106944815e-9
+  k1=0.88325
+  k2=-0.00834484262750002 lk2=-7.4229269745343e-9
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=77796.1053695 lvsat=0.00877022869474586
+  ua=-2.8572090550946e-10 lua=8.46861685631195e-17
+  ub=1.0505226157e-18 lub=4.25224007162523e-25
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0362910518205 lu0=4.52641254946819e-9
+  a0=1.1222
+  keta=-0.01066
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.75091767705+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.95987911429764e-8
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=1.031604579 lpclm=-2.36922928524877e-9
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.674704005e-05 lalpha0=3.81709162623463e-13
+  alpha1=0.0
+  beta0=32.3580179100001 lbeta0=1.94540049088779e-6
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.37073
+  kt2=-0.019151
+  at=9131.64299999998 lat=0.012372641822967
+  ute=-1.13718994 lute=-6.84444015738602e-8
+  ua1=2.0117e-9
+  ub1=-1.6583655e-18 lub1=1.31623849180501e-25
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.02e-6
+  sbref=2.01e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.23 nmos
* DC IV MOS Parameters
+  lmin=5e-07 lmax=6e-07 wmin=1.0e-05 wmax=1.5e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.944065847361234+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-6.1792639399861e-08 wvth0=-1.88871524746907e-08 pvth0=7.98418485277983e-15
+  k1=0.88325
+  k2=0.000624627716505122 lk2=-1.12146001425259e-08 wk2=-6.93400638801579e-08 pk2=2.93121945441231e-14
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=76973.7384678477 lvsat=0.00911786867744824 wvsat=0.157373565850651 pvsat=-6.65266848656117e-8
+  ua=2.06868275181716e-10 lua=-1.23546548379642e-16 wua=-7.41344948929643e-16 pua=3.13389491605977e-22
+  ub=2.92689173000701e-18 lub=-3.67975384897591e-25 wub=-1.04198967344985e-23 pub=4.40481336647125e-30
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0425737092891022 lu0=1.8705384751085e-09 wu0=1.58942652363933e-08 pu0=-6.71899863764567e-15
+  a0=1.1222
+  keta=-0.01066
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.46884482213206+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-2.83891268824708e-07 wnfactor=-6.40419754680268e-07 pnfactor=2.70725283315739e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=2.18168857600595 lpclm=-4.88545387423572e-07 wpclm=-1.99138387117761e-05 ppclm=8.41819695246782e-12
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=2.792252773e-05 lalpha0=-4.34251591983062e-12
+  alpha1=0.0
+  beta0=36.96
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.435276200000001 lkt1=2.72856796721998e-8
+  kt2=-0.019151
+  at=79101.9518433424 lat=-0.017205976804688 wat=-0.768658677123809 pat=3.24935851239225e-7
+  ute=-1.300713655 lute=6.82141991804604e-10
+  ua1=-1.192050637e-09 lua1=1.35432471052965e-15
+  ub1=6.41629420500001e-18 lub1=-3.28178512257386e-24
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=1.81e-6
+  sbref=1.81e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.24 nmos
* DC IV MOS Parameters
+  lmin=2.0e-05 lmax=1.0e-04 wmin=7e-06 wmax=1.0e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.791968+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+  k1=0.88325
+  k2=-0.0388233
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=105660.0
+  ua=-6.02229e-11
+  ub=1.73106e-18
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0426101
+  a0=0.9440931
+  keta=-0.02132
+  a1=0.0
+  a2=0.65972622
+  ags=0.1460627
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.93087+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.33405
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.4467e-5
+  alpha1=0.0
+  beta0=24.0
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.40273
+  kt2=-0.019151
+  at=160000.0
+  ute=-1.2986
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.25 nmos
* DC IV MOS Parameters
+  lmin=8e-06 lmax=2.0e-05 wmin=7e-06 wmax=1.0e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.791968+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+  k1=0.88325
+  k2=-0.0388233
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=105660.0
+  ua=-6.02229e-11
+  ub=1.73106e-18
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0426101
+  a0=0.9440931
+  keta=-0.02132
+  a1=0.0
+  a2=0.65972622
+  ags=0.1460627
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.93087+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.33405
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.4467e-5
+  alpha1=0.0
+  beta0=24.0
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.40273
+  kt2=-0.019151
+  at=160000.0
+  ute=-1.2986
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.26 nmos
* DC IV MOS Parameters
+  lmin=4e-06 lmax=8e-06 wmin=7e-06 wmax=1.0e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.787009917893+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=3.87857425989748e-8
+  k1=0.88325
+  k2=-0.040038259480075 lk2=9.50430118852657e-9
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=110438.41375 lvsat=-0.037380245372951
+  ua=-1.026911477714e-10 lua=3.32217678357012e-16
+  ub=1.872940661065e-18 lub=-1.10989424561367e-24
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0426265377433 lu0=-1.2858804408272e-10
+  a0=1.03171951755192 la0=-6.85477893002312e-7
+  keta=-0.01729370857425 lketa=-3.14965947512487e-8
+  a1=0.0
+  a2=0.65972622
+  ags=0.158828805742775 lags=-9.98658111432839e-8
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.970406595367501+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-3.09284150215798e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.2603764168025 lpclm=5.76328623160164e-7
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.4467e-5
+  alpha1=0.0
+  beta0=21.51522485 lbeta0=1.94377275939346e-5
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.414198193 lkt1=8.97125888950823e-8
+  kt2=-0.019151
+  at=236454.62 lat=-0.59808392596722
+  ute=-1.33682731 lute=2.99041962983603e-7
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.27 nmos
* DC IV MOS Parameters
+  lmin=2e-06 lmax=4e-06 wmin=7e-06 wmax=1.0e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.803592063161+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-2.46033381635127e-8
+  k1=0.88325
+  k2=-0.04195453332085 lk2=1.68297006041463e-08 wk2=2.11758236813575e-22
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=93870.327025 lvsat=0.0259550933613946
+  ua=1.037893167889e-10 lua=-4.57101594412048e-16 wua=-9.86076131526265e-32 pua=3.76158192263132e-37
+  ub=1.535692017715e-18 lub=1.79316598028319e-25
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.04299289831795 lu0=-1.52908596997528e-09 wu0=-2.11758236813575e-22
+  a0=0.484478507841295 la0=1.40647727928978e-6
+  keta=-0.0390877390815 lketa=5.18161212837616e-8
+  a1=0.0
+  a2=0.65972622
+  ags=0.1175536953818 lags=5.79178327620362e-8
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.93082131177+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.57960259463844e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.598489405835 lpclm=-7.16186381517035e-7
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.4467e-5
+  alpha1=0.0
+  beta0=23.895067196 lbeta0=1.03402304827678e-5
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.407134579 lkt1=6.27102926852487e-8
+  kt2=-0.019151
+  at=138327.392 lat=-0.222969929547552
+  ute=-1.22214538 lute=-1.39356205967219e-7
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.28 nmos
* DC IV MOS Parameters
+  lmin=1e-06 lmax=2e-06 wmin=7e-06 wmax=1.0e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.788553847568+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=2.80728358253129e-9
+  k1=0.88325
+  k2=-0.0408446990747 lk2=1.4806771318827e-8
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=113605.84308 lvsat=-0.0100174435530516
+  ua=-1.457233283565e-10 lua=-2.30716121352835e-18
+  ub=1.62915829593e-18 lub=8.95271527121714e-27
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0413299526304 lu0=1.50201668603836e-09 wu0=2.11758236813575e-22
+  a0=1.24344551694185 la0=2.30845838249147e-8
+  keta=-0.01066
+  a1=0.0
+  a2=0.65972622
+  ags=0.186729528529 lags=-6.81711027661927e-8
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.88736983212+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-7.87599005099196e-8
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-0.21724791552 lpclm=7.70683321973685e-07 ppclm=8.07793566946316e-28
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.5418899767e-05 lalpha0=-1.73505721420369e-12
+  alpha1=0.0
+  beta0=26.908933408 lbeta0=4.84676310830273e-6
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.37273
+  kt2=-0.019151
+  at=9418.15199999999 lat=0.011996938386888
+  ute=-1.2986
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.81e-6
+  sbref=2.81e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.29 nmos
* DC IV MOS Parameters
+  lmin=8.0e-07 lmax=1e-06 wmin=7e-06 wmax=1.0e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.783036037460001+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=7.34695701049632e-9
+  k1=0.88325
+  k2=-0.030889548134 lk2=6.61636003023396e-9
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=131166.650712 lvsat=-0.0244652643769344
+  ua=-1.4478582114954e-10 lua=-3.07847745541804e-18
+  ub=1.3494737154e-18 lub=2.39057889895242e-25
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0418973720144999 lu0=1.03518316873834e-9
+  a0=1.73638514612 la0=-3.82472130228453e-7
+  keta=-0.01066
+  a1=0.0
+  a2=0.65972622
+  ags=-0.0716778688999997 lags=1.44428673727966e-7
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.82044130875+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-2.36957295491962e-8
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-0.240480973049999 lpclm=7.897978786284e-7
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=6.99697250000007e-07 lalpha0=1.03748869918102e-11
+  alpha1=0.0
+  beta0=24.44917729 lbeta0=6.87048071902103e-6
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.37895731 lkt1=5.12340098360974e-9
+  kt2=-0.019151
+  at=8431.72500000003 lat=0.012808502459025
+  ute=-1.4589532325 lute=1.31927575327956e-7
+  ua1=6.0953253185e-09 lua1=-2.54300007821482e-15
+  ub1=-1.09310316025e-17 lub1=5.90600048385643e-24
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.41e-6
+  sbref=2.41e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.30 nmos
* DC IV MOS Parameters
+  lmin=6e-07 lmax=8.0e-07 wmin=7e-06 wmax=1.0e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.788372556664999+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=4.02374106944815e-9
+  k1=0.88325
+  k2=-0.00834484262749999 lk2=-7.4229269745343e-9
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=77796.1053695001 lvsat=0.00877022869474592
+  ua=-2.8572090550946e-10 lua=8.46861685631195e-17
+  ub=1.0505226157e-18 lub=4.25224007162523e-25
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0362910518205 lu0=4.52641254946824e-9
+  a0=1.1222
+  keta=-0.01066
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.750917677049999+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.95987911429764e-8
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=1.031604579 lpclm=-2.36922928524877e-9
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.674704005e-05 lalpha0=3.81709162623463e-13
+  alpha1=0.0
+  beta0=32.35801791 lbeta0=1.94540049088779e-6
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.37073
+  kt2=-0.019151
+  at=9131.64300000004 lat=0.012372641822967
+  ute=-1.13718994 lute=-6.84444015738602e-8
+  ua1=2.0117e-9
+  ub1=-1.6583655e-18 lub1=1.316238491805e-25
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.02e-6
+  sbref=2.01e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.31 nmos
* DC IV MOS Parameters
+  lmin=5e-07 lmax=6e-07 wmin=7e-06 wmax=1.0e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.904633522594727+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-4.51233733189911e-08 wvth0=3.75528682288915e-07 pvth0=-1.58747615392671e-13
+  k1=0.88325
+  k2=-0.0223912797040854 lk2=-1.4850625827123e-09 wk2=1.60873051676371e-07 pk2=-6.80060260082039e-14
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=97233.929958093 lvsat=0.000553257668585383 wvsat=-0.0452759199814192 pvsat=1.91395349296657e-8
+  ua=1.38356425709113e-10 lua=-9.4584465740239e-17 wua=-5.60655883810525e-17 pua=2.37006622419106e-23
+  ub=4.80385025599818e-18 lub=-1.16142393954837e-24 wub=-2.91938890930292e-23 pub=1.23411619301853e-29
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0447917611813147 lu0=9.32899180661649e-10 wu0=-6.29146167157398e-09 pu0=2.65959588388594e-15
+  a0=1.1222
+  keta=-0.01066
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.9224723284691+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-4.75653678206073e-07 wnfactor=-5.17775993543558e-06 pnfactor=2.18879963526662e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.190772171999999 lpclm=3.53076694958269e-7
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=2.792252773e-05 lalpha0=-4.34251591983062e-12
+  alpha1=0.0
+  beta0=36.96
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.4352762 lkt1=2.72856796722e-8
+  kt2=-0.019151
+  at=-70061.8647164159 lat=0.0458501925334352 wat=0.723329725115057 pat=-3.05773898027614e-7
+  ute=-1.300713655 lute=6.82141991805451e-10
+  ua1=-1.19205063700001e-09 lua1=1.35432471052965e-15
+  ub1=7.922877386592e-18 lub1=-3.91866453751142e-24 wub1=-1.50693692732303e-23 pub1=6.37028954224194e-30
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=1.81e-6
+  sbref=1.81e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.32 nmos
* DC IV MOS Parameters
+  lmin=2.0e-05 lmax=1.0e-04 wmin=5.0e-06 wmax=7.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.776028018098001+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} wvth0=1.11617300391504e-7
+  k1=0.88325
+  k2=-0.0376359927022 wk2=-8.31393888213531e-9
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=119341.42178 wvsat=-0.0958020764383392
+  ua=-3.818978876704e-10 wua=2.25248020656385e-15
+  ub=2.18684893802e-18 wub=-3.19159275856647e-24
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0419270293806 wu0=4.78309818561439e-9
+  a0=1.2307971730372 wa0=-2.00760169242389e-6
+  keta=-0.016990467806 wketa=-3.03168910995915e-8
+  a1=0.0
+  a2=0.65972622
+  ags=0.17196595846056 wags=-1.81383630074785e-7
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.86478898292+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} wnfactor=4.62722277788102e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.6563262699 wpclm=-2.25669059398173e-6
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=2.3873915414e-05 walpha0=-6.58704953353921e-11
+  alpha1=0.0
+  beta0=26.71377379 wbeta0=-1.9002788470859e-5
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.40273
+  kt2=-0.019151
+  at=180009.392 wat=-0.140112726052416
+  ute=-1.2986
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.33 nmos
* DC IV MOS Parameters
+  lmin=8e-06 lmax=2.0e-05 wmin=5.0e-06 wmax=7.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.776028018098+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} wvth0=1.11617300391508e-7
+  k1=0.88325
+  k2=-0.0376359927021999 wk2=-8.3139388821352e-9
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=119341.42178 wvsat=-0.0958020764383396
+  ua=-3.818978876704e-10 wua=2.25248020656385e-15
+  ub=2.18684893802e-18 wub=-3.19159275856647e-24
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0419270293805999 wu0=4.78309818561439e-9
+  a0=1.2307971730372 wa0=-2.00760169242389e-6
+  keta=-0.016990467806 wketa=-3.03168910995915e-8
+  a1=0.0
+  a2=0.65972622
+  ags=0.17196595846056 wags=-1.81383630074786e-7
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.864788982919999+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} wnfactor=4.62722277788106e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.6563262699 wpclm=-2.25669059398172e-6
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=2.3873915414e-05 walpha0=-6.5870495335392e-11
+  alpha1=0.0
+  beta0=26.71377379 wbeta0=-1.9002788470859e-5
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.40273
+  kt2=-0.019151
+  at=180009.392 wat=-0.140112726052416
+  ute=-1.2986
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.34 nmos
* DC IV MOS Parameters
+  lmin=4e-06 lmax=8e-06 wmin=5.0e-06 wmax=7.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.76609805199018+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=7.76794537006013e-08 wvth0=1.46432162380885e-07 pvth0=-2.72347300145025e-13
+  k1=0.88325
+  k2=-0.0355441712559598 lk2=-1.63637564739681e-08 wk2=-3.14691696879567e-08 pk2=1.81137141836854e-13
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=142358.044629165 lvsat=-0.180052849077472 wvsat=-0.22351236344746 pvsat=9.99043221205142e-7
+  ua=-5.30719753909936e-10 lua=1.16419342650987e-15 wua=2.99720525413697e-15 pua=-5.8257837161267e-21
+  ub=2.47088245558924e-18 lub=-2.22191780292793e-24 wub=-4.18699652900322e-24 pub=7.78677593251241e-30
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0414852410840166 lu0=3.4559910031198e-09 wu0=7.9917563795395e-09 pu0=-2.51004699220233e-14
+  a0=1.5374306826202 la0=-2.39871146105371e-06 wa0=-3.54116556529356e-06 pa0=1.19966576487776e-11
+  keta=-0.00289372094974119 lketa=-1.10275058631608e-07 wketa=-1.00833724542504e-07 pketa=5.51634218995709e-13
+  a1=0.0
+  a2=0.65972622
+  ags=0.216743443729466 lags=-3.50282222115116e-07 wags=-4.05538449476832e-07 pags=1.7535028545358e-12
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.893712518208824+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-2.26261036133485e-07 wnfactor=5.37038617803899e-07 pnfactor=-5.81356736848089e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.398382235922076 lpclm=2.01782679086416e-06 wpclm=-9.66364771500327e-07 ppclm=-1.00938718116257e-11
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=3.56295526813255e-05 lalpha0=-9.19611880758626e-11 walpha0=-1.48187558442974e-10 palpha0=6.4394424140064e-16
+  alpha1=0.0
+  beta0=26.8487990558172 lbeta0=-1.05626633269107e-06 wbeta0=-3.73475426729554e-05 pbeta0=1.4350607738412e-10
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.414198193 lkt1=8.97125888950823e-8
+  kt2=-0.019151
+  at=275586.642772388 lat=-0.747675122511933 wat=-0.274016041396186 pat=1.04748961594248e-6
+  ute=-1.33682731 lute=2.9904196298361e-7
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.35 nmos
* DC IV MOS Parameters
+  lmin=2e-06 lmax=4e-06 wmin=5.0e-06 wmax=7.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.792617456874918+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-2.36970974538422e-08 wvth0=7.68480123781366e-08 pvth0=-6.34581282087204e-15
+  k1=0.88325
+  k2=-0.0464348021430451 lk2=2.52681958276506e-08 wk2=3.13724014265605e-08 pk2=-5.90892801513148e-14
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=73149.6607673882 lvsat=0.0845121853708424 wvsat=0.145093315927656 pvsat=-4.10037136118172e-7
+  ua=1.17870375291842e-10 lua=-1.31519216668377e-15 wua=-9.86004718459581e-17 pua=6.00864880256573e-21
+  ub=1.73364004840338e-18 lub=5.96361601536086e-25 wub=-1.3861009967947e-24 pub=-2.92029424622259e-30
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0442274290163249 lu0=-7.02665581354086e-09 wu0=-8.64461356670417e-09 pu0=3.84958971989523e-14
+  a0=0.282402129461553 la0=2.39892509499099e-06 wa0=1.41500912399463e-06 pa0=-6.94946497737973e-12
+  keta=-0.0509533314757667 lketa=7.34439043741559e-08 wketa=8.3087007170809e-08 pketa=-1.51445263667456e-13
+  a1=0.0
+  a2=0.65972622
+  ags=0.125423325374416 lags=-1.18997475559567e-09 wags=-5.5105887839532e-08 pags=4.13893437755475e-13
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.86337673144876+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.10295483676393e-07 wnfactor=4.72270422123277e-07 pnfactor=-3.33765347405714e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=1.58217464218495 lpclm=-2.50749313812152e-06 wpclm=-6.8881063473846e-06 ppclm=1.25433532844959e-11
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=8.93577904908678e-06 lalpha0=1.0081927895079e-11 walpha0=3.87315339631854e-11 palpha0=-7.05971676322509e-17
+  alpha1=0.0
+  beta0=23.8424799613759 lbeta0=1.04360828655213e-05 wbeta0=3.68234117195296e-07 pbeta0=-6.71191740669546e-13
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.407134579 lkt1=6.27102926852487e-8
+  kt2=-0.019151
+  at=147445.326772388 lat=-0.257825341457937 wat=-0.0638469523175615 pat=2.44069723879864e-7
+  ute=-1.22214538 lute=-1.39356205967222e-7
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.36 nmos
* DC IV MOS Parameters
+  lmin=1e-06 lmax=2e-06 wmin=5.0e-06 wmax=7.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.772059441820768+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=1.37746338838208e-08 wvth0=1.15499569095311e-07 pvth0=-7.67972034475343e-14
+  k1=0.88325
+  k2=-0.0391684962943441 lk2=1.20236749017418e-08 wk2=-1.17373551866199e-08 pk2=1.94882096299835e-14
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=125704.672891147 lvsat=-0.0112814644325093 wvsat=-0.0847202167304282 pvsat=8.85111407722944e-9
+  ua=-9.7971348799031e-10 lua=6.85407966020373e-16 wua=5.83988932633149e-15 pua=-4.81562064575605e-21
+  ub=2.37254127214367e-18 lub=-5.68183464913286e-25 wub=-5.20542629672385e-24 pub=4.04130837704257e-30
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0369952004021475 lu0=6.15575148060733e-09 wu0=3.03534435959992e-08 pu0=-3.258707053128e-14
+  a0=1.59039003104256 la0=1.48149991543372e-08 wa0=-2.42942622442409e-06 pa0=5.79065096788477e-14
+  keta=-0.01066
+  a1=0.0
+  a2=0.65972622
+  ags=0.150777410837121 lags=-4.7403652305118e-08 wags=2.51749239415493e-07 pags=-1.45420915201204e-13
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.83239112336181+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-5.38170552624582e-08 wnfactor=3.84980051315495e-07 pnfactor=-1.74658482532875e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.154574198787607 lpclm=9.46384456725589e-08 wpclm=-2.60362783847764e-06 ppclm=4.73390148747744e-12
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=4.75698636328951e-05 lalpha0=-6.03376157324504e-11 walpha0=-2.25132237524422e-10 palpha0=4.10355508435128e-16
+  alpha1=0.0
+  beta0=32.6707548893432 lbeta0=-5.65548752220742e-06 wbeta0=-4.03462791262406e-05 pbeta0=7.35404136980518e-11
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.37273
+  kt2=-0.019151
+  at=3529.04277238801 lat=0.00449533079366646 wat=0.0412375922217505 pat=5.25288669271798e-8
+  ute=-1.2986
+  ua1=3.0044e-9
+  ub1=-3.1351619841418e-18 lub1=-1.12524113898323e-24 wub1=-4.32281562066863e-24 pub1=7.87933003907695e-30
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.81e-6
+  sbref=2.81e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.37 nmos
* DC IV MOS Parameters
+  lmin=8.0e-07 lmax=1e-06 wmin=5.0e-06 wmax=7.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.774397233919526+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=1.18512598526184e-08 wvth0=6.04919086940245e-08 pvth0=-3.15406959979254e-14
+  k1=0.88325
+  k2=-0.0324574764400287 lk2=6.50231082598111e-09 wk2=1.09791796378636e-08 pk2=7.98612217301295e-16
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=197926.601083172 lvsat=-0.0707006836358625 wvsat=-0.467476404961681 pvsat=3.23756495576915e-7
+  ua=-1.3828407270095e-10 lua=-6.86209825005792e-18 wua=-4.55275052454843e-17 pua=2.64942295041049e-23
+  ub=1.174081169333e-18 lub=4.17826813932237e-25 wub=1.22815964416713e-24 pub=-1.25180221769259e-30
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0443842146673082 lu0=7.65803852172632e-11 wu0=-1.74137376762074e-08 pu0=6.71247028398351e-15
+  a0=3.12224725792007 la0=-1.24549142897182e-06 wa0=-9.70428878683901e-06 pa0=6.04316146051705e-12
+  keta=-0.01066
+  a1=0.0
+  a2=0.65972622
+  ags=-0.115735225298413 lags=1.71864555335306e-07 wags=3.08504941461718e-07 pags=-1.92115590701397e-13
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.819376745690837+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-4.31097233068422e-08 wnfactor=7.45444100818884e-09 pnfactor=1.35943540360869e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-3.65175328036066 lpclm=3.22622205891969e-06 wpclm=2.38869158185522e-05 ppclm=-1.70606899860143e-11
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=-0.000137517249337248 lalpha0=9.19392898085885e-11 walpha0=9.67843159501324e-10 palpha0=-5.71142332935261e-16
+  alpha1=0.0
+  beta0=-4.3599301167161 lbeta0=2.48108049835127e-05 wbeta0=0.000201731395631203 pbeta0=-1.25624393732815e-10
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.378957310000001 lkt1=5.12340098360974e-9
+  kt2=-0.019151
+  at=-53302.0765858201 lat=0.0512520544543643 wat=0.432281562066864 pat=-2.6919512942746e-7
+  ute=-1.4589532325 lute=1.31927575327956e-7
+  ua1=6.0953253185e-09 lua1=-2.54300007821482e-15
+  ub1=-1.25380410249067e-17 lub1=6.61079893710431e-24 wub1=1.12528392149707e-23 pub1=-4.93524403950343e-30
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.41e-6
+  sbref=2.41e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.38 nmos
* DC IV MOS Parameters
+  lmin=6e-07 lmax=8.0e-07 wmin=5.0e-06 wmax=7.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.783995817037795+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=5.87392458879556e-09 wvth0=3.06474539750749e-08 pvth0=-1.29556288663402e-14
+  k1=0.88325
+  k2=-0.0137970764584721 lk2=-5.11809871493364e-09 wk2=3.81784386618396e-08 pk2=-1.61392095539581e-14
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=54486.4623478138 lvsat=0.0186239373989464 wvsat=0.163222232193618 pvsat=-6.89990974374405e-8
+  ua=-2.84394807916967e-10 lua=8.41255860017476e-17 wua=-9.28579682459402e-18 pua=3.92539417745779e-24
+  ub=1.39825535786074e-18 lub=2.78226597336171e-25 wub=-2.43494567160378e-24 pub=1.02932701870274e-30
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0392412079630242 lu0=3.27929009318284e-09 wu0=-2.06580199642923e-08 pu0=8.732785437525e-15
+  a0=1.1222
+  keta=-0.01066
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.650533026169797+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=6.20344949942155e-08 wnfactor=7.02928259321684e-07 pnfactor=-2.97149565991316e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=2.59220040443708 lpclm=-6.6208146316809e-07 wpclm=-1.09278350570577e-05 ppclm=4.61953464150504e-12
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=-5.79083269222719e-06 lalpha0=9.90916664481787e-12 walpha0=1.57818028120789e-10 palpha0=-6.67145728455292e-17
+  alpha1=0.0
+  beta0=32.35801791 lbeta0=1.94540049088779e-6
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.37073
+  kt2=-0.019151
+  at=9131.64299999992 lat=0.012372641822967
+  ute=-1.13718994 lute=-6.84444015738594e-8
+  ua1=2.0117e-9
+  ub1=-3.1380461568843e-18 lub1=7.57130732945857e-25 wub1=1.03612388883725e-23 pub1=-4.38001687652058e-30
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.02e-6
+  sbref=2.01e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.39 nmos
* DC IV MOS Parameters
+  lmin=5e-07 lmax=6e-07 wmin=5.0e-06 wmax=7.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={1.02512339348845+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-9.6058176931766e-08 wvth0=-4.68183324184009e-07 pvth0=1.97915604815631e-13
+  k1=0.88325
+  k2=-8.95242876995939e-05 lk2=-1.09127059516365e-08 wk2=4.70839923995237e-09 pk2=-1.99038631910435e-15
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=98381.6808445817 lvsat=6.80677885890879e-05 wvsat=-0.0533128711059225 pvsat=2.25370033154777e-8
+  ua=1.40656959956311e-10 lua=-9.55569728830913e-17 wua=-7.21747297658531e-17 pua=3.05104956886496e-23
+  ub=2.64023953159718e-19 lub=7.57701373276843e-25 wub=2.59555453899915e-24 pub=-1.09722136582564e-30
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0371862044551142 lu0=4.14800378108516e-09 wu0=4.69652932590234e-08 pu0=-1.98536853846803e-14
+  a0=1.1222
+  keta=-0.01066
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={2.14482677345016+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-5.69649795087357e-07 wnfactor=-6.73476313853976e-06 pnfactor=2.84699315631805e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.190772172000003 lpclm=3.53076694958267e-7
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=2.792252773e-05 lalpha0=-4.34251591983064e-12
+  alpha1=0.0
+  beta0=36.96
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.435276200000001 lkt1=2.72856796722002e-8
+  kt2=-0.019151
+  at=110728.117074624 lat=-0.0305753372590729 wat=-0.542624642299468 pat=2.29384257663896e-7
+  ute=-1.300713655 lute=6.82141991804604e-10
+  ua1=-1.192050637e-09 lua1=1.35432471052965e-15
+  ub1=5.770832205e-18 lub1=-3.00892832585186e-24
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=1.81e-6
+  sbref=1.81e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.40 nmos
* DC IV MOS Parameters
+  lmin=2.0e-05 lmax=1.0e-04 wmin=3.0e-06 wmax=5.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.798699780586+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} wvth0=-1.79474534681639e-9
+  k1=0.88325
+  k2=-0.041738908924 wk2=1.22102758741536e-8
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=133465.022884 wvsat=-0.166453244173732
+  ua=3.947692489668e-10 wua=-1.63267909105897e-15
+  ub=1.249189664904e-18 wub=1.4989052309868e-24
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.04614916916614 wu0=-1.63375143263021e-8
+  a0=0.62735805610454 wa0=1.01101076728597e-6
+  keta=-0.012123954454 wketa=-5.4660884432942e-8
+  a1=0.0
+  a2=0.65972622
+  ags=0.10429923799464 wags=1.57108853714468e-7
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.9406269686+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} wnfactor=8.33542817977267e-8
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-0.83685494384 wpclm=5.21272146420814e-6
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=5.060084586e-06 walpha0=2.82428336793921e-11
+  alpha1=0.0
+  beta0=21.58646101 wbeta0=6.64581435954855e-6
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.40273
+  kt2=-0.019151
+  at=209645.0816 wat=-0.288360758651597
+  ute=-1.2986
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.41 nmos
* DC IV MOS Parameters
+  lmin=8e-06 lmax=2.0e-05 wmin=3.0e-06 wmax=5.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.798699780586+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} wvth0=-1.79474534681555e-9
+  k1=0.88325
+  k2=-0.041738908924 wk2=1.22102758741535e-8
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=133465.022884 wvsat=-0.166453244173732
+  ua=3.947692489668e-10 wua=-1.63267909105897e-15
+  ub=1.249189664904e-18 wub=1.49890523098681e-24
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.04614916916614 wu0=-1.63375143263021e-8
+  a0=0.62735805610454 wa0=1.01101076728597e-6
+  keta=-0.012123954454 wketa=-5.4660884432942e-8
+  a1=0.0
+  a2=0.65972622
+  ags=0.10429923799464 wags=1.57108853714469e-7
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.9406269686+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} wnfactor=8.33542817977267e-8
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-0.83685494384 wpclm=5.21272146420814e-6
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=5.060084586e-06 walpha0=2.82428336793921e-11
+  alpha1=0.0
+  beta0=21.58646101 wbeta0=6.64581435954855e-6
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.40273
+  kt2=-0.019151
+  at=209645.0816 wat=-0.288360758651597
+  ute=-1.2986
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.42 nmos
* DC IV MOS Parameters
+  lmin=4e-06 lmax=8e-06 wmin=3.0e-06 wmax=5.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.793977815715114+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=3.69386609763872e-08 wvth0=6.96788207098502e-09 pvth0=-6.85476771426777e-14
+  k1=0.88325
+  k2=-0.0450760620484701 lk2=2.61056511985391e-08 wk2=1.62126651541757e-08 pk2=-3.13096146948975e-14
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=138701.535465055 lvsat=-0.0409638292997088 wvsat=-0.205221232143392 pvsat=3.0327154129789e-7
+  ua=3.94811634571485e-10 lua=-3.31571183723714e-19 wua=-1.63262483597029e-15 pua=-4.24422964128786e-25
+  ub=1.3214761304438e-18 lub=-5.6547757485861e-25 wub=1.56273390277543e-24 pub=-4.993145294897e-31
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0461768115720998 lu0=-2.16239106016391e-10 wu0=-1.54771118683824e-08 pu0=-6.73069698004468e-15
+  a0=0.627864755942601 la0=-3.96377653089588e-09 wa0=1.00879972889027e-06 pa0=1.7296358600231e-14
+  keta=-0.012123954454 wketa=-5.46608844329421e-8
+  a1=0.0
+  a2=0.65972622
+  ags=0.100686011543886 lags=2.82652985663355e-08 wags=1.75021214301842e-07 pags=-1.4012357845003e-13
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.990044954536936+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-3.86583610546431e-07 wnfactor=5.51502476028439e-08 pnfactor=2.20632572621372e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-0.83685494384 wpclm=5.21272146420814e-6
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=-7.52621277122709e-06 lalpha0=9.84592185115985e-11 walpha0=6.76925985570713e-11 palpha0=-3.08604898651333e-16
+  alpha1=0.0
+  beta0=16.9122792731474 lbeta0=3.65648663725107e-05 wbeta0=1.23583871888432e-05 pbeta0=-4.46879205614811e-11
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.414198193 lkt1=8.97125888950823e-8
+  kt2=-0.019151
+  at=304851.727776492 lat=-0.744775982450879 wat=-0.420410180836297 pat=1.03298710845634e-6
+  ute=-1.33682731 lute=2.99041962983613e-7
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.43 nmos
* DC IV MOS Parameters
+  lmin=2e-06 lmax=4e-06 wmin=3.0e-06 wmax=5.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.808197364660361+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-1.74188495826241e-08 wvth0=-1.0881081725596e-09 pvth0=-3.7751793502973e-14
+  k1=0.88325
+  k2=-0.0407002493996922 lk2=9.37809653586388e-09 wk2=2.68617297995467e-09 pk2=2.03985262607549e-14
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=145535.509743893 lvsat=-0.0670882746286273 wvsat=-0.217005890928268 pvsat=3.48321121759255e-7
+  ua=4.6968531468265e-10 lua=-2.86553509228757e-16 wua=-1.85850123027769e-15 pua=8.6304027172297e-22
+  ub=1.14244723413934e-18 lub=1.18901736940237e-25 wub=1.57125119525339e-24 pub=-5.31873847481273e-31
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0464302606404529 lu0=-1.18510671653069e-09 wu0=-1.96639439359974e-08 pu0=9.27443575662109e-15
+  a0=0.187022990318489 la0=1.68125570701513e-06 wa0=1.89212876992866e-06 pa0=-3.35943294977749e-12
+  keta=-0.0403690368951649 lketa=1.07973352245397e-07 wketa=3.01406823441246e-08 pketa=-3.24173578167263e-13
+  a1=0.0
+  a2=0.65972622
+  ags=0.0198783102854944 lags=3.37171403205526e-07 wags=4.72867007300503e-07 pags=-1.27870792456559e-12
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.906206048959413+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-6.60900271891615e-08 wnfactor=2.58023271332498e-07 pnfactor=-5.54896424253705e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-0.836854943840001 wpclm=5.21272146420814e-6
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=2.16595411307164e-05 lalpha0=-1.31100676877318e-11 walpha0=-2.49171518383305e-11 palpha0=4.54172650874319e-17
+  alpha1=0.0
+  beta0=24.1149404514226 lbeta0=9.03103020382165e-06 wbeta0=-9.94708070268526e-07 pbeta0=6.35737063147799e-12
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.407134579 lkt1=6.27102926852487e-8
+  kt2=-0.019151
+  at=178386.59193097 lat=-0.261333787234989 wat=-0.218625928201064 pat=2.61620190595806e-7
+  ute=-1.22214538 lute=-1.3935620596722e-7
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.44 nmos
* DC IV MOS Parameters
+  lmin=1e-06 lmax=2e-06 wmin=3.0e-06 wmax=5.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.804975277380067+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-1.15458512121256e-08 wvth0=-4.91568950830722e-08 pvth0=4.98646745312077e-14
+  k1=0.88325
+  k2=-0.0461855968289395 lk2=1.93764093409232e-08 wk2=2.33646236384126e-08 pk2=-1.72927267863867e-14
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=123016.696134823 lvsat=-0.026042534980152 wvsat=-0.0712740215793801 pvsat=8.26911258090888e-8
+  ua=6.93929683953229e-10 lua=-6.95290672673689e-16 wua=-2.53225624755393e-15 pua=2.09111442811791e-21
+  ub=8.38919166452132e-19 lub=6.72151755283805e-25 wub=2.46628517643801e-24 pub=-2.1632800310399e-30
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0473175156701152 lu0=-2.80233396400218e-09 wu0=-2.12823695400881e-08 pu0=1.22243902763913e-14
+  a0=1.09398826116445 la0=2.81019919207959e-08 wa0=5.37481763221227e-08 pa0=-8.55965201245845e-15
+  keta=0.043161769716436 lketa=-4.42808384205731e-08 wketa=-2.69235222097474e-07 pketa=2.21508163511477e-13
+  a1=0.0
+  a2=0.65972622
+  ags=0.268348640459815 lags=-1.15723170183443e-07 wags=-3.36382965945132e-07 pags=1.96337088418399e-13
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.994522832221622+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-2.2706776586147e-07 wnfactor=-4.26059178235965e-07 pnfactor=6.92001863130672e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-2.26529280080043 lpclm=2.60365796345534e-06 wpclm=9.50138900717756e-06 ppclm=-7.81708727926421e-12
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=-9.94292616198666e-06 lalpha0=4.44927291231641e-11 walpha0=6.25667514804244e-11 palpha0=-1.14042357492665e-16
+  alpha1=0.0
+  beta0=21.7244614970318 lbeta0=1.33882302988374e-05 wbeta0=1.44108897322017e-05 pbeta0=-2.17228900566161e-11
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.37273
+  kt2=-0.019151
+  at=31724.679544776 lat=0.00599142699061089 wat=-0.0998067949953312 pat=4.50448731085871e-8
+  ute=-1.2986
+  ua1=3.0044e-9
+  ub1=-3.9993193e-18 lub1=4.49885189508299e-25 wub1=-5.87747175411144e-39
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.81e-6
+  sbref=2.81e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.45 nmos
* DC IV MOS Parameters
+  lmin=8.0e-07 lmax=1e-06 wmin=3.0e-06 wmax=5.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.777072586230272+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=1.14105577802381e-08 wvth0=4.71088654130779e-08 pvth0=-2.93361508675494e-14
+  k1=0.88325
+  k2=-0.032191838640235 lk2=7.8633106725722e-09 wk2=9.65036692134118e-09 pk2=-6.00958264329371e-15
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=80434.7155192338 lvsat=0.00899098051369196 wvsat=0.120258893805318 pvsat=-7.48889411982797e-8
+  ua=-1.55130376037617e-10 lua=3.25735954264059e-18 wua=3.87435665580859e-17 pua=-2.41268199462835e-23
+  ub=1.55372557869567e-18 lub=8.40583609322689e-26 wub=-6.70953807719372e-25 pub=4.17823735634889e-31
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0461858959602269 lu0=-1.87131534846603e-09 wu0=-2.64263744884755e-08 pu0=1.64565226115829e-14
+  a0=1.14665659908444 la0=-1.52298824044541e-08 wa0=1.78303194206081e-07 pa0=-1.11034926431151e-13
+  keta=-0.01066
+  a1=0.0
+  a2=0.65972622
+  ags=0.0263146619035055 lags=8.34056870281681e-08 wags=-4.02078027683027e-07 pags=2.50386452257079e-13
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.479557443675287+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.96610223222644e-07 wnfactor=1.70734884680708e-06 pnfactor=-1.06321905472102e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=1.12338747725 lpclm=-1.8431435038537e-7
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=0.000118497909324933 lalpha0=-6.11795278978249e-11 walpha0=-3.12833757402122e-10 palpha0=1.94811278580781e-16
+  alpha1=0.0
+  beta0=45.8293844437591 lbeta0=-6.44363706204655e-06 wbeta0=-4.93330216817607e-05 pbeta0=3.07212019249043e-11
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.37895731 lkt1=5.12340098360974e-9
+  kt2=-0.019151
+  at=70165.52658582 lat=-0.0256350495363142 wat=-0.185346355723583 pat=1.15420921446103e-7
+  ute=-1.4589532325 lute=1.31927575327958e-7
+  ua1=6.0953253185e-09 lua1=-2.54300007821482e-15
+  ub1=-1.02885295525e-17 lub1=5.62421342975788e-24
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.41e-6
+  sbref=2.41e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.46 nmos
* DC IV MOS Parameters
+  lmin=6e-07 lmax=8.0e-07 wmin=3.0e-06 wmax=5.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.784125528945466+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=7.01847171026114e-09 wvth0=2.99985898731643e-08 pvth0=-1.86810518703037e-14
+  k1=0.88325
+  k2=-0.00247798867421287 lk2=-1.06404248306188e-08 wk2=-1.84435774775739e-08 pk2=1.14853874461871e-14
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=83481.59055986 lvsat=0.00709359697276779 wvsat=0.0181785105723455 pvsat=-1.13203220672271e-8
+  ua=-4.8919599447988e-10 lua=2.11290376180809e-16 wua=1.01520100917602e-15 pua=-6.32197139645191e-22
+  ub=1.46939705427746e-18 lub=1.36572347271746e-25 wub=-2.79082119439054e-24 pub=1.73793087320401e-30
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0307972642037701 lu0=7.71166269386406e-09 wu0=2.15815252119252e-08 pu0=-1.34394847767474e-14
+  a0=1.1222
+  keta=-0.01066
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.910070567050685+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-7.14836446100404e-08 wnfactor=-5.95368839228742e-07 pnfactor=3.70754632621752e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=1.22882231888504 lpclm=-2.49971894751598e-07 wpclm=-4.10774341755258e-06 ppclm=2.55801916615594e-12
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=2.75919307721007e-05 lalpha0=-4.56955696764102e-12 walpha0=-9.17417192946443e-12 palpha0=5.71304125980731e-18
+  alpha1=0.0
+  beta0=32.35801791 lbeta0=1.94540049088779e-6
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.37073
+  kt2=-0.019151
+  at=9131.64299999998 lat=0.012372641822967
+  ute=-1.13718994 lute=-6.84444015738602e-8
+  ua1=2.0117e-9
+  ub1=-1.59348306254102e-18 lub1=2.09538434019232e-25 wub1=2.63479678251055e-24 pub1=-1.64076963516958e-30
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.02e-6
+  sbref=2.01e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.47 nmos
* DC IV MOS Parameters
+  lmin=5e-07 lmax=6e-07 wmin=3.0e-06 wmax=5.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.932502668413154+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-5.57051448340536e-08 wvth0=-4.86222534505521e-09 pvth0=-3.94430459229243e-15
+  k1=0.88325
+  k2=0.0187817979052611 lk2=-1.96275956711463e-08 wk2=-8.96925215893597e-08 pk2=4.16045248395064e-14
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=97586.4682913488 lvsat=0.00113102790445785 wvsat=-0.0493349411806827 pvsat=1.7219706905782e-8
+  ua=5.43056588087452e-10 lua=-2.25074790300462e-16 wua=-2.08511770474841e-15 pua=6.78403690610796e-22
+  ub=-3.72204248885243e-19 lub=9.15074307759015e-25 wub=5.77818941304231e-24 pub=-1.88445554988668e-30
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0512118196040274 lu0=-9.18202725042151e-10 wu0=-2.3195714629913e-08 pu0=5.48924259883255e-15
+  a0=1.1222
+  keta=-0.01066
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.15448589471109+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.74805580487252e-07 wnfactor=-1.78073342446117e-06 pnfactor=8.71844989101646e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-1.45155395867007 lpclm=8.83106249435551e-07 wpclm=8.21548683510517e-06 ppclm=-2.65139228178033e-12
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=2.42545814257987e-05 lalpha0=-3.15875594112944e-12 walpha0=1.83483438589289e-11 palpha0=-5.92157936193599e-18
+  alpha1=0.0
+  beta0=36.96
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.4352762 lkt1=2.72856796722e-8
+  kt2=-0.019151
+  at=2254.12799999997 lat=0.015279980616432
+  ute=-1.300713655 lute=6.82141991804604e-10
+  ua1=-1.192050637e-09 lua1=1.35432471052965e-15
+  ub1=6.82425623008204e-18 lub1=-3.34890091489061e-24 wub1=-5.26959356502109e-24 pub1=1.70066120083282e-30
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=1.81e-6
+  sbref=1.81e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.48 nmos
* DC IV MOS Parameters
+  lmin=2.0e-05 lmax=1.0e-04 wmin=1.5e-06 wmax=3.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.796161967949333+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} wvth0=5.82465134725489e-9
+  k1=0.88325
+  k2=-0.040337165352 wk2=8.00175386424651e-9
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=39808.2731413333 wvsat=0.114736911102664
+  ua=-1.48608538959733e-10 wua=-1.26987623332263e-18
+  ub=1.86201551506133e-18 wub=-3.41011234581363e-25
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.04215561309632 wu0=-4.34746924719019e-9
+  a0=0.749243386399547 wa0=6.45068589645414e-7
+  keta=-0.0351905965626667 wketa=1.45932023687291e-8
+  a1=0.0
+  a2=0.65972622
+  ags=0.157906297991467 wags=-3.83819565288392e-9
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.930480752133333+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} wnfactor=1.13816754513992e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=1.36005000637333 wpclm=-1.38315171925496e-6
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.4467e-5
+  alpha1=0.0
+  beta0=20.8954605333333 wbeta0=8.72043825866772e-6
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.414748784 wkt1=3.60845721048317e-8
+  kt2=-0.019151
+  at=157268.248533333 wat=-0.131107278647556
+  ute=-1.414280796 wute=3.47314006509008e-7
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.49 nmos
* DC IV MOS Parameters
+  lmin=8e-06 lmax=2.0e-05 wmin=1.5e-06 wmax=3.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.796161967949334+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} wvth0=5.82465134725531e-9
+  k1=0.88325
+  k2=-0.040337165352 wk2=8.00175386424651e-9
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=39808.2731413333 wvsat=0.114736911102664
+  ua=-1.48608538959733e-10 wua=-1.26987623332273e-18
+  ub=1.86201551506133e-18 wub=-3.41011234581364e-25
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.04215561309632 wu0=-4.34746924719017e-9
+  a0=0.749243386399546 wa0=6.45068589645415e-7
+  keta=-0.0351905965626667 wketa=1.45932023687292e-8
+  a1=0.0
+  a2=0.65972622
+  ags=0.157906297991467 wags=-3.83819565288392e-9
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.930480752133334+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} wnfactor=1.13816754513991e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=1.36005000637333 wpclm=-1.38315171925497e-6
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.4467e-5
+  alpha1=0.0
+  beta0=20.8954605333333 wbeta0=8.72043825866774e-6
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.414748784 wkt1=3.60845721048317e-8
+  kt2=-0.019151
+  at=157268.248533333 wat=-0.131107278647556
+  ute=-1.414280796 wute=3.47314006509008e-7
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.50 nmos
* DC IV MOS Parameters
+  lmin=4e-06 lmax=8e-06 wmin=1.5e-06 wmax=3.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.792552398370418+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=2.82366918416435e-08 wvth0=1.12474809849996e-08 pvth0=-4.24213375149116e-14
+  k1=0.88325
+  k2=-0.0443484358379496 lk2=3.13790899798229e-08 wk2=1.40280780562719e-08 pk2=-4.71423130730071e-14
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=24444.16987803 lvsat=0.120189246885045 wvsat=0.137819140912082 pvsat=-1.80566074679253e-7
+  ua=-1.48487531343643e-10 lua=-9.46610029625242e-19 wua=-1.45167178334062e-18 pua=1.42213768478728e-24
+  ub=2.04925404641407e-18 lub=-1.46471666360753e-24 wub=-6.22308667682088e-25 pub=2.20051415013745e-30
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0427845428164322 lu0=-4.91994801834344e-09 wu0=-5.29234055434136e-09 pu0=7.39147406546218e-15
+  a0=0.748783553632681 la0=3.59714804017444e-09 wa0=6.45759418483049e-07 pa0=-5.4041681638619e-15
+  keta=-0.0351905965626667 wketa=1.45932023687291e-8
+  a1=0.0
+  a2=0.65972622
+  ags=0.16261576291107 lags=-3.68408772199924e-08 wags=-1.09134508559199e-08 pags=5.53478182097011e-14
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.0105913901646+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-6.26683971556982e-07 wnfactor=-6.53730231100917e-09 pnfactor=9.41497411300687e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=1.36005000637333 wpclm=-1.38315171925496e-6
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.55745467865354e-05 lalpha0=-8.66404058098122e-12 walpha0=-1.66392069965795e-12 palpha0=1.30164040387559e-17
+  alpha1=0.0
+  beta0=15.3481622933458 lbeta0=4.33950219081959e-05 wbeta0=1.70544106749165e-05 pbeta0=-6.51944243737342e-11
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.437703121544776 lkt1=1.79565607895983e-07 wkt1=7.05699752065509e-08 pkt1=-2.69770031891313e-13
+  kt2=-0.019151
+  at=259797.622899999 lat=-0.802059715268725 wat=-0.285142079168568 pat=1.20497280911454e-6
+  ute=-1.49079525448259 lute=5.98552026319943e-07 wute=4.62265350181406e-07 pute=-8.99233439637715e-13
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.51 nmos
* DC IV MOS Parameters
+  lmin=2e-06 lmax=4e-06 wmin=1.5e-06 wmax=3.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.814039318728968+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-5.39020247075175e-08 wvth0=-1.86276872865354e-08 pvth0=7.17833943669031e-14
+  k1=0.88325
+  k2=-0.0416045364057562 lk2=2.08899005594949e-08 wk2=5.40115726403674e-09 pk2=-1.41639155259853e-14
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=25656.7766350079 lvsat=0.115553777444336 wvsat=0.142911783663729 pvsat=-2.00033877997901e-7
+  ua=-1.4830393267259e-10 lua=-1.64845836101704e-18 wua=-3.08244945917678e-18 pua=7.65616206031499e-24
+  ub=1.67434946563874e-18 lub=-3.15573006356879e-26 wub=-2.57044056843893e-26 pub=-8.01434569332721e-32
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0412862290757887 lu0=8.07702365740615e-10 wu0=-4.21977105589111e-09 pu0=3.29132939408195e-15
+  a0=0.401233044200054 la0=1.33218925451407e-06 wa0=1.24899564307745e-06 pa0=-2.31141398424384e-12
+  keta=-0.027309549650734 lketa=-3.01271223426993e-08 wketa=-9.06844306521807e-09 pketa=9.04521055113584e-14
+  a1=0.0
+  a2=0.65972622
+  ags=0.199399120299584 lags=-1.77453757793143e-07 wags=-6.61169376036776e-08 pags=2.66375898308444e-13
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.926284842035236+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-3.04402716519862e-07 wnfactor=1.97739747098885e-07 pnfactor=1.60601201932954e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=1.36005000637333 wpclm=-1.38315171925496e-6
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.11958059778781e-05 lalpha0=8.07470764923814e-12 walpha0=6.49862247032318e-12 palpha0=-1.81868027759692e-17
+  alpha1=0.0
+  beta0=22.8060300707575 lbeta0=1.48855995615832e-05 wbeta0=2.93509639330062e-06 pbeta0=-1.12200839706584e-11
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.407134579 lkt1=6.27102926852491e-8
+  kt2=-0.019151
+  at=95552.6216666667 lat=-0.174195257459025 wat=0.0300704767540267
+  ute=-1.27184026728806 lute=-2.38453990833174e-07 wute=1.49201345459533e-07 pute=2.9752603619673e-13
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.52 nmos
* DC IV MOS Parameters
+  lmin=1e-06 lmax=2e-06 wmin=1.5e-06 wmax=3.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.778372980349092+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=1.11081159139711e-08 wvth0=3.07124582032825e-08 pvth0=-1.81504183618959e-14
+  k1=0.88325
+  k2=-0.0370837429359244 lk2=1.26497101574349e-08 wk2=-3.96230919357353e-09 pk2=2.90316505376118e-15
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=80830.3141159705 lvsat=0.0149872602981232 wvsat=0.0553841781021562 pvsat=-4.04945979850502e-8
+  ua=-1.50165656267154e-10 lua=1.74496294822505e-18 wua=2.01170896605923e-18 pua=-1.62911842027393e-24
+  ub=1.67256043883212e-18 lub=-2.82963860154129e-26 wub=-3.65960304094844e-26 pub=-6.02909549064711e-32
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0414867843109361 lu0=4.42144121425288e-10 wu0=-3.77648490531938e-09 pu0=2.48333798556425e-15
+  a0=1.12265679986659 la0=1.72278109242424e-08 wa0=-3.23247535131724e-08 pa0=2.40884235541804e-14
+  keta=-0.0711347726271313 lketa=4.97544701582924e-08 wketa=7.39227732146505e-08 pketa=-6.08185571296626e-14
+  a1=0.0
+  a2=0.65972622
+  ags=0.107130098106346 lags=-9.27215070184144e-09 wags=1.47651202252721e-07 pags=-1.23265917020149e-13
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.769856297530521+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.92755591662412e-08 wnfactor=2.48467942860789e-07 pnfactor=6.81373469436648e-14
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=1.95079735887845 lpclm=-1.07677351257901e-06 wpclm=-3.15678085155401e-06 ppclm=3.23284880194457e-12
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=2.03999974269822e-05 lalpha0=-8.70205743497871e-12 walpha0=-2.8533264471069e-11 palpha0=4.56669035406015e-17
+  alpha1=0.0
+  beta0=29.6982592420596 lbeta0=2.32291979194649e-06 wbeta0=-9.52922597998709e-06 pbeta0=1.14990228131267e-11
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.37273
+  kt2=-0.019151
+  at=-19774.07581592 lat=0.0360142891701077 wat=0.0548103901643438 pat=-4.50942071103007e-8
+  ute=-1.48827819646741 lute=1.56054132257828e-07 wute=5.69479953807531e-07 pute=-4.68528811876024e-13
+  ua1=3.0044e-9
+  ub1=-4.2465249544776e-18 lub1=9.00474599299911e-25 wub1=7.42197402309513e-25 pub1=-1.35282621330902e-30
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.81e-6
+  sbref=2.81e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.53 nmos
* DC IV MOS Parameters
+  lmin=8.0e-07 lmax=1e-06 wmin=1.5e-06 wmax=3.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.781745515415132+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=8.33342676655244e-09 wvth0=3.30791058207669e-08 pvth0=-2.00975327228765e-14
+  k1=0.88325
+  k2=-0.0264430990948728 lk2=3.89532260944269e-09 wk2=-7.60934975519792e-09 pk2=5.903698382067e-15
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=132130.850841691 lvsat=-0.0272192815827659 wvsat=-0.0349508946877917 pvsat=3.38268667864965e-8
+  ua=-1.38753039054786e-10 lua=-7.64455102352388e-18 wua=-1.04268983776454e-17 pua=8.60450943821939e-24
+  ub=1.31648529090036e-18 lub=2.64657676517634e-25 wub=4.13240958623141e-26 pub=-1.24398258314197e-31
+  uc=6.49659440235399e-11 luc=1.01858703156899e-18 wuc=3.71707488481302e-18 puc=-3.05815273705705e-24
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0372362186179289 lu0=3.93921628459876e-09 wu0=4.43671380818123e-10 pu0=-9.88715415885969e-16
+  a0=1.21021817167643 la0=-5.48116440662348e-08 wa0=-1.25307661423247e-08 pa0=7.80329653057541e-15
+  keta=-0.01066
+  a1=0.0
+  a2=0.65972622
+  ags=-0.104627703533545 lags=1.64947557199148e-07 wags=-8.94347869782957e-09 pags=5.56938143297816e-15
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.3129828502261+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-4.66122610992023e-07 wnfactor=-7.94884255699929e-07 pnfactor=9.2653554461772e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.689692470758196 lpclm=-3.92234268709418e-08 wpclm=1.30210333535066e-06 ppclm=-4.35613444031696e-13
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.52656073913924e-05 lalpha0=-4.47783558660792e-12 walpha0=-2.8944621565594e-12 palpha0=2.45730660735827e-17
+  alpha1=0.0
+  beta0=27.9134705980921 lbeta0=3.79132073778657e-06 wbeta0=4.45678642095024e-06 pbeta0=-7.70315550897992e-15
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.37895731 lkt1=5.12340098361016e-9
+  kt2=-0.019151
+  at=8431.72500000001 lat=0.012808502459025
+  ute=-1.4589532325 lute=1.31927575327958e-7
+  ua1=6.0953253185e-09 lua1=-2.54300007821482e-15
+  ub1=-1.07496047118238e-17 lub1=6.25075991114113e-24 wub1=1.38430808244559e-24 pub1=-1.88111057528806e-30
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.41e-6
+  sbref=2.41e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.54 nmos
* DC IV MOS Parameters
+  lmin=6e-07 lmax=8.0e-07 wmin=1.5e-06 wmax=3.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.781928197326944+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=8.21966507692823e-09 wvth0=3.65957440633712e-08 pvth0=-2.22874523723322e-14
+  k1=0.88325
+  k2=0.000911237264600392 lk2=-1.31390706260284e-08 wk2=-2.8619213196518e-08 pk2=1.89871916527436e-14
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=68614.0445328244 lvsat=0.0123346027267611 wvsat=0.0628160576515235 pvsat=-2.70556452107176e-8
+  ua=-1.54981435230088e-10 lua=2.46137435511848e-18 wua=1.17725956415233e-17 pua=-5.21980367183172e-24
+  ub=-3.2097659373646e-19 lub=1.2843559533994e-24 wub=2.58450354697674e-24 pub=-1.70811494108614e-30
+  uc=5.28667617651555e-11 luc=8.55312289851497e-18 wuc=4.00430305399089e-17 puc=-2.56794514281107e-23
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0368093991750178 lu0=4.20500998310225e-09 wu0=3.53100380526958e-09 pu0=-2.91129302389706e-15
+  a0=1.1222
+  keta=-0.01066
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.570252283461086+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-3.60126241988183e-09 wnfactor=4.24883904869925e-07 pnfactor=1.66948098217895e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.214818984948731 lpclm=2.56495013820672e-07 wpclm=-1.06335253591558e-06 ppclm=1.0374292561378e-12
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=-1.03218001983088e-05 lalpha0=1.14562363291343e-11 walpha0=1.04656042422083e-10 palpha0=-4.24019671931796e-17
+  alpha1=0.0
+  beta0=27.7488321840351 lbeta0=3.89384618201066e-06 wbeta0=1.38383795459792e-05 pbeta0=-5.84991202385135e-12
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.37073
+  kt2=-0.019151
+  at=9131.64300000004 lat=0.012372641822967
+  ute=-1.13718994 lute=-6.84444015738598e-8
+  ua1=2.0117e-9
+  ub1=3.71090209504428e-19 lub1=-6.74441557912535e-25 wub1=-3.26353585166856e-24 pub1=1.01324592564678e-30
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.02e-6
+  sbref=2.01e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.55 nmos
* DC IV MOS Parameters
+  lmin=5e-07 lmax=6e-07 wmin=1.5e-06 wmax=3.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.933882035449781+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-5.60159328665771e-08 wvth0=-9.00356520873894e-09 pvth0=-3.01121076442311e-15
+  k1=0.88325
+  k2=-0.0139257595891757 lk2=-6.8670121090348e-09 wk2=8.50694823894731e-09 pk2=3.29281230296799e-15
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=88185.4049455505 lvsat=0.00406118196812905 wvsat=-0.0211096774465513 pvsat=8.42236471302674e-9
+  ua=-1.47031238351019e-10 lua=-8.99420321767371e-19 wua=-1.32338992165188e-17 pua=5.35121690600349e-24
+  ub=3.235758758219e-18 lub=-2.19186338668085e-25 wub=-5.05417110541111e-24 pub=1.52098963339244e-30
+  uc=9.53545884226091e-11 luc=-9.40779855221711e-18 wuc=-8.75202108494439e-17 puc=2.82454851676519e-23
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0455109030782561 lu0=5.26614536582367e-10 wu0=-6.0795793005965e-09 pu0=1.15139838302881e-15
+  a0=1.1222
+  keta=-0.01066
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.0144051996922716+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=2.31372531148793e-07 wnfactor=1.64218557006719e-06 pnfactor=-3.47643052012611e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-0.673391306529668 lpclm=6.31969038547626e-07 wpclm=5.87917175277674e-06 ppclm=-1.89739097894539e-12
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=2.42394203250304e-05 lalpha0=-3.15386298391739e-12 walpha0=1.83938627594983e-11 palpha0=-5.93626972223563e-18
+  alpha1=0.0
+  beta0=36.96
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.4352762 lkt1=2.72856796722e-8
+  kt2=-0.019151
+  at=2254.12799999997 lat=0.015279980616432
+  ute=-1.300713655 lute=6.82141991804604e-10
+  ua1=-1.192050637e-09 lua1=1.35432471052965e-15
+  ub1=5.64284418623082e-18 lub1=-2.90297538824806e-24 wub1=-1.72258347798845e-24 pub1=3.61837587768613e-31
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=1.81e-6
+  sbref=1.81e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.56 nmos
* DC IV MOS Parameters
+  lmin=2.0e-05 lmax=1.0e-04 wmin=1e-06 wmax=1.5e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.792208657424+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} wvth0=1.17638995083681e-8
+  k1=0.88325
+  k2=-0.028938775816 wk2=-9.12259385838404e-9
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=124760.09888 wvsat=-0.0128902943921702
+  ua=-1.466700791344e-10 wua=-4.18211747499243e-18
+  ub=1.402449179472e-18 wub=3.494173305586e-25
+  uc=9.3383668368e-11 wuc=-4.08333204133281e-17
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.03898470082496 wu0=4.16344461863004e-10
+  a0=1.2875694210256 wa0=-1.63684451822969e-7
+  keta=-0.032772088744 wketa=1.09597619843709e-8
+  a1=0.0
+  a2=0.65972622
+  ags=0.17451138202 wags=-2.87848104329829e-8
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.76902432232+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} wnfactor=3.56380498931193e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-0.74019317336 wpclm=1.77214442133105e-6
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=-1.8305770208e-05 walpha0=4.92361057764484e-11
+  alpha1=0.0
+  beta0=26.166750864 wbeta0=8.01125772971351e-7
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.386720608 wkt1=-6.02350205241582e-9
+  kt2=-0.019151
+  at=-90375.6800000001 wat=0.24094008209664
+  ute=-1.2119676224 wute=4.33692147773948e-8
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.57 nmos
* DC IV MOS Parameters
+  lmin=8e-06 lmax=2.0e-05 wmin=1e-06 wmax=1.5e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.792208657424+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} wvth0=1.17638995083681e-8
+  k1=0.88325
+  k2=-0.028938775816 wk2=-9.12259385838401e-9
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=124760.09888 wvsat=-0.0128902943921703
+  ua=-1.466700791344e-10 wua=-4.18211747499243e-18
+  ub=1.402449179472e-18 wub=3.494173305586e-25
+  uc=9.3383668368e-11 wuc=-4.08333204133281e-17
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.03898470082496 wu0=4.16344461863031e-10
+  a0=1.2875694210256 wa0=-1.63684451822968e-7
+  keta=-0.032772088744 wketa=1.09597619843709e-8
+  a1=0.0
+  a2=0.65972622
+  ags=0.17451138202 wags=-2.87848104329829e-8
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.769024322319999+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} wnfactor=3.56380498931192e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-0.74019317336 wpclm=1.77214442133105e-6
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=-1.8305770208e-05 walpha0=4.92361057764484e-11
+  alpha1=0.0
+  beta0=26.166750864 wbeta0=8.0112577297131e-7
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.386720608 wkt1=-6.02350205241603e-9
+  kt2=-0.019151
+  at=-90375.68 wat=0.24094008209664
+  ute=-1.2119676224 wute=4.33692147773948e-8
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.58 nmos
* DC IV MOS Parameters
+  lmin=4e-06 lmax=8e-06 wmin=1e-06 wmax=1.5e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.78820643970024+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=3.13082726563984e-08 wvth0=1.77766233012224e-08 pvth0=-4.70359208087985e-14
+  k1=0.88325
+  k2=-0.0253312238897967 lk2=-2.82209082872203e-08 wk2=-1.45423922796117e-08 pk2=4.23976251234888e-14
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=124760.09888 wvsat=-0.0128902943921703
+  ua=-1.46902472150145e-10 lua=1.81794804845443e-18 wua=-3.83298229257352e-18 pua=-2.73119061469981e-24
+  ub=9.35521223895571e-19 lub=3.65265179285436e-24 wub=1.05090561076294e-24 pub=-5.48755411569116e-30
+  uc=9.3383668368e-11 wuc=-4.0833320413328e-17
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0378840085692306 lu0=8.61041943035447e-09 wu0=2.06996727087357e-09 pu0=-1.29358464103541e-14
+  a0=1.2922123001217 la0=-3.63199942343311e-08 wa0=-1.70659671947238e-07 pa0=5.45652706979584e-14
+  keta=-0.032772088744 wketa=1.09597619843709e-8
+  a1=0.0
+  a2=0.65972622
+  ags=0.127379472866241 lags=3.68700246826291e-07 wags=4.20237190203479e-08 pags=-5.53916078418985e-13
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.570637704179611+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.55192514771198e-06 wnfactor=6.54426237921171e-07 pnfactor=-2.3315316418148e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-0.74019317336 wpclm=1.77214442133105e-6
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=-3.57668579697721e-05 lalpha0=1.36593392527735e-10 walpha0=7.54687360531712e-11 palpha0=-2.05210810077258e-16
+  alpha1=0.0
+  beta0=28.320170070082 lbeta0=-1.68456191794135e-05 wbeta0=-2.43405926444762e-06 pbeta0=2.53079822829535e-11
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.382888901227612 lkt1=-2.99744113512698e-08 wkt1=-1.17800590584997e-08 pkt1=4.50319969447573e-14
+  kt2=-0.019151
+  at=-301119.55248134 lat=1.64859262431983 wat=0.557550717431236 pat=-2.47675983196164e-6
+  ute=-1.2119676224 wute=4.33692147773956e-8
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.59 nmos
* DC IV MOS Parameters
+  lmin=2e-06 lmax=4e-06 wmin=1e-06 wmax=1.5e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.795270009468324+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=4.30614553328502e-09 wvth0=9.57034694257454e-09 pvth0=-1.5665533778026e-14
+  k1=0.88325
+  k2=-0.0353667058430187 lk2=1.01420396753019e-08 wk2=-3.97023500623083e-09 pk2=1.98311177766038e-15
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=135117.578588022 lvsat=-0.0395938587617275 wvsat=-0.0215364332287783 pvsat=3.30518629610057e-8
+  ua=-1.4764682457355e-10 lua=4.66340713232725e-18 wua=-4.06965449755442e-18 pua=-1.82645643988027e-24
+  ub=2.23149945195267e-18 lub=-1.3015243548646e-24 wub=-8.62737573323145e-25 pub=1.82778900705342e-30
+  uc=1.17428957143398e-10 luc=-9.19186708056678e-17 wuc=-7.69577119144704e-17 puc=1.38093831247553e-22
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0418318844241591 lu0=-6.4812479844325e-09 wu0=-5.03953527720469e-09 pu0=1.42418693747639e-14
+  a0=1.44086346683731 la0=-6.04573417424254e-07 wa0=-3.12891043110788e-07 pa0=5.98277542417362e-13
+  keta=-0.056415229479798 lketa=9.03813670280978e-08 wketa=3.46584168146165e-08 pketa=-9.05935824778797e-14
+  a1=0.0
+  a2=0.65972622
+  ags=0.245315286636944 lags=-8.21366444852025e-08 wags=-1.35098998268279e-07 pags=1.23176423764486e-13
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.12983943215205+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-5.85752633061822e-07 wnfactor=-1.08070084253928e-07 pnfactor=5.83286686349932e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-0.740193173360001 wpclm=1.77214442133105e-6
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=-9.02542620708921e-06 lalpha0=3.43680923441428e-11 walpha0=3.68779502009445e-11 palpha0=-5.76886166855899e-17
+  alpha1=0.0
+  beta0=20.7837913976754 lbeta0=1.19639291993343e-05 wbeta0=5.9732026193281e-06 pbeta0=-6.83071834527452e-12
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.407134579 lkt1=6.27102926852496e-8
+  kt2=-0.019151
+  at=230519.47817164 lat=-0.383720378967271 wat=-0.172696710182507 pat=3.14779647247671e-7
+  ute=-1.1802024576403 lute=-1.21429680047017e-07 wute=1.15294654108392e-08 pute=1.21714796935766e-13
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.60 nmos
* DC IV MOS Parameters
+  lmin=1e-06 lmax=2e-06 wmin=1e-06 wmax=1.5e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.796019009055702+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=2.94092076638461e-09 wvth0=4.20198226796447e-09 pvth0=-5.88044906630961e-15
+  k1=0.88325
+  k2=-0.0364117836669904 lk2=1.20469354224677e-08 wk2=-4.97182585733798e-09 pk2=3.80874247128966e-15
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=129163.93639985 lvsat=-0.0287419705824383 wvsat=-0.0172297426687857 pvsat=2.52019245698997e-8
+  ua=-1.45296124319302e-10 lua=3.7871290720167e-19 wua=-5.30402261673255e-18 pua=4.23464596357483e-25
+  ub=1.5052171686533e-18 lub=2.22928776559645e-26 wub=2.14811796857124e-25 pub=-1.36293634004635e-31
+  uc=3.48973919084798e-11 luc=5.85141716265406e-17 wuc=4.70334200530791e-17 puc=-8.79086487147901e-23
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0365322403897227 lu0=3.17857748609983e-09 wu0=3.66696424562757e-09 pu0=-1.62773720698782e-15
+  a0=1.08088450784044 la0=5.15713904870688e-08 wa0=3.04317658677358e-08 pa0=-2.75075845148699e-14
+  keta=-0.00367810815684387 lketa=-5.7442188580117e-09 wketa=-2.74206117389569e-08 pketa=2.25597873166038e-14
+  a1=0.0
+  a2=0.65972622
+  ags=0.280197298357686 lags=-1.45717168590961e-07 wags=-1.12355959910479e-07 pags=8.1721982715534e-14
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.751966009699182+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.03008968119112e-07 wnfactor=2.75345381003625e-07 pnfactor=-1.15576568054434e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-2.51243523087537 lpclm=3.23032053773704e-06 wpclm=3.54854770319746e-06 ppclm=-3.23790533035965e-12
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=-3.0275611234253e-06 lalpha0=2.3435597722331e-11 walpha0=6.66308126201857e-12 palpha0=-2.61503840967236e-18
+  alpha1=0.0
+  beta0=20.6550487354105 lbeta0=1.2198592440867e-05 wbeta0=4.05682323825611e-06 pbeta0=-3.33767423963368e-12
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.37273
+  kt2=-0.019151
+  at=16709.076 lat=0.00599846919344399
+  ute=-0.861492961059723 lute=-7.02351359458826e-07 wute=-3.72169591036734e-07 pute=8.21094961793507e-13
+  ua1=3.0044e-9
+  ub1=-3.00980870718737e-18 lub1=-1.35372644283967e-24 wub1=-1.11578077837448e-24 pub1=2.03376821394728e-30
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.81e-6
+  sbref=2.81e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.61 nmos
* DC IV MOS Parameters
+  lmin=8.0e-07 lmax=1e-06 wmin=1e-06 wmax=1.5e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.811828988608955+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-1.00664395214428e-08 wvth0=-1.21167399650264e-08 pvth0=7.54546959516161e-15
+  k1=0.88325
+  k2=-0.0305704289907948 lk2=7.24107184836665e-09 wk2=-1.40866394071927e-09 pk2=8.77218704468062e-16
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=72169.177208734 lvsat=0.0181493846416279 wvsat=0.0551324057713347 pvsat=-3.4332658178389e-8
+  ua=-1.32579570725209e-10 lua=-1.00835899478199e-17 wua=-1.97015961756481e-17 pua=1.22687946880577e-23
+  ub=1.20940666709628e-18 lub=2.65665347412466e-25 wub=2.0219345217712e-25 pub=-1.2591213066771e-31
+  uc=2.3122639425898e-10 luc=-1.03011784806289e-16 wuc=-2.46063980005501e-16 puc=1.53231668332805e-22
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0329081478992339 lu0=6.16023072489216e-09 wu0=6.94593976890822e-09 pu0=-4.32545201823193e-15
+  a0=1.21009927153571 la0=-5.47376012627047e-08 wa0=-1.23521367537137e-08 pa0=7.69205847277619e-15
+  keta=-0.01066
+  a1=0.0
+  a2=0.65972622
+  ags=-0.0749140393292189 lags=1.46443937375524e-07 wags=-5.35837426878701e-08 pags=3.33682576677601e-14
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.414604233074654+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=3.80566959963188e-07 wnfactor=5.54793063020306e-07 pnfactor=-3.45486838927698e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=2.61609633001858 lpclm=-9.89081361888799e-07 wpclm=-1.59202564980146e-06 ppclm=9.91403724926515e-13
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=3.79763348847082e-06 lalpha0=1.78202985340911e-11 walpha0=1.43344255005471e-11 palpha0=-8.92649112638115e-18
+  alpha1=0.0
+  beta0=30.88001791 lbeta0=3.78619332688779e-6
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.37895731 lkt1=5.12340098361016e-9
+  kt2=-0.019151
+  at=8431.72500000003 lat=0.012808502459025
+  ute=-3.17260247352226 lute=1.19907008083899e-06 wute=2.57449750995131e-06 pute=-1.60321940886949e-12
+  ua1=6.0953253185e-09 lua1=-2.54300007821482e-15
+  ub1=-1.35416314655632e-17 lub1=7.31113062698161e-24 wub1=5.57890389187236e-24 pub1=-3.47415639948957e-30
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.41e-6
+  sbref=2.41e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.62 nmos
* DC IV MOS Parameters
+  lmin=6e-07 lmax=8.0e-07 wmin=1e-06 wmax=1.5e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.80628723003+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-6.61541465981143e-9
+  k1=0.88325
+  k2=-0.01813841913759 lk2=-5.00726079529443e-10
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=110425.966705 lvsat=-0.00567430413817138
+  ua=-1.471453042927e-10 lua=-1.01305611760265e-18
+  ub=1.3993329131e-18 lub=1.47392386312324e-25
+  uc=7.95203936399999e-11 luc=-8.53975533483086e-18
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.03915972267215 lu0=2.26718131497936e-9
+  a0=1.1222
+  keta=-0.01066
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.853065523050001+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.07523522395551e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-0.4929747725 lpclm=9.47033594853697e-7
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=5.9339851045e-05 lalpha0=-1.67675621471039e-11
+  alpha1=0.0
+  beta0=36.96
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.37073
+  kt2=-0.019151
+  at=9131.64299999998 lat=0.012372641822967
+  ute=-1.13718994 lute=-6.84444015738594e-8
+  ua1=2.0117e-9
+  ub1=-1.8012e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.02e-6
+  sbref=2.01e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.63 nmos
* DC IV MOS Parameters
+  lmin=5e-07 lmax=6e-07 wmin=1e-06 wmax=1.5e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.925540511192462+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-5.70274734589009e-08 wvth0=3.5283070761935e-09 pvth0=-1.4915247786269e-15
+  k1=0.88325
+  k2=0.0130597615589074 lk2=-1.36891642035405e-08 wk2=-3.2034695486833e-08 pk2=1.35420588578444e-14
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=96765.5558562644 lvsat=0.000100375000325392 wvsat=-0.0340000500069608 pvsat=1.43728751394926e-8
+  ua=-1.33142135900223e-10 lua=-6.9326294953226e-18 wua=-3.41001645052665e-17 pua=1.44151966414756e-23
+  ub=-1.5280938005684e-18 lub=1.38490640840808e-24 wub=2.10279325857802e-24 pub=-8.88915896991946e-31
+  uc=-9.13972395179613e-11 luc=6.37124266476674e-17 wuc=1.93046024353417e-16 puc=-8.16065389209441e-23
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0441029472885234 lu0=1.77527029675238e-10 wu0=-3.96433973580302e-09 pu0=1.67584930085575e-15
+  a0=1.1222
+  keta=-0.01066
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.60643362873125+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-2.10948530287191e-07 wnfactor=-7.49595156242661e-07 pnfactor=3.16877109993616e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=3.239930875 lpclm=-6.30981342419626e-7
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=3.648283048e-05 lalpha0=-7.10519098664088e-12
+  alpha1=0.0
+  beta0=36.96
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.4352762 lkt1=2.72856796722002e-8
+  kt2=-0.019151
+  at=-54058.7974973031 lat=0.0390851999248324 wat=0.0846016109950224 pat=-3.57637236175368e-8
+  ute=-0.292722640238988 lute=-4.25426907669131e-07 wute=-1.51435328504417e-06 pute=6.40164078540008e-13
+  ua1=-1.19205063700001e-09 lua1=1.35432471052965e-15
+  ub1=1.73911594479305e-17 lub1=-8.1132053017831e-24 wub1=-1.93726414147724e-23 pub1=8.18941607790815e-30
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=1.81e-6
+  sbref=1.81e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.64 nmos
* DC IV MOS Parameters
+  lmin=2.0e-05 lmax=1.0e-04 wmin=7.5e-07 wmax=1.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.808702848752+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} wvth0=-4.76902018087055e-9
+  k1=0.88325
+  k2=-0.032620085008 wk2=-5.43264095240124e-9
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=144702.3728 wvsat=-0.0328793927713344
+  ua=-1.521420059352e-10 wua=1.3026574099359e-18
+  ub=2.403117039776e-18 wub=-6.53600097881393e-25
+  uc=3.9537088448e-11 wuc=1.31396912763241e-17
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.040014738316 wu0=-6.16111557205976e-10
+  a0=2.0761041806528 wa0=-9.54070691065773e-7
+  keta=-0.026604876928 wketa=4.77806955502695e-9
+  a1=0.0
+  a2=0.65972622
+  ags=0.102290229248 wags=4.36059176057256e-8
+  b0=-3.080311136e-07 wb0=3.41764697338733e-13
+  b1=9.79346438559999e-11 wb1=-9.81645943997738e-17
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.18180863584+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} wnfactor=-5.73730321569527e-8
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=3.50221238416 wpclm=-2.48022230443801e-6
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=3.9087818608e-05 walpha0=-8.2922431860916e-12
+  alpha1=0.0
+  beta0=21.66947008 wbeta0=5.30896617225215e-6
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.398748784 wkt1=6.03291610483197e-9
+  kt2=-0.019151
+  at=420845.28 wat=-0.27148122471744
+  ute=-1.277038112 wute=1.08592489886977e-7
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.65 nmos
* DC IV MOS Parameters
+  lmin=8e-06 lmax=2.0e-05 wmin=7.5e-07 wmax=1.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.811804462995799+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-6.14824648205887e-08 wvth0=-7.87791701491265e-09 pvth0=6.16268256479819e-14
+  k1=0.88325
+  k2=-0.0290868735892264 lk2=-7.00378995204777e-08 wk2=-8.97414835158611e-09 pk2=7.02023485085515e-14
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=166086.051014676 lvsat=-0.423882901040091 wvsat=-0.0543132798624588 pvsat=4.24878178091733e-7
+  ua=-1.52989211571623e-10 lua=1.67939294324928e-17 wua=2.15185228519289e-18 pua=-1.68333615787999e-23
+  ub=2.82819709740899e-18 lub=-8.42624763592337e-24 wub=-1.07967824348971e-24 pub=8.44603246537252e-30
+  uc=3.09914643834926e-11 luc=1.69397607057856e-16 wuc=2.1705380466135e-17 puc=-1.69795352639228e-22
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0404154370568576 lu0=-7.94294335205864e-09 wu0=-1.01775113870711e-09 pu0=7.96159338304928e-15
+  a0=2.69660045300462 la0=-1.22999306933329e-05 wa0=-1.57602388866508e-06 pa0=1.23288109306009e-11
+  keta=-0.0297123765878209 lketa=6.15991298392204e-08 wketa=7.89286562404907e-09 pketa=-6.1743764596083e-14
+  a1=0.0
+  a2=0.65972622
+  ags=0.0739303712414532 lags=5.62169836461978e-07 wags=7.2032364558872e-08 pags=-5.6348981123799e-13
+  b0=-5.30303658712187e-07 lb0=4.40604887044425e-12 wb0=5.64559138386843e-13 pb0=-4.41639427319205e-18
+  b1=1.61777675061524e-10 lb1=-1.26554323381171e-15 wb1=-1.62157529042569e-16 pb1=1.2685147293247e-21
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.21912217342194+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-7.39656218145193e-07 wnfactor=-9.47741819251351e-08 pnfactor=7.41392930945391e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=5.1152675895227 lpclm=-3.19751594240545e-05 wpclm=-4.09706496342289e-06 ppclm=3.20502370983822e-11
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=4.44808214898482e-05 lalpha0=-1.06904045409102e-10 walpha0=-1.36979088387064e-11 palpha0=1.07155056107723e-16
+  alpha1=0.0
+  beta0=18.2166926801991 lbeta0=6.84434775991337e-05 wbeta0=8.76985069338783e-06 pbeta0=-6.86041828845365e-11
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.402672394681592 lkt1=7.77766790899245e-08 wkt1=9.96573942430446e-09 pkt1=-7.79592987324291e-14
+  kt2=-0.019151
+  at=597407.76067164 lat=-3.49995055904662 wat=-0.448458274093697 pat=3.50816844295926e-6
+  ute=-1.34766310426866 lute=1.39998022361865e-06 wute=1.79383309637479e-07 pute=-1.4032673771837e-12
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.66 nmos
* DC IV MOS Parameters
+  lmin=4e-06 lmax=8e-06 wmin=7.5e-07 wmax=1.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.807402441468123+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-2.70466345533712e-08 wvth0=-1.46445067880999e-09 pvth0=1.14560037231033e-14
+  k1=0.88325
+  k2=-0.0504348231167274 lk2=9.69613670347398e-08 wk2=1.06201501983038e-08 pk2=-8.30785781809274e-14
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=80551.3381559709 lvsat=0.245232148815804 wvsat=0.031422268502039 pvsat=-2.45807953901224e-7
+  ua=-1.49135602994441e-10 lua=-1.33518138460927e-17 wua=-1.59460805705536e-18 pua=1.24741898807765e-23
+  ub=2.06173277802987e-18 lub=-2.43040344432239e-24 wub=-7.79502881004715e-26 pub=6.09784135182482e-31
+  uc=6.51739606415222e-11 luc=-9.80028660772151e-17 wuc=-1.25573762931084e-17 puc=9.82329768067643e-23
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0410140266048861 lu0=-1.26255483656968e-08 wu0=-1.06740004712962e-09 pu0=8.3499834380824e-15
+  a0=0.205329605405133 la0=7.18861099557992e-06 wa0=9.18775023336525e-07 pa0=-7.18732985708037e-12
+  keta=-0.0172823779485374 lketa=-3.56374058462599e-08 wketa=-4.56631865203943e-09 pketa=3.5721082475187e-14
+  a1=0.0
+  a2=0.65972622
+  ags=0.281633621575158 lags=-1.06263681872426e-06 wags=-1.12592618429737e-07 pags=8.80781766561477e-13
+  b0=3.5878652173656e-07 lb0=-2.54906444594776e-12 wb0=-3.26618625805597e-13 pb0=2.55504964926685e-18
+  b1=-9.35944497605726e-11 lb1=7.32164203569974e-16 wb1=9.38142095286104e-17 pb1=-7.33883325119956e-22
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.46664125937496+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-2.67593144492152e-06 wnfactor=-2.43681133621775e-07 pnfactor=1.9062519580982e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-1.33695323192808 lpclm=1.8498828414754e-05 wpclm=2.37030567251665e-06 ppclm=-1.85422636638719e-11
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=5.78309854859996e-05 lalpha0=-2.11338787156879e-10 walpha0=-1.83488751390347e-11 palpha0=1.43538314365256e-16
+  alpha1=0.0
+  beta0=27.7209638672388 lbeta0=-5.90587924812868e-06 wbeta0=-1.83344612544005e-06 pbeta0=1.43425558423099e-11
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.394641365500001 lkt1=1.49520981491815e-8
+  kt2=-0.019151
+  at=312645.58294776 lat=-1.27233264373851 wat=-0.0576555385358514 pat=4.51023768626098e-7
+  ute=-1.06516313519403 lute=-8.09941041960453e-07 wute=-1.03779969364533e-07 pute=8.11842783526978e-13
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.67 nmos
* DC IV MOS Parameters
+  lmin=2e-06 lmax=4e-06 wmin=7.5e-07 wmax=1.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.810093696386089+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-3.73345781571817e-08 wvth0=-5.28814599207406e-09 pvth0=2.60729623316669e-14
+  k1=0.88325
+  k2=-0.0255642081467986 lk2=1.88769620012919e-09 wk2=-1.37957489670416e-08 pk2=1.02568364513127e-14
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=179071.574182834 lvsat=-0.131384211571404 wvsat=-0.0655936328052471 pvsat=1.25057739519079e-7
+  ua=-1.54160957669918e-10 lua=5.85876525784815e-18 wua=2.45977378332423e-18 pua=-3.0246212662794e-24
+  ub=1.31364299036314e-18 lub=4.29342577774629e-25 wub=5.72740152381968e-26 pub=9.28579988563541e-32
+  uc=-8.55348910279702e-12 luc=1.83837341611336e-16 wuc=4.93205411155111e-17 puc=-1.38309656286605e-22
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0373124883548525 lu0=1.52443665039237e-09 wu0=-5.09527665927325e-10 pu0=6.21738739241654e-15
+  a0=1.72456767343709 la0=1.38097253653403e-06 wa0=-5.97261387187664e-07 pa0=-1.39193047344082e-12
+  keta=-0.026604876928 wketa=4.77806955502692e-9
+  a1=0.0
+  a2=0.65972622
+  ags=-0.0390859133532448 lags=1.63387689752131e-07 wags=1.49969975739487e-07 pags=-1.22924401609636e-13
+  b0=-4.36113150891039e-07 lb0=4.89623174495612e-13 wb0=4.70147471253331e-13 pb0=-4.90772809709328e-19
+  b1=2.83955290092932e-10 lb1=-7.11106891009954e-16 wb1=-2.8462201711407e-16 pb1=7.12776569990046e-22
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.565641978592248+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=7.68346436704248e-07 wnfactor=4.57452104926832e-07 pnfactor=-7.73991808031948e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=3.50221238416 wpclm=-2.48022230443801e-6
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=2.68637333004843e-05 lalpha0=-9.29593122424921e-11 walpha0=9.04522946847233e-13 palpha0=6.99377526470145e-17
+  alpha1=0.0
+  beta0=27.6265376446715 lbeta0=-5.54491319990785e-06 wbeta0=-8.8561039585596e-07 pbeta0=1.07192348159211e-11
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.407134579 lkt1=6.27102926852487e-8
+  kt2=-0.019151
+  at=-56813.65089552 lat=0.140010622710442 wat=0.115311077071703 pat=-2.10181074821982e-7
+  ute=-1.37577372961194 lute=3.77439706249293e-07 wute=2.07559938729065e-07 pute=-3.78325934679567e-13
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.68 nmos
* DC IV MOS Parameters
+  lmin=1e-06 lmax=2e-06 wmin=7.5e-07 wmax=1.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.768474749470466+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=3.8525566573279e-08 wvth0=3.18109157747067e-08 pvth0=-4.15486476215581e-14
+  k1=0.88325
+  k2=-0.0293014148413765 lk2=8.69961869574382e-09 wk2=-1.20988898289544e-08 pk2=7.1639186976879e-15
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=103765.730211941 lvsat=0.00587808471550688 wvsat=0.00822809850725281 pvsat=-9.499418617885e-9
+  ua=-1.50611637252012e-10 lua=-6.10691096803309e-19 wua=2.39711403433281e-20 pua=1.41519172096362e-24
+  ub=1.63301466910097e-18 lub=-1.52786081582842e-25 wub=8.67142278784027e-26 pub=3.91964106304618e-32
+  uc=1.5650964136704e-10 luc=-1.17028343253081e-16 wuc=-7.48643749672099e-17 puc=8.8046039989769e-23
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0384824954043378 lu0=-6.08171468923196e-10 wu0=1.71213003223818e-09 pu0=2.16790303458163e-15
+  a0=3.54052395048844 la0=-1.92902726429206e-06 wa0=-2.43498291019161e-06 pa0=1.95774151590568e-12
+  keta=-0.0397232214678504 lketa=2.3911213261466e-08 wketa=8.7091354981038e-09 pketa=-7.16527575749044e-15
+  a1=0.0
+  a2=0.65972622
+  ags=0.191741898815005 lags=-2.57349319149115e-07 wags=-2.3692867089671e-08 pags=1.93616245563198e-13
+  b0=-3.95864753737438e-08 lb0=-2.33138289296704e-13 wb0=7.26897511019213e-14 pb0=2.33685697999973e-19
+  b1=5.83311906154261e-10 lb1=-1.25675347516004e-15 wb1=-5.84681522509911e-16 pb1=1.25970433231971e-21
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.984020528881793+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=5.75488335643733e-09 wnfactor=4.27459978099756e-08 pnfactor=-1.80941307007336e-14
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=6.1742996224072 lpclm=-4.87049624385756e-06 wpclm=-5.15858360352061e-06 ppclm=4.88193216903814e-12
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=-6.99479501716981e-05 lalpha0=8.35023443844425e-11 walpha0=7.37405993837767e-11 palpha0=-6.28228217929465e-17
+  alpha1=0.0
+  beta0=15.6186920457019 lbeta0=1.63421592165476e-05 wbeta0=9.10500529347218e-06 pbeta0=-7.49097011010365e-12
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.37273
+  kt2=-0.019151
+  at=16709.076 lat=0.00599846919344402
+  ute=-1.7472869395089 lute=1.05460835083801e-06 wute=5.15704231673847e-07 pute=-9.39990089903103e-13
+  ua1=3.0044e-9
+  ub1=-4.49510655875966e-18 lub1=1.35357199545456e-24 wub1=3.73004552553316e-25 pub1=-6.79886961080058e-31
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.81e-6
+  sbref=2.81e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.69 nmos
* DC IV MOS Parameters
+  lmin=8.0e-07 lmax=1e-06 wmin=7.5e-07 wmax=1.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.774721653570436+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=3.33860449162044e-08 wvth0=2.50777230961617e-08 pvth0=-3.60090412759464e-14
+  k1=0.88325
+  k2=-0.0306768302821886 lk2=9.83121561677868e-09 wk2=-1.30201281909329e-09 pk2=-1.71900672151221e-15
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=169603.386799398 lvsat=-0.0482885963263484 wvsat=-0.0425305793434483 pvsat=3.22613191688999e-8
+  ua=-1.71471912808448e-10 lua=1.6551704272019e-17 wua=1.92820651268025e-17 pua=-1.44290392026096e-23
+  ub=1.25457791138648e-18 lub=1.58565570528353e-25 wub=1.56916145805325e-25 pub=-1.85608835074709e-32
+  uc=-2.0023459379401e-10 luc=1.76476198085205e-16 wuc=1.86410078447438e-16 puc=-1.26912552342518e-22
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0333562083091468 lu0=3.60938383919048e-09 wu0=6.49682731315283e-09 pu0=-1.76861574404258e-15
+  a0=1.42521408908625 la0=-1.88696266710766e-07 wa0=-2.27972043895858e-07 pa0=1.41965258867311e-13
+  keta=0.0472741247908106 lketa=-4.76642004232684e-08 wketa=-5.80701541158193e-08 pketa=4.77761159658622e-14
+  a1=0.0
+  a2=0.65972622
+  ags=-0.996949788725737 lags=7.20624181632967e-07 wags=8.70616946648231e-07 pags=-5.421601618032e-13
+  b0=-1.4310785489521e-06 lb0=9.11685375890489e-13 wb0=1.46744904806904e-12 pb0=-9.1382601315308e-19
+  b1=-3.88422343648918e-09 lb1=2.41882634482834e-15 wb1=3.89334359311805e-15 pb1=-2.424505749086e-21
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.48711708308097+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-4.08158247776411e-07 wnfactor=-5.20238047157829e-07 pnfactor=4.45090295599674e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-1.43131424375202 lpclm=1.38687805786148e-06 wpclm=2.46488824399635e-06 ppclm=-1.39013444754134e-12
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=2.773828919182e-05 lalpha0=3.13284698665589e-12 walpha0=-9.66244286239364e-12 palpha0=5.79544655728748e-18
+  alpha1=0.0
+  beta0=30.88001791 lbeta0=3.78619332688774e-6
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.378957310000001 lkt1=5.12340098361059e-9
+  kt2=-0.019151
+  at=8431.72499999998 lat=0.012808502459025
+  ute=1.96834524954453 lute=-2.00235743569411e-06 wute=-2.57852115836924e-06 pute=1.60572505947243e-12
+  ua1=6.0953253185e-09 lua1=-2.54300007821482e-15
+  ub1=-6.11514220770167e-18 lub1=2.68642554494427e-24 wub1=-1.86502276276659e-24 pub1=1.1614074900804e-30
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.41e-6
+  sbref=2.41e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.70 nmos
* DC IV MOS Parameters
+  lmin=6e-07 lmax=8.0e-07 wmin=7.5e-07 wmax=1.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.837252490774+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-5.55384586640858e-09 wvth0=-3.1037967176229e-08 pvth0=-1.06406135693082e-15
+  k1=0.88325
+  k2=-0.00530596074401637 lk2=-5.96801134159689e-09 wk2=-1.28625890058817e-08 pk2=5.48012244786277e-15
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=154253.099561557 lvsat=-0.0387294966044405 wvsat=-0.0439300389645044 pvsat=3.31328060581799e-8
+  ua=-1.24787343635771e-10 lua=-1.25202241734516e-17 wua=-2.2410457148552e-17 pua=1.1534186886444e-23
+  ub=2.04765559675248e-18 lub=-3.35308489557303e-25 wub=-6.49844945313701e-25 pub=4.83834257526168e-31
+  uc=1.68689517031658e-10 luc=-5.32642823733743e-17 wuc=-8.93784924933818e-17 puc=4.48295402280299e-23
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0341118594669004 lu0=3.13881643807134e-09 wu0=5.05971558805553e-09 pu0=-8.73681722361004e-16
+  a0=1.1222
+  keta=-0.0292664688576 wketa=1.86501568464776e-8
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.606861232018368+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.40004358611658e-07 wnfactor=2.46782378706974e-07 pnfactor=-3.25571012195421e-14
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-5.30160632986333 lpclm=3.79702891893766e-06 wpclm=4.81992222426001e-06 ppclm=-2.85668711310491e-12
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=5.8556373156851e-05 lalpha0=-1.60585292589718e-11 walpha0=7.85317494230447e-13 palpha0=-7.10697697353413e-19
+  alpha1=0.0
+  beta0=34.6701060788064 lbeta0=1.4259879314388e-06 wbeta0=2.29527059212057e-06 pbeta0=-1.42933615110183e-12
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.37073
+  kt2=-0.019151
+  at=9131.64299999998 lat=0.012372641822967
+  ute=-1.13718994 lute=-6.84444015738594e-8
+  ua1=2.0117e-9
+  ub1=-1.8012e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.02e-6
+  sbref=2.01e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.71 nmos
* DC IV MOS Parameters
+  lmin=5e-07 lmax=6e-07 wmin=7.5e-07 wmax=1.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={1.02032486314634+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-8.29442129117407e-08 wvth0=-9.14785985360731e-08 pvth0=2.44860671784477e-14
+  k1=0.88325
+  k2=-0.00522767670481988 lk2=-6.00110443177043e-09 wk2=-1.37043183180624e-08 pk2=5.83594752173023e-15
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=-60262.8507423664 lvsat=0.0519530455834875 wvsat=0.123397059290363 pvsat=-3.76015455141986e-8
+  ua=-2.00831595879396e-10 lua=1.96260386217487e-17 wua=3.37482303259377e-17 pua=-1.22058312283345e-23
+  ub=-1.37147325068622e-18 lub=1.11006326724931e-24 wub=1.94580496364471e-24 pub=-6.13427424137732e-31
+  uc=-5.01226823710712e-11 luc=3.9234417492341e-17 wuc=1.51674554546345e-16 puc=-5.70710554001211e-23
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0333884482263436 lu0=3.44462479520319e-09 wu0=6.77531697017472e-09 pu0=-1.59891961022562e-15
+  a0=1.1222
+  keta=-0.089315311866421 lketa=2.53845074539619e-08 wketa=7.88399945386834e-08 pketa=-2.54441102774638e-14
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={-0.145055675685168+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=4.57862944922081e-07 wnfactor=1.00600664506053e-06 pnfactor=-3.53504734559446e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=11.412307847082 lpclm=-3.26846073499664e-06 wpclm=-8.1915657132125e-06 ppclm=2.64367219419078e-12
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=4.02611554499695e-05 lalpha0=-8.3245735825241e-12 walpha0=-3.78719647699893e-12 palpha0=1.22224570621835e-18
+  alpha1=0.0
+  beta0=41.5397878423872 lbeta0=-1.47803951016146e-06 wbeta0=-4.59054118424109e-06 pbeta0=1.48150994693133e-12
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.435276200000001 lkt1=2.72856796721998e-8
+  kt2=-0.019151
+  at=30344.6342399999 lat=0.00340525282309057
+  ute=-1.803528553 lute=2.13237586638243e-7
+  ua1=-1.192050637e-09 lua1=1.35432471052965e-15
+  ub1=-4.26606814883525e-18 lub1=1.04197617742527e-24 wub1=2.33543735239053e-24 pub1=-9.87261767413401e-31
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=1.81e-6
+  sbref=1.81e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.72 nmos
* DC IV MOS Parameters
+  lmin=2.0e-05 lmax=1.0e-04 wmin=7e-07 wmax=7.5e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.802364+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+  k1=0.88325
+  k2=-0.039841
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=101000.0
+  ua=-1.5041055e-10
+  ub=1.53437e-18
+  uc=5.7002e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.03919582
+  a0=0.80798
+  keta=-0.020254
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=1.46233e-7
+  b1=-3.2543e-11
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.10555+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.20557
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=2.8066e-5
+  alpha1=0.0
+  beta0=28.726
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.39073
+  kt2=-0.019151
+  at=60000.0
+  ute=-1.1327
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.73 nmos
* DC IV MOS Parameters
+  lmin=8e-06 lmax=2.0e-05 wmin=7e-07 wmax=7.5e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.801333355190753+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=2.04301948102928e-8
+  k1=0.88325
+  k2=-0.0410150615442501 lk2=2.32731061691134e-8
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=93894.3526750002 lvsat=0.140853335504342
+  ua=-1.50129029468138e-10 lua=-5.58050577409135e-18
+  ub=1.3931188576985e-18 lub=2.79998339728529e-24
+  uc=5.98416513530003e-11 luc=-5.62896449043049e-17
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0390626705994377 lu0=2.63938475016236e-9
+  a0=0.601793410698303 la0=4.08718129553509e-6
+  keta=-0.0192213995080001 lketa=-2.04689617833831e-8
+  a1=0.0
+  a2=0.65972622
+  ags=0.169673783278 lags=-1.86805120922095e-7
+  b0=2.20092618525e-07 lb0=-1.46409934978369e-12
+  b1=-5.375759457775e-11 lb1=4.20531201588797e-16
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.093150971365+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=2.45782609292891e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-0.3304370091775 lpclm=1.06251227570401e-5
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=2.62739427067501e-05 lalpha0=3.55234696606833e-11
+  alpha1=0.0
+  beta0=29.8733338800001 lbeta0=-2.27432908704254e-5
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.389426211500002 lkt1=-2.58446487163942e-8
+  kt2=-0.019151
+  at=1329.51750000007 lat=1.16300919223771
+  ute=-1.109231807 lute=-4.65203676895096e-7
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.74 nmos
* DC IV MOS Parameters
+  lmin=4e-06 lmax=8e-06 wmin=7e-07 wmax=7.5e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.805455934427748+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-1.18196335869371e-8
+  k1=0.88325
+  k2=-0.03631881536725 lk2=-1.34643643833373e-8
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=122316.941975 lvsat=-0.0814889349130361
+  ua=-1.51255111595588e-10 lua=3.22853179286087e-18
+  ub=1.9581234269045e-18 lub=-1.61989536138408e-24
+  uc=4.84830459410001e-11 luc=3.25656697689155e-17
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0395952682016876 lu0=-1.52698302348489e-9
+  a0=1.4265397679051 la0=-2.36458760012362e-6
+  keta=-0.023351801476 lketa=1.1842061734151e-8
+  a1=0.0
+  a2=0.65972622
+  ags=0.131978650166 lags=1.08073765422278e-7
+  b0=-7.53458555750002e-08 lb0=8.47036360151077e-13
+  b1=3.110078373325e-11 lb1=-2.43293065034391e-16
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.142747085905+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.42194453398709e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=1.8135910275325 lpclm=-6.14703183060035e-06 wpclm=-3.3881317890172e-21
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=3.34421718797501e-05 lalpha0=-2.05516589060489e-11
+  alpha1=0.0
+  beta0=25.2839983600001 lbeta0=1.31578463712788e-5
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.3946413655 lkt1=1.49520981491781e-8
+  kt2=-0.019151
+  at=236011.447500001 lat=-0.672844416713122
+  ute=-1.203104579 lute=2.69137766685274e-7
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.75 nmos
* DC IV MOS Parameters
+  lmin=2e-06 lmax=4e-06 wmin=7e-07 wmax=7.5e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.803064840069499+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-2.67912305971303e-9
+  k1=0.88325
+  k2=-0.0439011333024999 lk2=1.55207974395987e-8
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=91886.3450000002 lvsat=0.0348390514918053
+  ua=-1.50891494890295e-10 lua=1.83852294141966e-18
+  ub=1.3897700156735e-18 lub=5.5276684268443e-25
+  uc=5.7002e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.036635238377545 lu0=9.78841474618902e-9
+  a0=0.930704478229998 la0=-4.69142667388643e-7
+  keta=-0.020254
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=1.8879376885e-07 lb0=-1.62698370466729e-13
+  b1=-9.43563650375001e-11 lb1=2.36295866743168e-16 pb1=1.88079096131566e-37
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.173674571125+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-2.60421909901236e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.20557
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=2.8066e-5
+  alpha1=0.0
+  beta0=26.4494089809999 lbeta0=8.70279506265284e-6
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.407134578999999 lkt1=6.27102926852513e-8
+  kt2=-0.019151
+  at=96454.6199999999 lat=-0.13935620596722 wat=2.22044604925031e-16
+  ute=-1.099890842 lute=-1.25420585370503e-7
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.76 nmos
* DC IV MOS Parameters
+  lmin=1e-06 lmax=2e-06 wmin=7e-07 wmax=7.5e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.810756932415998+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-1.66997382345467e-8
+  k1=0.88325
+  k2=-0.0453829221079001 lk2=1.82216998306546e-8
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=114702.2895 lvsat=-0.00674827784262488
+  ua=-1.50579775480142e-10 lua=1.2703423092318e-18
+  ub=1.748272804802e-18 lub=-1.00687304646557e-25
+  uc=5.7002e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.04075821094055 lu0=2.27334484345046e-9
+  a0=0.30401250872 la0=6.73148212888284e-7
+  keta=-0.028147281214 lketa=1.43873283604754e-8
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=5.70307165400001e-08 lb0=7.74702296333292e-14
+  b1=-1.93830483417999e-10 lb1=4.17610426012975e-16 wb1=1.97215226305253e-31 pb1=1.88079096131566e-37
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.0408373182+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.82953310400041e-8
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-0.682345977130002 lpclm=1.61843197691014e-06 ppclm=1.21169035041947e-27
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=2.8066e-5
+  alpha1=0.0
+  beta0=27.720811402 lbeta0=6.3853704564211e-6
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.37273
+  kt2=-0.019151
+  at=16709.076 lat=0.00599846919344404
+  ute=-1.0618272431 lute=-1.94800287057094e-7
+  ua1=3.0044e-9
+  ub1=-3.9993193e-18 lub1=4.4988518950829e-25
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.81e-6
+  sbref=2.81e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.77 nmos
* DC IV MOS Parameters
+  lmin=8.0e-07 lmax=1e-06 wmin=7e-07 wmax=7.5e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.808054264405001+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-1.44761694791893e-8
+  k1=0.88325
+  k2=-0.0324074294452001 lk2=7.54635977677883e-9
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=113072.925705002 lvsat=-0.00540774973820035
+  ua=-1.458427290706e-10 lua=-2.62697262033675e-18
+  ub=1.46314648046001e-18 lub=1.33894961305667e-25
+  uc=4.75364888000007e-11 luc=7.78756949508693e-18
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0419916101619502 lu0=1.25858906862885e-9
+  a0=1.1222
+  keta=-0.0299111061340001 lketa=1.5838481800732e-8
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=5.194138403e-07 lb0=-3.0294670016086e-13
+  b1=1.2907003928e-09 lb1=-8.03759146308737e-16
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.795631165450011+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.83443372218159e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=1.8449465345 lpclm=-4.60849918475712e-7
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.48952393500001e-05 lalpha0=1.0835993080335e-11
+  alpha1=0.0
+  beta0=30.8800179100003 lbeta0=3.78619332688768e-6
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.378957310000004 lkt1=5.12340098360889e-9
+  kt2=-0.019151
+  at=8431.72500000009 lat=0.0128085024590251
+  ute=-1.45895323249999 lute=1.31927575327965e-7
+  ua1=6.09532531850002e-09 lua1=-2.54300007821482e-15
+  ub1=-8.5940785015e-18 lub1=4.23013602211759e-24
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.41e-6
+  sbref=2.41e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.78 nmos
* DC IV MOS Parameters
+  lmin=6e-07 lmax=8.0e-07 wmin=7e-07 wmax=7.5e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.795997689570001+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-6.96816657561652e-9
+  k1=0.88325
+  k2=-0.02240255567865 lk2=1.31601473126139e-9
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=95862.5157299992 lvsat=0.00530970607594128
+  ua=-1.54574698887e-10 lua=2.81069567540024e-18
+  ub=1.183899801145e-18 lub=3.07790525162176e-25
+  uc=4.9890115035e-11 luc=6.32189347613917e-18
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0408370924549 lu0=1.97754303485763e-9
+  a0=1.1222
+  keta=-0.0044772
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.934877494049992+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=9.67303667627495e-8
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=1.1049
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=5.960019529e-05 lalpha0=-1.7003168837137e-11
+  alpha1=0.0
+  beta0=37.7209158000003 lbeta0=-4.73845857049734e-7
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.37073
+  kt2=-0.019151
+  at=9131.64299999969 lat=0.012372641822967
+  ute=-1.13718993999999 lute=-6.84444015738594e-8
+  ua1=2.0117e-9
+  ub1=-1.8012e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.02e-6
+  sbref=2.01e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.79 nmos
* DC IV MOS Parameters
+  lmin=5e-07 lmax=6e-07 wmin=7e-07 wmax=7.5e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.898734058709998+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-5.03980146385351e-8
+  k1=0.88325
+  k2=-0.0234430747893 lk2=1.75587441542561e-9
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=103753.08243 lvsat=0.00197411892428345
+  ua=-1.55974388408999e-10 lua=3.40238782672487e-18
+  ub=1.21483649379999e-18 lub=2.94712626139433e-25
+  uc=1.51478909640001e-10 luc=-3.66228392560267e-17
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0423940107720999 lu0=1.3193853977094e-9
+  a0=1.1222
+  keta=0.015476612268 lketa=-8.43509501386391e-9
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.192100328+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.20056990557692e-8
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.524306931000012 lpclm=2.45434688651439e-7
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=3.52273194100001e-05 lalpha0=-6.69999864350872e-12
+  alpha1=0.0
+  beta0=35.4381684 lbeta0=4.91142234099748e-7
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.435276200000001 lkt1=2.72856796721994e-8
+  kt2=-0.019151
+  at=30344.63424 lat=0.00340525282309057
+  ute=-1.80352855299999 lute=2.13237586638246e-7
+  ua1=-1.19205063699998e-09 lua1=1.35432471052965e-15
+  ub1=-1.16186988900001e-18 lub1=-2.70264657153139e-25
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=1.81e-6
+  sbref=1.81e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.80 nmos
* DC IV MOS Parameters
+  lmin=2.0e-05 lmax=1.0e-04 wmin=4.2e-07 wmax=7.0e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.829863379957143+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} wvth0=-1.93141345141393e-8
+  k1=0.88325
+  k2=-0.0303668293285714 wk2=-6.65416482273651e-9
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=59217.7157142857 wvsat=0.0293457038035029
+  ua=-3.83702537663571e-10 wua=1.63852160951534e-16
+  ub=1.10028675914286e-18 wub=3.04877496049533e-25
+  uc=2.51494188714286e-11 wuc=2.23715966504899e-17
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.033313145882 wu0=4.13168440142906e-9
+  a0=0.361467660857143 wa0=3.13607048372307e-7
+  keta=-0.0283449809714286 wketa=5.68268430332091e-9
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=2.52240839614286e-07 wb0=-7.44543941374143e-14
+  b1=-2.47784296963e-08 wb1=1.73802240293729e-14
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.685826591142857+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} wnfactor=2.94791896763996e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-0.238498754285714 wpclm=3.11890801435063e-7
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.39535432571429e-05 walpha0=9.91185576843222e-12
+  alpha1=0.0
+  beta0=35.4503835142857 wbeta0=-4.72285731249154e-6
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.395255157142857 wkt1=3.17823506897152e-9
+  kt2=-0.019151
+  at=-241677.142857143 wat=0.211882337931429
+  ute=-1.27418658 wute=9.93728164898401e-8
+  ua1=3.0044e-9
+  ub1=-4.20531739142857e-18 wub1=3.18035389235074e-25
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.81 nmos
* DC IV MOS Parameters
+  lmin=8e-06 lmax=2.0e-05 wmin=4.2e-07 wmax=7.0e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.830040237339873+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-3.50579632321709e-09 wvth0=-2.01622212636721e-08 pvth0=1.6811395500651e-14
+  k1=0.88325
+  k2=-0.0350365507201248 lk2=9.25666309897083e-08 wk2=-4.19899512030268e-09 pk2=-4.8668168570696e-14
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=41394.0114735032 lvsat=0.353314494588591 wvsat=0.0368735096421888 pvsat=-1.49221670160502e-7
+  ua=-3.83472984958131e-10 lua=-4.55036153027141e-18 wua=1.63888660450486e-16 pua=-7.23519749355789e-25
+  ub=5.73305531446006e-19 lub=1.04462071186844e-23 wub=5.75794250066786e-25 pub=-5.3703099382772e-30
+  uc=3.22723597588459e-11 luc=-1.41196141140175e-16 wuc=1.93632368125709e-17 puc=5.96339078182704e-23
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0325932074479978 lu0=1.42711459137877e-08 wu0=4.5438145054874e-09 pu0=-8.16954418975049e-15
+  a0=-0.351465119514047 la0=1.41322747263802e-05 wa0=6.69519222177582e-07 pa0=-7.05515128096721e-12
+  keta=-0.0257548206487314 lketa=-5.13440513236997e-08 wketa=4.58873527135039e-09 pketa=2.16850573884619e-14
+  a1=0.0
+  a2=0.65972622
+  ags=0.18388848334906 lags=-4.68579296676391e-07 wags=-9.9836661655087e-09 pags=1.9790352879268e-13
+  b0=4.26221859352303e-07 lb0=-3.44877895337241e-12 wb0=-1.44774460036575e-13 pb0=1.39393575022133e-18
+  b1=-4.09112978563748e-08 lb1=3.19797505795628e-13 wb1=2.86962116877927e-14 pb1=-2.24313779352174e-19
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.478850580627578+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=4.10282977989755e-06 wnfactor=4.31452650833646e-07 pnfactor=-2.70898936617983e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-1.58301107886357 lpclm=2.66519061362915e-05 wpclm=8.7974289269587e-07 ppclm=-1.12563792528504e-11
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=-6.89600587874757e-06 lalpha0=4.13295003992038e-10 walpha0=2.32968470491271e-11 palpha0=-2.65327081594559e-16
+  alpha1=0.0
+  beta0=39.3224637900319 lbeta0=-7.67552057165222e-05 wbeta0=-6.63657749405106e-06 pbeta0=3.79351603683258e-11
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.406734372303882 lkt1=2.27549394228119e-07 wkt1=1.2156352124285e-08 pkt1=-1.77970799273993e-13
+  kt2=-0.019151
+  at=-455710.285237293 lat=4.24272140648641 wat=0.321000991372932 pat=-2.16302971425315e-6
+  ute=-1.29191899110746 lute=3.51504815364543e-07 wute=1.28309978383505e-07 pute=-5.73613576121564e-13
+  ua1=3.0044e-9
+  ub1=-4.50050644520086e-18 lub1=5.85145320707254e-24 wub1=5.25360830773931e-25 pub1=-4.10975645708097e-30
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.82 nmos
* DC IV MOS Parameters
+  lmin=4e-06 lmax=8e-06 wmin=4.2e-07 wmax=7.0e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.825094685478934+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=3.51819255314485e-08 wvth0=-1.37932375232973e-08 pvth0=-3.30114510436738e-14
+  k1=0.88325
+  k2=-0.0136677548587363 lk2=-7.45957108278474e-08 wk2=-1.59089270460336e-08 pk2=4.2935478912609e-14
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=104039.599191698 lvsat=-0.136745086467747 wvsat=0.012837055149167 pvsat=3.88090475321497e-8
+  ua=-3.8312220969584e-10 lua=-7.29438204862381e-18 wua=1.62851392616516e-16 pua=7.39074749073964e-24
+  ub=2.49460890589185e-18 lub=-4.58363234899766e-24 wub=-3.76799503195806e-25 pub=2.08157474577644e-30
+  uc=-3.1699983691757e-11 luc=3.59242293113505e-16 wuc=5.63163904965077e-17 puc=-2.29440673052826e-22
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0349806758861491 lu0=-4.40537744886079e-09 wu0=3.24104968363374e-09 pu0=2.02163456787375e-15
+  a0=2.2133134063879 la0=-5.93129775632726e-06 wa0=-5.52588891441116e-07 pa0=2.5050717447893e-12
+  keta=-0.0444619681608831 lketa=9.49969314411826e-08 wketa=1.48266833507943e-08 pketa=-5.84036564289943e-14
+  a1=0.0
+  a2=0.65972622
+  ags=0.0893345499528206 lags=2.71090689274304e-07 wags=2.99509984965261e-08 pags=-1.14494610433624e-13
+  b0=-2.97254339359509e-07 lb0=2.21078073405265e-12 wb0=1.55856979769082e-13 pb0=-9.5782313352102e-19
+  b1=2.46170943585901e-09 lb1=-1.94978629125554e-14 wb1=-1.70713312560322e-15 pb1=1.35234086232667e-20
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.840734150971558+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.27191195577701e-06 wnfactor=2.12118180824633e-07 pnfactor=-9.9319480827175e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=3.79503821944784 lpclm=-1.54191268291375e-05 wpclm=-1.39166547234736e-06 ppclm=6.51223737803255e-12
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=4.36625087600007e-05 lalpha0=1.77893442135483e-11 walpha0=-7.17823316717034e-12 palpha0=-2.69287268590427e-17
+  alpha1=0.0
+  beta0=26.8094775473051 lbeta0=2.11305196670302e-05 wbeta0=-1.07141725624535e-06 pbeta0=-5.59959114392443e-12
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.365142126282251 lkt1=-9.7815558084927e-08 wkt1=-2.07187316661081e-08 pkt1=7.92021378207134e-14
+  kt2=-0.019151
+  at=140945.406935236 lat=-0.424755572998083 wat=0.0667694434585811 pat=-1.7424470320557e-7
+  ute=-1.35620563054012 lute=8.54401902540276e-07 wute=1.07530217347102e-07 pute=-4.11059095289506e-13
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.83 nmos
* DC IV MOS Parameters
+  lmin=2e-06 lmax=4e-06 wmin=4.2e-07 wmax=7.0e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.828706914689571+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=2.13733449488423e-08 wvth0=-1.80096598252579e-08 pvth0=-1.68932028008778e-14
+  k1=0.88325
+  k2=-0.039432867350833 lk2=2.38973834141779e-08 wk2=-3.13827765462142e-09 pk2=-5.88327840607348e-15
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=42658.0865916858 lvsat=0.0978999245752087 wvsat=0.0345753688365627 pvsat=-4.42906780883824e-8
+  ua=-4.95338611218774e-10 lua=4.21678734761542e-16 wua=2.41921743259075e-16 pua=-2.94873933091439e-22
+  ub=9.80320658020081e-19 lub=1.20508427907743e-24 wub=2.87575937449164e-25 pub=-4.5815384681575e-31
+  uc=7.23050598093979e-11 luc=-3.83410108347095e-17 wuc=-1.0748073451011e-17 puc=2.69287322777365e-23
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0323195500644227 lu0=5.76739072475335e-09 wu0=3.0311150553448e-09 pu0=2.82415817940729e-15
+  a0=0.836277238788978 la0=-6.67258910325673e-07 wa0=6.63207827669228e-08 pa0=1.39146546994335e-13
+  keta=-0.0196114276857143 wketa=-4.51309379793941e-10
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=4.2676755444091e-07 lb0=-5.56960204056926e-13 wb0=-1.67140412362205e-13 pb0=2.76909010298408e-19
+  b1=8.83699715181148e-09 lb1=-4.38688728982461e-14 wb1=-6.27291827985186e-15 pb1=3.09771770717527e-20
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.26557044870923+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-3.52122929510027e-07 wnfactor=-6.45428858295311e-08 pnfactor=6.44060277201906e-14
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-0.238498754285714 wpclm=3.11890801435063e-7
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=5.00660594762677e-05 lalpha0=-6.68970761959775e-12 walpha0=-1.54516977730377e-11 palpha0=4.69850276720925e-18
+  alpha1=0.0
+  beta0=31.5630213168573 lbeta0=2.95900053930625e-06 wbeta0=-3.59153539686469e-06 pbeta0=4.03414259588348e-12
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.407134579 lkt1=6.27102926852491e-8
+  kt2=-0.019151
+  at=38793.0917004286 lat=-0.0342547508282139 wat=0.0404984590781474 pat=-7.38177968139707e-8
+  ute=-1.099890842 lute=-1.25420585370499e-7
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.84 nmos
* DC IV MOS Parameters
+  lmin=1e-06 lmax=2e-06 wmin=4.2e-07 wmax=7.0e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.82550588050513+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=2.72079691888823e-08 wvth0=-1.03588941925044e-08 pvth0=-3.08384904934318e-14
+  k1=0.88325
+  k2=-0.0337785900796947 lk2=1.35911569494788e-08 wk2=-8.15027939134591e-09 pk2=3.25225253150811e-15
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=109440.465509034 lvsat=-0.0238263877311877 wvsat=0.00369563155640729 pvsat=1.19947763240126e-8
+  ua=-2.61621187577944e-10 lua=-4.32525854873159e-18 wua=7.79897137040678e-17 pua=3.93005907138902e-24
+  ub=1.64503250918819e-18 lub=-6.50661811407619e-27 wub=7.25106151437669e-26 pub=-6.61476168247137e-32
+  uc=5.12701342857143e-11 wuc=4.02576442069713e-18
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0342049949863969 lu0=2.33073181667854e-09 wu0=4.60263811896757e-09 pu0=-4.03056258728715e-17
+  a0=-0.0662191907906005 la0=9.77749309258342e-07 wa0=2.60031493687871e-07 pa0=-2.13935970833316e-13
+  keta=-0.0269760447370097 lketa=1.34237158025247e-08 wketa=-8.22615597141188e-10 pketa=6.7679135285157e-16
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=1.52785413629952e-07 lb0=-5.75644625544266e-14 wb0=-6.72531199917333e-14 pb0=9.4841345988686e-20
+  b1=-2.4398393366071e-08 lb1=1.67103036958044e-14 wb1=1.70000263315056e-14 pb1=-1.14431405326515e-20
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.949326724901382+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=2.24304309429983e-07 wnfactor=6.42722821820981e-08 pnfactor=-1.70389372284815e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-1.6760517212323 lpclm=2.62027235699552e-06 wpclm=6.97927241958765e-07 ppclm=-7.03640587272208e-13
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=4.46001824407663e-05 lalpha0=3.2731158951988e-12 walpha0=-1.16127499689073e-11 palpha0=-2.29886640276109e-18
+  alpha1=0.0
+  beta0=27.6281323584481 lbeta0=1.01312446253563e-05 wbeta0=6.50929408805778e-08 pbeta0=-2.63090723080329e-12
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.37273
+  kt2=-0.019151
+  at=16709.076 lat=0.00599846919344402
+  ute=-1.0618272431 lute=-1.94800287057094e-7
+  ua1=3.0044e-9
+  ub1=-4.37161800613e-18 lub1=1.12848558243134e-24 wub1=2.61483251652993e-25 pub1=-4.76613628768712e-31
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.81e-6
+  sbref=2.81e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.85 nmos
* DC IV MOS Parameters
+  lmin=8.0e-07 lmax=1e-06 wmin=4.2e-07 wmax=7.0e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.9502414186827+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-7.54158248714876e-08 wvth0=-9.98648634326337e-08 pvth0=4.2800845085469e-14
+  k1=0.88325
+  k2=-0.036633482656502 lk2=1.5939965574088e-08 wk2=2.96816002085153e-09 pk2=-5.8952322445285e-15
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=47296.6147484926 lvsat=0.0273012847488832 wvsat=0.0461978604476812 pvsat=-2.29731249539341e-8
+  ua=-3.88716722579163e-10 lua=1.00240178058357e-16 wua=1.70582063592752e-16 pua=-7.22485375448784e-23
+  ub=3.03979129562241e-19 lub=1.09681956995896e-24 wub=8.14138870568339e-25 pub=-6.76308173038426e-31
+  uc=-1.24504160297532e-11 luc=5.24248720815948e-17 wuc=4.21316826333675e-17 puc=-3.13509201970285e-23
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0402734029207484 lu0=-2.66193551155848e-09 wu0=1.20677941944345e-09 pu0=2.75357259784529e-15
+  a0=1.1222
+  keta=-0.0589491996107237 lketa=3.97290214849303e-08 wketa=2.03948468771899e-08 pketa=-1.67794727661174e-14
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=2.38142167818785e-07 lb0=-1.2779011028496e-13 wb0=1.97550596623836e-13 pb0=-1.23020880586158e-19
+  b1=-1.68150543832829e-08 lb1=1.04712556311561e-14 wb1=1.27165406554723e-14 pb1=-7.91898407892289e-21
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.01618125680964+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.69301013538566e-07 wnfactor=-1.54902915566264e-07 pnfactor=9.93285733389253e-15
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=2.91385884361788 lpclm=-1.15598935193423e-06 wpclm=-7.50748422484323e-07 ppclm=4.88229790810718e-13
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=-6.20121687575445e-06 lalpha0=4.50690019562792e-11 walpha0=1.48170538372462e-11 palpha0=-2.40434853180016e-17
+  alpha1=0.0
+  beta0=28.3987504251882 lbeta0=9.49723325268927e-06 wbeta0=1.74271325542266e-06 pbeta0=-4.01113746980679e-12
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.37895731 lkt1=5.12340098360974e-9
+  kt2=-0.019151
+  at=8431.72500000001 lat=0.012808502459025
+  ute=-1.4589532325 lute=1.31927575327958e-7
+  ua1=6.0953253185e-09 lua1=-2.54300007821482e-15
+  ub1=-6.73258497085e-18 lub1=3.07092629428239e-24 wub1=-1.30741625826497e-24 pub1=8.14168633925601e-31
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.41e-6
+  sbref=2.41e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.86 nmos
* DC IV MOS Parameters
+  lmin=6e-07 lmax=8.0e-07 wmin=4.2e-07 wmax=7.0e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.813398532560909+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=9.80048244602145e-09 wvth0=-1.22214472729793e-08 pvth0=-1.17774271030487e-14
+  k1=0.88325
+  k2=0.00276616484055717 lk2=-8.59541631140312e-09 wk2=-1.76772005192241e-08 pk2=6.96127376995335e-15
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=63054.8854495002 lvsat=0.0174881210769738 wvsat=0.0230423735122485 pvsat=-8.55348541914514e-9
+  ua=-2.40767086464583e-10 lua=8.10735321108734e-18 wua=6.05370510303399e-17 pua=-3.72009682687469e-24
+  ub=1.93648646732793e-18 lub=8.02066430047961e-26 wub=-5.28577739820248e-25 pub=1.59843084465469e-31
+  uc=4.6270162837865e-11 luc=1.58577472827842e-17 wuc=2.54246618575341e-18 puc=-6.69748784938932e-24
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0320679037535301 lu0=2.44788319034262e-09 wu0=6.1590221460298e-09 pu0=-3.30342467524536e-16
+  a0=1.1222
+  keta=0.00484884719428572 wketa=-6.55013059481218e-9
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.966101666153628+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=2.00487127107379e-07 wnfactor=-2.19302348286379e-08 pnfactor=-7.28733531145297e-14
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=2.43420447416318 lpclm=-8.5729370678934e-07 wpclm=-9.33634338819565e-07 ppclm=6.0211852037608e-13
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=0.000134661383131218 lalpha0=-4.26505058086625e-11 walpha0=-5.27190751579035e-11 palpha0=1.8013355827277e-17
+  alpha1=0.0
+  beta0=49.7062182813655 lbeta0=-3.77158751285595e-06 wbeta0=-8.41785322718211e-06 pbeta0=2.31616225647214e-12
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.37073
+  kt2=-0.019151
+  at=9131.64299999998 lat=0.012372641822967
+  ute=-1.13718994 lute=-6.84444015738602e-8
+  ua1=2.0117e-9
+  ub1=-1.8012e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.02e-6
+  sbref=2.01e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.87 nmos
* DC IV MOS Parameters
+  lmin=5e-07 lmax=6e-07 wmin=4.2e-07 wmax=7.0e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=8.86345e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.174e-9
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.11128e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.11128e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.913698747061291+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-3.25995275299398e-08 wvth0=-1.05104189341533e-08 pvth0=-1.25007318237489e-14
+  k1=0.88325
+  k2=0.00860863579909676 lk2=-1.10652099021775e-08 wk2=-2.25114548283393e-08 pk2=9.0048629282999e-15
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=117634.619845754 lvsat=-0.00558442462408915 wvsat=-0.00974967004088034 pvsat=5.30872794411253e-9
+  ua=-4.91558500800461e-10 lua=1.14124658584708e-16 wua=2.35696830169918e-16 pua=-7.77655654223276e-23
+  ub=7.04880950984635e-20 lub=8.69022000895732e-25 wub=8.03730809131227e-25 pub=-4.03365040741338e-31
+  uc=2.31534787583976e-10 luc=-6.24593528007643e-17 wuc=-5.62270857621959e-17 puc=1.81462236151193e-23
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0242708432803261 lu0=5.74394236124058e-09 wu0=1.27287704415124e-08 pu0=-3.1075787342222e-15
+  a0=1.1222
+  keta=0.0549007048328759 lketa=-2.11584718314189e-08 wketa=-2.76894325647555e-08 pketa=8.93623826105611e-15
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={2.12439448710056+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-2.89159155384341e-07 wnfactor=-6.54794938055964e-07 pnfactor=1.94658175745461e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-0.302893278965829 lpclm=2.99762363488641e-07 wpclm=5.8098241306908e-07 ppclm=-3.8156933766559e-14
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=9.60608596678027e-05 lalpha0=-2.63328679244496e-11 walpha0=-4.27263153329872e-11 palpha0=1.37891064737303e-17
+  alpha1=0.0
+  beta0=53.1263408744397 lbeta0=-5.21737935674879e-06 wbeta0=-1.24232525610778e-05 pbeta0=4.0093687222892e-12
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.362255775506429 lkt1=-3.58231739439185e-09 wkt1=-5.1285749102211e-08 pkt1=2.16800760037267e-14
+  kt2=-0.019151
+  at=72715.9525594697 lat=-0.0145064169414172 wat=-0.0297594106790429 pat=1.25802254357625e-8
+  ute=-2.56196736207323 lute=5.33853182836577e-07 wute=5.32687980674964e-07 pute=-2.25183722758708e-13
+  ua1=-1.192050637e-09 lua1=1.35432471052965e-15
+  ub1=-9.69649710380863e-18 lub1=3.33758683999013e-24 wub1=5.99427835506641e-24 pub1=-2.53396728331558e-30
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.461036368e-10
+  cgso=2.461036368e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=4.0116e-11
+  cgdl=4.0116e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=7.81225e-8
+  dwc=-2.252e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000741207936
+  mjs=0.295
+  pbs=0.72468
+  cjsws=7.232371132e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.583682e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=1.81e-6
+  sbref=1.81e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.ends sky130_fd_pr__nfet_g5v0d10v5
