* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 68
.param
+  sky130_fd_pr__pfet_01v8_hvt__toxe_mult=0.948
+  sky130_fd_pr__pfet_01v8_hvt__rshp_mult=1.0
+  sky130_fd_pr__pfet_01v8_hvt__overlap_mult=0.91064
+  sky130_fd_pr__pfet_01v8_hvt__lint_diff=1.7325e-8
+  sky130_fd_pr__pfet_01v8_hvt__wint_diff=-3.2175e-8
+  sky130_fd_pr__pfet_01v8_hvt__dlc_diff=1.7325e-8
+  sky130_fd_pr__pfet_01v8_hvt__dwc_diff=-3.2175e-8
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 000, W = 1.26, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_0=1.6702
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_0=-0.098011
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_0=0.00097522
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_0=6.9012e-20
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_0=0.00086508
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_0=-29674.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_0=-0.030352
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_0=1.8215e-10
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_0=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 001, W = 1.68, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_1=1.7209
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_1=-0.12703
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_1=-2.6856e-20
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_1=-0.0068783
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_1=0.00054806
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_1=-23641.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_1=-0.059296
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_1=1.9021e-10
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_1=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 002, W = 1.0, L = 1.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_2=0.88917
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_2=-0.16742
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_2=0.22697
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_2=-0.05321
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_2=1.7862e-19
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_2=-0.0030523
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_2=0.0021726
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_2=0.02652
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_2=2.0425e-10
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 003, W = 1.0, L = 2.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_3=-5.5786e-11
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_3=0.56532
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_3=-0.11759
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_3=0.1273
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_3=-0.04025
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_3=5.1865e-19
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_3=-0.0062951
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_3=0.0020197
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_3=0.036899
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_3=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 004, W = 1.0, L = 4.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_4=-6.1212e-11
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_4=0.3705
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_4=-0.085417
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_4=0.18515
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_4=-0.063572
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_4=4.5105e-19
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_4=-0.0087946
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_4=0.0016238
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_4=0.029425
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_4=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 005, W = 1.0, L = 8.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_5=3.4914e-11
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_5=0.58901
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_5=-0.052472
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_5=0.051784
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_5=-0.063375
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_5=4.024e-19
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_5=-0.010302
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_5=0.0021038
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_5=0.025149
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_5=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 006, W = 1.0, L = 0.15
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_6=4.112e-10
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_6=2.3478
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_6=-0.15288
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_6=-1.3862e-19
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_6=-0.013041
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_6=0.0015364
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_6=-27670.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_6=-0.053351
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 007, W = 1.0, L = 0.18
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_7=0.0010756
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_7=3.3792e-19
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_7=-15990.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_7=-0.059438
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_7=1.0152e-10
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_7=1.0669
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_7=-0.11315
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_7=0.013182
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 008, W = 1.0, L = 0.25
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_8=0.0065099
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_8=0.0021339
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_8=3.4578e-19
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_8=-29944.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_8=0.037342
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_8=4.1649e-10
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_8=1.2977
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_8=-0.045339
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 009, W = 1.0, L = 0.5
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_9=-0.073336
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_9=-0.012277
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_9=0.0045307
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_9=4.1908e-20
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_9=-10537.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_9=0.045267
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_9=7.7724e-10
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_9=1.4783
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 010, W = 3.0, L = 1.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_10=7.2706e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_10=-0.071099
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_10=-0.0037068
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_10=0.00973
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_10=0.2504
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_10=0.0023319
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_10=0.020152
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_10=-0.010112
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_10=-1.437e-10
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 011, W = 3.0, L = 2.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_11=-1.3981e-10
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_11=9.452e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_11=-0.10271
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_11=0.025822
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_11=-0.010134
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_11=-0.17771
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_11=0.0035013
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_11=0.013621
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_11=-0.011751
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 012, W = 3.0, L = 4.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_12=-0.010705
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_12=-1.7178e-10
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_12=1.079e-18
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_12=-0.067375
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_12=0.067597
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_12=-0.042239
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_12=0.27193
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_12=0.0041731
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_12=-0.017373
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 013, W = 3.0, L = 8.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_13=0.27144
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_13=0.0048327
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_13=0.00227
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_13=-0.00843
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_13=-3.3818e-10
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_13=1.4661e-18
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_13=-0.066337
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_13=0.037844
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_13=-0.021169
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_13=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 014, W = 3.0, L = 0.15
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_14=-24444.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_14=1.2545
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_14=0.00041791
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_14=-0.049892
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_14=-0.0042041
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_14=9.4745e-11
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_14=4.124e-20
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_14=-0.12375
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_14=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 015, W = 3.0, L = 0.18
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_15=-6505.6
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_15=0.66146
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_15=0.00089379
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_15=-0.071254
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_15=-8.1586e-5
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_15=1.6305e-10
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_15=1.0152e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_15=-0.093754
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_15=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 016, W = 3.0, L = 0.25
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_16=-28762.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_16=0.70713
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_16=0.0012256
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_16=-0.001682
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_16=0.0028259
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_16=1.3012e-10
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_16=2.539e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_16=-0.04469
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_16=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 017, W = 3.0, L = 0.5
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_17=0.52823
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_17=0.0026198
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_17=13859.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_17=0.016554
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_17=-0.006883
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_17=1.1056e-10
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_17=5.0826e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_17=-0.073286
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_17=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 018, W = 5.0, L = 1.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_18=-0.008952
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_18=0.011728
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_18=0.28249
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_18=0.0023179
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_18=0.016121
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_18=-0.011899
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_18=-1.6357e-10
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_18=7.6564e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_18=-0.06502
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 019, W = 5.0, L = 2.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_19=-0.077046
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_19=0.038942
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_19=-0.039498
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_19=0.12738
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_19=0.0031187
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_19=0.0029058
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_19=-0.0081995
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_19=-2.5441e-10
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_19=1.0061e-18
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_19=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 020, W = 5.0, L = 4.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_20=-0.066055
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_20=0.016281
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_20=-0.015815
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_20=0.26745
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_20=0.0046376
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_20=0.0014783
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_20=-0.0077373
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_20=-3.3629e-10
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_20=1.4023e-18
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 021, W = 5.0, L = 8.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_21=1.3543e-18
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_21=-0.04378
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_21=-0.038207
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_21=-0.044188
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_21=0.36554
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_21=0.0039903
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_21=0.01708
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_21=-0.0066951
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_21=-4.1477e-10
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 022, W = 5.0, L = 0.15
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_22=1.324e-10
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_22=-4.5976e-20
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_22=-0.084594
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_22=-26795.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_22=1.0827
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_22=0.00042769
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_22=-0.071575
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_22=0.00045233
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 023, W = 5.0, L = 0.18
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_23=0.0076182
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_23=1.5074e-10
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_23=7.5942e-20
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_23=-0.048212
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_23=-20619.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_23=0.71624
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_23=0.00066193
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_23=-0.050276
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 024, W = 5.0, L = 0.25
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_24=0.31532
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_24=0.00084832
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_24=-0.0077162
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_24=0.001811
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_24=-2.852e-13
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_24=3.5019e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_24=-0.050657
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_24=-11016.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 025, W = 5.0, L = 0.5
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_25=-2879.9
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_25=0.28888
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_25=0.00033371
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_25=0.028527
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_25=-0.0086212
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_25=-1.3033e-11
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_25=1.7081e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_25=-0.056202
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_25=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 026, W = 7.0, L = 1.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_26=0.11511
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_26=0.0033142
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_26=0.0065868
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_26=-0.0096254
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_26=-2.915e-10
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_26=1.086e-18
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_26=-0.066547
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_26=0.017504
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_26=-0.021718
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_26=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 027, W = 7.0, L = 2.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_27=-0.025453
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_27=0.004512
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_27=0.0029878
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_27=-0.010442
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_27=-3.7793e-10
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_27=1.4138e-18
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_27=-0.058137
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_27=0.045741
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_27=-0.048361
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_27=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 028, W = 7.0, L = 4.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_28=0.36762
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_28=0.0049774
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_28=0.017746
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_28=-0.0066393
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_28=-4.132e-10
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_28=1.5608e-18
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_28=-0.045427
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_28=-0.0082778
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_28=0.0056012
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 029, W = 7.0, L = 8.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_29=-0.00067009
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_29=0.0017417
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_29=0.97578
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_29=0.0092277
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_29=0.008761
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_29=-0.011014
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_29=-5.3257e-11
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_29=1.8573e-18
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_29=-0.034623
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 030, W = 7.0, L = 0.15
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_30=-0.088188
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_30=-18897.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_30=1.1748
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_30=0.00083903
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_30=-0.073728
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_30=-0.019298
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_30=2.86e-10
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_30=-1.7396e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_30=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 031, W = 7.0, L = 0.18
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_31=-0.086699
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_31=-4248.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_31=0.42507
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_31=0.00024638
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_31=-0.085301
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_31=0.0015551
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_31=-1.6895e-11
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_31=1.885e-19
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 032, W = 7.0, L = 0.25
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_32=2.5238e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_32=-0.06692
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_32=-11755.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_32=0.35759
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_32=0.00068645
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_32=-0.0035656
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_32=8.2421e-5
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_32=2.8428e-11
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 033, W = 7.0, L = 0.5
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_33=1.9174e-10
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_33=1.8e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_33=-0.047344
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_33=-32711.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_33=0.97073
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_33=0.0021523
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_33=0.013441
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_33=-0.0091659
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 034, W = 0.42, L = 1.0
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_34=-0.011769
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_34=-1.0721e-10
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_34=1.3365e-18
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_34=-0.12761
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_34=7.2095e-8
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_34=5.0779e-8
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_34=1.0947
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_34=0.0050028
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_34=0.046227
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 035, W = 0.42, L = 20.0
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_35=0.49911
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_35=0.003451
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_35=-0.0087503
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_35=-0.017093
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_35=-1.9758e-10
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_35=9.821e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_35=-0.094876
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_35=-1.0283e-7
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_35=2.3178e-9
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_35=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 036, W = 0.42, L = 2.0
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_36=0.69604
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_36=0.0062132
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_36=0.013867
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_36=-0.018297
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_36=6.1158e-11
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_36=1.2575e-18
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_36=-0.099857
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_36=5.6678e-8
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_36=1.5052e-8
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 037, W = 0.42, L = 4.0
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_37=-1.0273e-9
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_37=0.74962
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_37=0.0031442
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_37=0.033856
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_37=-0.012048
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_37=1.0374e-10
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_37=4.574e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_37=-0.076379
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_37=9.5235e-8
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_37=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 038, W = 0.42, L = 8.0
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_38=1.91e-8
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_38=-2.6206e-7
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_38=0.5372
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_38=0.0060424
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_38=0.0034632
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_38=-0.016469
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_38=7.736e-10
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_38=3.488e-20
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_38=-0.087212
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_38=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 039, W = 0.42, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_39=2.2787
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_39=0.0025449
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_39=-50000.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_39=0.040102
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_39=-0.0018016
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_39=5.933e-10
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_39=2.2929e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_39=-0.19968
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_39=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 040, W = 0.42, L = 0.18
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_40=-45149.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_40=1.9521
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_40=0.0021813
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_40=0.00501
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_40=-0.0085993
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_40=5.5697e-10
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_40=6.3421e-20
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_40=-0.19674
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_40=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 041, W = 0.42, L = 0.5
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_41=-0.093014
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_41=-38889.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_41=1.6445
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_41=0.0057123
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_41=0.091479
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_41=-0.023719
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_41=4.3063e-10
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_41=8.5174e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_41=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 042, W = 0.55, L = 1.0
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_42=-0.08843
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_42=1.0665e-7
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_42=9.4459e-9
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_42=1.3174
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_42=0.0047
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_42=0.034666
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_42=-0.014806
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_42=7.2762e-10
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_42=-4.3961e-20
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 043, W = 0.55, L = 2.0
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_43=2.8498e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_43=-0.061848
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_43=1.1443e-7
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_43=-1.6295e-9
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_43=0.73413
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_43=0.003296
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_43=0.041686
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_43=-0.0061916
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_43=2.8632e-10
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 044, W = 0.55, L = 4.0
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_44=-4.6452e-11
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_44=5.5996e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_44=-0.069356
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_44=9.4887e-8
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_44=2.3137e-9
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_44=0.4916
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_44=0.0024626
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_44=0.03279
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_44=-0.0078584
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 045, W = 0.55, L = 8.0
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_45=-0.0088326
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_45=-1.474e-10
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_45=5.7719e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_45=-0.067651
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_45=7.7369e-8
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_45=7.0231e-10
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_45=0.3621
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_45=0.0019517
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_45=0.026283
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 046, W = 0.55, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_46=2.0889
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_46=0.0012322
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_46=-0.039462
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_46=-0.016442
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_46=2.1814e-10
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_46=1.5922e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_46=-0.13831
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_46=-40582.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 047, W = 0.55, L = 0.5
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_47=-50000.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_47=3.6882
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_47=0.015631
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_47=0.074708
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_47=-0.0080946
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_47=2.0e-9
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_47=1.1367e-18
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_47=-0.075714
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_47=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 048, W = 0.64, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_48=-24472.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_48=2.5262
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_48=0.0012175
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_48=-0.023234
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_48=-0.007354
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_48=2.5998e-10
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_48=1.7343e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_48=-0.19561
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_48=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 049, W = 0.84, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_49=-30755.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_49=1.8113
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_49=0.001795
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_49=-0.012419
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_49=-0.0068842
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_49=5.2165e-10
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_49=-1.2533e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_49=-0.15886
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_49=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 050, W = 0.64, L = 0.18
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_50=-29893.59829279
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_50=0.00124944
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_50=1.72013046
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_50=-0.04127798
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_50=0.0010617
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_50=3.46701e-10
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_50=1.396e-20
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_50=-0.103349
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_50=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 051, W = 2.0, L = 0.15
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_51=-14190.02188706
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_51=3.06099e-5
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_51=0.96707997
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_51=-0.07541995
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_51=0.00703588
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_51=5.6917e-11
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_51=-2.9419e-20
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_51=-0.082426
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_51=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 052, W = 1.12, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_52=-0.072042
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_52=-7.6647e-8
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_52=-26609.98832683
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_52=0.0003282
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_52=1.21669943
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_52=-0.05314867
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_52=0.012422
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_52=6.42999e-11
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_52=1.03621e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_52=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 053, W = 1.65, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_53=-0.09478604
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_53=-16214.19463122
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_53=-0.00051934
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_53=1.11233043
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_53=-0.071217
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_53=0.00941368
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_53=-1.5565e-10
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_53=2.02164e-19
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 054, W = 0.84, L = 0.18
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_54=-2.0137e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_54=-0.109857
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_54=-24608.56214497
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_54=0.00160218
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_54=0.39679982
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_54=-0.06057999
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_54=0.00330583
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_54=5.29585e-10
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 055, W = 1.68, L = 0.18
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_55=1.77615e-10
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_55=-1.065e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_55=-0.036074
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_55=-39429.59956441
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_55=0.00036125
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_55=0.53532009
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_55=-0.0623438
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_55=0.01331141
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 056, W = 0.36, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_56=-0.0066348
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_56=-30180.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_56=-0.001025
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_56=0.08346
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 057, W = 0.54, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_57=-0.00056441
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_57=0.0086191
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_57=0.0054426
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_57=-37723.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_57=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 058, W = 0.63, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_58=-30636.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_58=-0.00052667
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_58=-0.00043348
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_58=0.0051619
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_58=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 059, W = 0.7, L = 0.15
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_59=-27201.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_59=0.00143932
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_59=0.0013145
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_59=1.243108
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_59=-0.044733
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_59=-0.005647
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_59=4.11678e-10
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_59=-6.27298e-20
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_59=-0.00026826
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_59=-0.00136297
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_59=-0.10590279
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_59=4.2886e-12
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_59=-7.09239e-5
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_59=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 060, W = 0.75, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_60=-7.29796e-5
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_60=-25393.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_60=0.0012886
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_60=0.00148104
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_60=0.90432662
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_60=-0.05008
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_60=-0.0047585
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_60=4.5847e-10
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_60=-1.17829e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_60=-0.00027604
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_60=-0.10757491
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_60=-0.00140248
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_60=4.41291e-12
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 061, W = 0.79, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_61=3.018e-12
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_61=-4.9911e-5
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_61=-23783.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_61=0.00101288
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_61=0.0013326
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_61=0.66438835
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_61=-0.052569
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_61=-0.0044981
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_61=4.91938e-10
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_61=-1.57174e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_61=-0.00018878
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_61=-0.10868729
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_61=-0.00095916
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_61=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 062, W = 0.82, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_62=1.34608e-12
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_62=-2.22611e-5
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_62=-21900.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_62=0.00045176
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_62=0.0013726
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_62=0.49989482
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_62=-0.054622
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_62=-0.0029267
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_62=5.1504e-10
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_62=-1.84303e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_62=-8.42008e-5
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_62=-0.10941523
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_62=-0.0004278
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 063, W = 0.82, L = 0.18
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_63=-0.0004278
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_63=-0.10941523
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_63=1.34608e-12
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_63=-2.22613e-5
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_63=-23535.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_63=0.00045176
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_63=0.0015171
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_63=0.49989469
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_63=-0.034774
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_63=-0.013873
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_63=5.1504e-10
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_63=-1.84303e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_63=-8.42007e-5
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_63=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 064, W = 0.82, L = 0.25
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_64=-0.0001157
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_64=-434810.89830208
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_64=-0.00046359
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_64=0.00047433
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_64=-0.0245589
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_64=1.562e-12
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_64=3.46622e-5
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_64=-19223.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_64=0.0022188
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_64=0.81033175
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_64=0.019208
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_64=0.0049685
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_64=2.61701e-10
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_64=3.89042e-19
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 065, W = 0.82, L = 0.5
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_65=-15187.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_65=-0.00058999
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_65=0.046929
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_65=-0.0016053
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_65=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 066, W = 0.86, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_66=4.61965e-10
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_66=-1.56897e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_66=0.00031999
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_66=-0.10432908
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_66=-4.53896e-13
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_66=1.91787e-6
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_66=-18965.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_66=2.59995e-5
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_66=0.0012435
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_66=0.51671158
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_66=-0.056768
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_66=-0.0024326
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 067, W = 0.94, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_67=-0.0012624
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_67=2.20238e-10
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_67=1.67256e-21
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_67=7.9727e-5
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_67=0.00057533
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_67=-0.08465745
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_67=-8.16075e-13
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_67=3.44709e-6
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_67=-17711.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_67=4.67463e-5
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_67=0.00053342
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_67=0.94327401
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_67=-0.047237
.include "sky130_fd_pr__pfet_01v8_hvt__fs.pm3.spice"
