* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 18
.param
+  sky130_fd_pr__rf_nfet_01v8_lvt_b__toxe_mult=1.0365
+  sky130_fd_pr__rf_nfet_01v8_lvt_b__rbpb_mult=1.2
+  sky130_fd_pr__rf_nfet_01v8_lvt_b__overlap_mult=9.6320e-1
+  sky130_fd_pr__rf_nfet_01v8_lvt_b__ajunction_mult=1.1229e+0
+  sky130_fd_pr__rf_nfet_01v8_lvt_b__pjunction_mult=1.0009e+0
+  sky130_fd_pr__rf_nfet_01v8_lvt_b__lint_diff=-1.21275e-8
+  sky130_fd_pr__rf_nfet_01v8_lvt_b__wint_diff=2.252e-8
+  sky130_fd_pr__rf_nfet_01v8_lvt_b__rshg_diff=7.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_b__dlc_diff=-1.1228e-8
+  sky130_fd_pr__rf_nfet_01v8_lvt_b__dwc_diff=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_b__xgw_diff=4.504e-8
+  sky130_fd_pr__rf_nfet_01v8_lvt__aw_cap_mult_p42=1.1125
+  sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_dist_mult_p42=1.245
+  sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_stub_mult_p42=1.245
+  sky130_fd_pr__rf_nfet_01v8_lvt__aw_cap_mult=1.1125
+  sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_dist_mult=1.245
+  sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_stub_mult=1.245
+  sky130_fd_pr__rf_nfet_01v8_lvt__aw_rd_mult=1.0
+  sky130_fd_pr__rf_nfet_01v8_lvt__aw_rs_mult=1.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 000, W = 1.65, L = 0.15
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_0=0.035472
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ags_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_0=-0.0035791
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_0=11669.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b1_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__voff_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b0_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ub_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ua_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__a0_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__pclm_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__kt1_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__nfactor_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__rdsw_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_0=-0.023208
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 001, W = 1.65, L = 0.18
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__kt1_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__nfactor_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__rdsw_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_1=-0.015447
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_1=0.031659
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ags_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_1=-0.0022517
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_1=16627.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b1_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__voff_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b0_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ub_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ua_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__a0_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__pclm_diff_1=0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 002, W = 1.65, L = 0.25
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__kt1_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__nfactor_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__rdsw_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_2=-0.00027242
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_2=0.006014
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ags_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_2=-0.0024036
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_2=7476.5
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b1_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__voff_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b0_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ub_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ua_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__a0_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__pclm_diff_2=0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 003, W = 3.01, L = 0.15
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__pclm_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__kt1_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__nfactor_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__rdsw_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_3=-0.025698
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_3=0.022412
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ags_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_3=-0.0067063
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_3=14950.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b1_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__voff_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b0_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ub_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ua_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__a0_diff_3=0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 004, W = 3.01, L = 0.18
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__pclm_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__kt1_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__nfactor_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__rdsw_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_4=-0.018667
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_4=0.0074967
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ags_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_4=-0.0031604
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_4=14641.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b1_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__voff_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b0_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ub_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ua_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__a0_diff_4=0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 005, W = 3.01, L = 0.25
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__a0_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__pclm_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__kt1_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__nfactor_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__rdsw_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_5=-0.0050153
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_5=0.005408
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ags_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_5=-0.0036655
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_5=14592.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b1_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__voff_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b0_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ub_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ua_diff_5=0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 006, W = 5.05, L = 0.15
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ua_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__a0_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__pclm_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__kt1_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__nfactor_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__rdsw_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_6=-0.031185
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_6=0.019026
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ags_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_6=-0.0097006
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_6=9042.7
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b1_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__voff_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b0_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ub_diff_6=0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 007, W = 5.05, L = 0.18
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ub_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ua_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__a0_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__pclm_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__kt1_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__nfactor_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__rdsw_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_7=-0.018406
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_7=0.005177
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ags_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_7=-0.0054184
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_7=13962.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b1_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__voff_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b0_diff_7=0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 008, W = 5.05, L = 0.25
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__voff_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b0_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ub_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ua_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__a0_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__pclm_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__kt1_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__nfactor_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__rdsw_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_8=-0.0045172
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_8=0.0026993
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ags_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_8=-0.0049523
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_8=16409.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b1_diff_8=0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 000, W = 1.65, L = 0.15
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ua_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__pclm_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__nfactor_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__a0_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__voff_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b0_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_0=-0.022384
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_0=0.032174
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_0=-0.0088162
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_0=18475.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__kt1_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b1_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__rdsw_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ags_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ub_diff_0=0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 001, W = 1.65, L = 0.18
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ags_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ub_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ua_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__pclm_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__nfactor_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__a0_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__voff_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b0_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_1=-0.015672
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_1=0.024627
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_1=-0.0052084
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_1=17204.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__kt1_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b1_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__rdsw_diff_1=0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 002, W = 1.65, L = 0.25
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ags_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ub_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ua_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__pclm_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__nfactor_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__a0_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__voff_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b0_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_2=-0.0053553
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_2=0.00058529
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_2=-0.0047533
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_2=14144.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__kt1_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b1_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__rdsw_diff_2=0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 003, W = 3.01, L = 0.15
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__kt1_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b1_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__rdsw_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ags_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ub_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ua_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__pclm_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__nfactor_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__a0_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__voff_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b0_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_3=-0.026679
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_3=0.025797
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_3=-0.0070348
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_3=14175.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 004, W = 3.01, L = 0.18
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_4=-0.007826
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_4=18436.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__kt1_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b1_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__rdsw_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ags_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ub_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ua_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__pclm_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__nfactor_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__a0_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__voff_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b0_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_4=-0.019062
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_4=0.0093971
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 005, W = 3.01, L = 0.25
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_5=-0.0078718
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_5=-0.0066522
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_5=26781.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__kt1_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b1_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__rdsw_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ags_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ub_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ua_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__pclm_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__nfactor_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__a0_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__voff_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b0_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_5=-0.0060231
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 006, W = 5.05, L = 0.15
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__voff_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b0_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_6=-0.03107
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_6=0.017691
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_6=-0.0077169
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_6=12148.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__kt1_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b1_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__rdsw_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ags_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ub_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ua_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__pclm_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__nfactor_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__a0_diff_6=0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 007, W = 5.05, L = 0.18
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__nfactor_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__a0_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__voff_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b0_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_7=-0.019933
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_7=0.0024544
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_7=-0.0097882
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_7=13883.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__kt1_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b1_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__rdsw_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ags_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ub_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ua_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__pclm_diff_7=0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 008, W = 5.05, L = 0.25
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__pclm_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__nfactor_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__a0_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__voff_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b0_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_8=-0.0057624
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_8=-0.0093065
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_8=39684.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_8=-0.014919
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__kt1_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b1_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__rdsw_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ags_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ub_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ua_diff_8=0.0
.include "sky130_fd_pr__rf_nfet_01v8_lvt_b.pm3.spice"
