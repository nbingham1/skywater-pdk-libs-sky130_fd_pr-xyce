* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 38
.param
+  sky130_fd_pr__nfet_01v8_lvt__toxe_mult=1.052
+  sky130_fd_pr__nfet_01v8_lvt__rshn_mult=1.0
+  sky130_fd_pr__nfet_01v8_lvt__overlap_mult=0.98026
+  sky130_fd_pr__nfet_01v8_lvt__ajunction_mult=1.1755
+  sky130_fd_pr__nfet_01v8_lvt__pjunction_mult=1.0477
+  sky130_fd_pr__nfet_01v8_lvt__lint_diff=-1.7325e-8
+  sky130_fd_pr__nfet_01v8_lvt__wint_diff=3.2175e-8
+  sky130_fd_pr__nfet_01v8_lvt__dlc_diff=-1.5633e-8
+  sky130_fd_pr__nfet_01v8_lvt__dwc_diff=3.2175e-8
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 000, W = 1.0, L = 1.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8_lvt__a0_diff_0=-0.055949
+  sky130_fd_pr__nfet_01v8_lvt__voff_diff_0=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b0_diff_0=0.0
+  sky130_fd_pr__nfet_01v8_lvt__k2_diff_0=0.0085425
+  sky130_fd_pr__nfet_01v8_lvt__u0_diff_0=-0.00221
+  sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_0=0.0
+  sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_0=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ags_diff_0=-0.102
+  sky130_fd_pr__nfet_01v8_lvt__ua_diff_0=-3.9896e-13
+  sky130_fd_pr__nfet_01v8_lvt__vsat_diff_0=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b1_diff_0=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pdits_diff_0=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pclm_diff_0=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ub_diff_0=-4.3129e-20
+  sky130_fd_pr__nfet_01v8_lvt__kt1_diff_0=0.0
+  sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_0=1.0438
+  sky130_fd_pr__nfet_01v8_lvt__keta_diff_0=0.0
+  sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_0=0.0
+  sky130_fd_pr__nfet_01v8_lvt__vth0_diff_0=-0.00077506
+  sky130_fd_pr__nfet_01v8_lvt__eta0_diff_0=0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 001, W = 1.0, L = 2.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8_lvt__eta0_diff_1=0.0
+  sky130_fd_pr__nfet_01v8_lvt__a0_diff_1=-0.070509
+  sky130_fd_pr__nfet_01v8_lvt__voff_diff_1=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b0_diff_1=0.0
+  sky130_fd_pr__nfet_01v8_lvt__k2_diff_1=0.0069185
+  sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_1=0.0
+  sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_1=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ags_diff_1=-0.15419
+  sky130_fd_pr__nfet_01v8_lvt__u0_diff_1=-0.0030873
+  sky130_fd_pr__nfet_01v8_lvt__ua_diff_1=5.5145e-12
+  sky130_fd_pr__nfet_01v8_lvt__vsat_diff_1=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b1_diff_1=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pdits_diff_1=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pclm_diff_1=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ub_diff_1=-1.3823e-20
+  sky130_fd_pr__nfet_01v8_lvt__kt1_diff_1=0.0
+  sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_1=0.3961
+  sky130_fd_pr__nfet_01v8_lvt__keta_diff_1=0.0
+  sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_1=0.0
+  sky130_fd_pr__nfet_01v8_lvt__vth0_diff_1=-0.001839
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 002, W = 1.0, L = 4.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8_lvt__vth0_diff_2=-0.0064743
+  sky130_fd_pr__nfet_01v8_lvt__eta0_diff_2=0.0
+  sky130_fd_pr__nfet_01v8_lvt__a0_diff_2=0.0022663
+  sky130_fd_pr__nfet_01v8_lvt__voff_diff_2=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b0_diff_2=0.0
+  sky130_fd_pr__nfet_01v8_lvt__k2_diff_2=0.009606
+  sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_2=0.0
+  sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_2=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ags_diff_2=0.060976
+  sky130_fd_pr__nfet_01v8_lvt__u0_diff_2=-0.0033168
+  sky130_fd_pr__nfet_01v8_lvt__ua_diff_2=-1.8322e-13
+  sky130_fd_pr__nfet_01v8_lvt__vsat_diff_2=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b1_diff_2=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pdits_diff_2=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pclm_diff_2=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ub_diff_2=-1.0299e-21
+  sky130_fd_pr__nfet_01v8_lvt__kt1_diff_2=0.0
+  sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_2=1.0086
+  sky130_fd_pr__nfet_01v8_lvt__keta_diff_2=0.0
+  sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_2=0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 003, W = 1.0, L = 0.15
* ----------------------------------
+  sky130_fd_pr__nfet_01v8_lvt__kt1_diff_3=0.0
+  sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_3=1.6908
+  sky130_fd_pr__nfet_01v8_lvt__keta_diff_3=0.0
+  sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_3=0.0
+  sky130_fd_pr__nfet_01v8_lvt__vth0_diff_3=0.072735
+  sky130_fd_pr__nfet_01v8_lvt__eta0_diff_3=0.0
+  sky130_fd_pr__nfet_01v8_lvt__a0_diff_3=0.0
+  sky130_fd_pr__nfet_01v8_lvt__voff_diff_3=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b0_diff_3=0.0
+  sky130_fd_pr__nfet_01v8_lvt__k2_diff_3=-0.018829
+  sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_3=0.0
+  sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_3=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ags_diff_3=0.0
+  sky130_fd_pr__nfet_01v8_lvt__u0_diff_3=0.0031047
+  sky130_fd_pr__nfet_01v8_lvt__ua_diff_3=7.7027e-11
+  sky130_fd_pr__nfet_01v8_lvt__vsat_diff_3=31179.0
+  sky130_fd_pr__nfet_01v8_lvt__b1_diff_3=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pdits_diff_3=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pclm_diff_3=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ub_diff_3=3.4943e-20
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 004, W = 1.0, L = 0.18
* ----------------------------------
+  sky130_fd_pr__nfet_01v8_lvt__pdits_diff_4=0.0
+  sky130_fd_pr__nfet_01v8_lvt__kt1_diff_4=0.0
+  sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_4=1.7097
+  sky130_fd_pr__nfet_01v8_lvt__keta_diff_4=0.0
+  sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_4=0.0
+  sky130_fd_pr__nfet_01v8_lvt__vth0_diff_4=0.026404
+  sky130_fd_pr__nfet_01v8_lvt__eta0_diff_4=0.0
+  sky130_fd_pr__nfet_01v8_lvt__a0_diff_4=0.0
+  sky130_fd_pr__nfet_01v8_lvt__voff_diff_4=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b0_diff_4=0.0
+  sky130_fd_pr__nfet_01v8_lvt__k2_diff_4=-0.014357
+  sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_4=0.0
+  sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_4=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ags_diff_4=0.0
+  sky130_fd_pr__nfet_01v8_lvt__u0_diff_4=-0.00066451
+  sky130_fd_pr__nfet_01v8_lvt__ua_diff_4=-5.6442e-12
+  sky130_fd_pr__nfet_01v8_lvt__vsat_diff_4=21392.0
+  sky130_fd_pr__nfet_01v8_lvt__b1_diff_4=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pclm_diff_4=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ub_diff_4=-1.266e-19
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 005, W = 1.0, L = 0.25
* ----------------------------------
+  sky130_fd_pr__nfet_01v8_lvt__pclm_diff_5=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ub_diff_5=-3.145e-19
+  sky130_fd_pr__nfet_01v8_lvt__pdits_diff_5=0.0
+  sky130_fd_pr__nfet_01v8_lvt__kt1_diff_5=0.0
+  sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_5=0.80567
+  sky130_fd_pr__nfet_01v8_lvt__keta_diff_5=0.0
+  sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_5=0.0
+  sky130_fd_pr__nfet_01v8_lvt__vth0_diff_5=0.012126
+  sky130_fd_pr__nfet_01v8_lvt__eta0_diff_5=0.0
+  sky130_fd_pr__nfet_01v8_lvt__a0_diff_5=0.0
+  sky130_fd_pr__nfet_01v8_lvt__voff_diff_5=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b0_diff_5=0.0
+  sky130_fd_pr__nfet_01v8_lvt__k2_diff_5=0.0068689
+  sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_5=0.0
+  sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_5=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ags_diff_5=0.0
+  sky130_fd_pr__nfet_01v8_lvt__u0_diff_5=-0.0062064
+  sky130_fd_pr__nfet_01v8_lvt__ua_diff_5=-3.0184e-11
+  sky130_fd_pr__nfet_01v8_lvt__vsat_diff_5=1072.2
+  sky130_fd_pr__nfet_01v8_lvt__b1_diff_5=0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 006, W = 1.0, L = 0.5
* ---------------------------------
+  sky130_fd_pr__nfet_01v8_lvt__pclm_diff_6=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ub_diff_6=-1.3619e-19
+  sky130_fd_pr__nfet_01v8_lvt__pdits_diff_6=0.0
+  sky130_fd_pr__nfet_01v8_lvt__kt1_diff_6=0.0
+  sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_6=0.9044
+  sky130_fd_pr__nfet_01v8_lvt__keta_diff_6=0.0
+  sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_6=0.0
+  sky130_fd_pr__nfet_01v8_lvt__vth0_diff_6=-0.00022243
+  sky130_fd_pr__nfet_01v8_lvt__eta0_diff_6=0.0
+  sky130_fd_pr__nfet_01v8_lvt__a0_diff_6=0.0
+  sky130_fd_pr__nfet_01v8_lvt__voff_diff_6=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b0_diff_6=0.0
+  sky130_fd_pr__nfet_01v8_lvt__k2_diff_6=0.004307
+  sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_6=0.0
+  sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_6=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ags_diff_6=0.0
+  sky130_fd_pr__nfet_01v8_lvt__u0_diff_6=-0.0019441
+  sky130_fd_pr__nfet_01v8_lvt__ua_diff_6=-1.4067e-11
+  sky130_fd_pr__nfet_01v8_lvt__vsat_diff_6=28850.0
+  sky130_fd_pr__nfet_01v8_lvt__b1_diff_6=0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 007, W = 3.0, L = 1.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8_lvt__b1_diff_7=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pclm_diff_7=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ub_diff_7=9.2338e-21
+  sky130_fd_pr__nfet_01v8_lvt__pdits_diff_7=0.0
+  sky130_fd_pr__nfet_01v8_lvt__kt1_diff_7=0.0
+  sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_7=0.91994
+  sky130_fd_pr__nfet_01v8_lvt__keta_diff_7=0.0
+  sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_7=0.0
+  sky130_fd_pr__nfet_01v8_lvt__vth0_diff_7=0.00047059
+  sky130_fd_pr__nfet_01v8_lvt__eta0_diff_7=0.0
+  sky130_fd_pr__nfet_01v8_lvt__a0_diff_7=-0.0728
+  sky130_fd_pr__nfet_01v8_lvt__voff_diff_7=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b0_diff_7=0.0
+  sky130_fd_pr__nfet_01v8_lvt__k2_diff_7=0.0063087
+  sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_7=0.0
+  sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_7=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ags_diff_7=-0.092159
+  sky130_fd_pr__nfet_01v8_lvt__u0_diff_7=7.7658e-5
+  sky130_fd_pr__nfet_01v8_lvt__ua_diff_7=-1.7373e-12
+  sky130_fd_pr__nfet_01v8_lvt__vsat_diff_7=0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 008, W = 3.0, L = 2.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_8=0.0
+  sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_8=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ags_diff_8=-0.11278
+  sky130_fd_pr__nfet_01v8_lvt__u0_diff_8=0.0005698
+  sky130_fd_pr__nfet_01v8_lvt__ua_diff_8=3.5055e-13
+  sky130_fd_pr__nfet_01v8_lvt__vsat_diff_8=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b1_diff_8=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pclm_diff_8=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ub_diff_8=1.1995e-19
+  sky130_fd_pr__nfet_01v8_lvt__pdits_diff_8=0.0
+  sky130_fd_pr__nfet_01v8_lvt__kt1_diff_8=0.0
+  sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_8=0.41301
+  sky130_fd_pr__nfet_01v8_lvt__keta_diff_8=0.0
+  sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_8=0.0
+  sky130_fd_pr__nfet_01v8_lvt__vth0_diff_8=-0.0063199
+  sky130_fd_pr__nfet_01v8_lvt__eta0_diff_8=0.0
+  sky130_fd_pr__nfet_01v8_lvt__a0_diff_8=-0.073197
+  sky130_fd_pr__nfet_01v8_lvt__voff_diff_8=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b0_diff_8=0.0
+  sky130_fd_pr__nfet_01v8_lvt__k2_diff_8=0.0051108
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 009, W = 3.0, L = 4.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_9=0.0
+  sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_9=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ags_diff_9=-0.0084268
+  sky130_fd_pr__nfet_01v8_lvt__u0_diff_9=-0.0003352
+  sky130_fd_pr__nfet_01v8_lvt__ua_diff_9=-1.3364e-12
+  sky130_fd_pr__nfet_01v8_lvt__vsat_diff_9=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b1_diff_9=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pclm_diff_9=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ub_diff_9=4.2918e-20
+  sky130_fd_pr__nfet_01v8_lvt__pdits_diff_9=0.0
+  sky130_fd_pr__nfet_01v8_lvt__kt1_diff_9=0.0
+  sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_9=0.58828
+  sky130_fd_pr__nfet_01v8_lvt__keta_diff_9=0.0
+  sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_9=0.0
+  sky130_fd_pr__nfet_01v8_lvt__vth0_diff_9=-0.0055555
+  sky130_fd_pr__nfet_01v8_lvt__eta0_diff_9=0.0
+  sky130_fd_pr__nfet_01v8_lvt__a0_diff_9=0.0081032
+  sky130_fd_pr__nfet_01v8_lvt__voff_diff_9=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b0_diff_9=0.0
+  sky130_fd_pr__nfet_01v8_lvt__k2_diff_9=0.0072177
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 010, W = 3.0, L = 0.15
* ----------------------------------
+  sky130_fd_pr__nfet_01v8_lvt__pdits_diff_10=0.0
+  sky130_fd_pr__nfet_01v8_lvt__eta0_diff_10=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ua_diff_10=-4.6287e-12
+  sky130_fd_pr__nfet_01v8_lvt__ub_diff_10=-2.4778e-21
+  sky130_fd_pr__nfet_01v8_lvt__a0_diff_10=0.0
+  sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_10=0.0
+  sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_10=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ags_diff_10=0.0
+  sky130_fd_pr__nfet_01v8_lvt__u0_diff_10=-0.00062201
+  sky130_fd_pr__nfet_01v8_lvt__vsat_diff_10=27925.0
+  sky130_fd_pr__nfet_01v8_lvt__vth0_diff_10=0.017771
+  sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_10=1.5215
+  sky130_fd_pr__nfet_01v8_lvt__kt1_diff_10=0.0
+  sky130_fd_pr__nfet_01v8_lvt__voff_diff_10=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b0_diff_10=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b1_diff_10=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_10=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pclm_diff_10=0.0
+  sky130_fd_pr__nfet_01v8_lvt__keta_diff_10=0.0
+  sky130_fd_pr__nfet_01v8_lvt__k2_diff_10=-0.022548
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 011, W = 3.0, L = 0.18
* ----------------------------------
+  sky130_fd_pr__nfet_01v8_lvt__keta_diff_11=0.0
+  sky130_fd_pr__nfet_01v8_lvt__k2_diff_11=-0.015748
+  sky130_fd_pr__nfet_01v8_lvt__pdits_diff_11=0.0
+  sky130_fd_pr__nfet_01v8_lvt__eta0_diff_11=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ua_diff_11=-1.308e-11
+  sky130_fd_pr__nfet_01v8_lvt__ub_diff_11=9.2336e-20
+  sky130_fd_pr__nfet_01v8_lvt__a0_diff_11=0.0
+  sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_11=0.0
+  sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_11=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ags_diff_11=0.0
+  sky130_fd_pr__nfet_01v8_lvt__u0_diff_11=0.0012153
+  sky130_fd_pr__nfet_01v8_lvt__vsat_diff_11=22649.0
+  sky130_fd_pr__nfet_01v8_lvt__vth0_diff_11=0.021254
+  sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_11=1.5828
+  sky130_fd_pr__nfet_01v8_lvt__kt1_diff_11=0.0
+  sky130_fd_pr__nfet_01v8_lvt__voff_diff_11=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b0_diff_11=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b1_diff_11=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_11=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pclm_diff_11=0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 012, W = 3.0, L = 0.25
* ----------------------------------
+  sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_12=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pclm_diff_12=0.0
+  sky130_fd_pr__nfet_01v8_lvt__keta_diff_12=0.0
+  sky130_fd_pr__nfet_01v8_lvt__k2_diff_12=0.0020207
+  sky130_fd_pr__nfet_01v8_lvt__pdits_diff_12=0.0
+  sky130_fd_pr__nfet_01v8_lvt__eta0_diff_12=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ua_diff_12=-2.023e-10
+  sky130_fd_pr__nfet_01v8_lvt__ub_diff_12=9.3908e-20
+  sky130_fd_pr__nfet_01v8_lvt__a0_diff_12=0.0
+  sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_12=0.0
+  sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_12=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ags_diff_12=0.0
+  sky130_fd_pr__nfet_01v8_lvt__u0_diff_12=-0.0050513
+  sky130_fd_pr__nfet_01v8_lvt__vsat_diff_12=22072.0
+  sky130_fd_pr__nfet_01v8_lvt__vth0_diff_12=0.011709
+  sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_12=1.0754
+  sky130_fd_pr__nfet_01v8_lvt__kt1_diff_12=0.0
+  sky130_fd_pr__nfet_01v8_lvt__voff_diff_12=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b0_diff_12=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b1_diff_12=0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 013, W = 3.0, L = 0.5
* ---------------------------------
+  sky130_fd_pr__nfet_01v8_lvt__b1_diff_13=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_13=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pclm_diff_13=0.0
+  sky130_fd_pr__nfet_01v8_lvt__keta_diff_13=0.0
+  sky130_fd_pr__nfet_01v8_lvt__k2_diff_13=0.009986
+  sky130_fd_pr__nfet_01v8_lvt__pdits_diff_13=0.0
+  sky130_fd_pr__nfet_01v8_lvt__eta0_diff_13=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ua_diff_13=-4.0028e-12
+  sky130_fd_pr__nfet_01v8_lvt__ub_diff_13=9.0364e-20
+  sky130_fd_pr__nfet_01v8_lvt__a0_diff_13=0.0
+  sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_13=0.0
+  sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_13=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ags_diff_13=0.0
+  sky130_fd_pr__nfet_01v8_lvt__u0_diff_13=0.0012156
+  sky130_fd_pr__nfet_01v8_lvt__vsat_diff_13=22472.0
+  sky130_fd_pr__nfet_01v8_lvt__vth0_diff_13=0.0015895
+  sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_13=1.2534
+  sky130_fd_pr__nfet_01v8_lvt__kt1_diff_13=0.0
+  sky130_fd_pr__nfet_01v8_lvt__voff_diff_13=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b0_diff_13=0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 014, W = 5.0, L = 1.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8_lvt__kt1_diff_14=0.0
+  sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_14=0.74152
+  sky130_fd_pr__nfet_01v8_lvt__voff_diff_14=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b0_diff_14=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b1_diff_14=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_14=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pclm_diff_14=0.0
+  sky130_fd_pr__nfet_01v8_lvt__keta_diff_14=0.0
+  sky130_fd_pr__nfet_01v8_lvt__k2_diff_14=0.003644
+  sky130_fd_pr__nfet_01v8_lvt__pdits_diff_14=0.0
+  sky130_fd_pr__nfet_01v8_lvt__eta0_diff_14=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ua_diff_14=-1.6542e-12
+  sky130_fd_pr__nfet_01v8_lvt__ub_diff_14=1.0391e-19
+  sky130_fd_pr__nfet_01v8_lvt__a0_diff_14=-0.072509
+  sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_14=0.0
+  sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_14=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ags_diff_14=-0.10562
+  sky130_fd_pr__nfet_01v8_lvt__u0_diff_14=0.0012428
+  sky130_fd_pr__nfet_01v8_lvt__vsat_diff_14=0.0
+  sky130_fd_pr__nfet_01v8_lvt__vth0_diff_14=-0.0046668
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 015, W = 5.0, L = 2.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8_lvt__vth0_diff_15=-0.0019576
+  sky130_fd_pr__nfet_01v8_lvt__kt1_diff_15=0.0
+  sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_15=0.75726
+  sky130_fd_pr__nfet_01v8_lvt__voff_diff_15=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b0_diff_15=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b1_diff_15=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_15=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pclm_diff_15=0.0
+  sky130_fd_pr__nfet_01v8_lvt__keta_diff_15=0.0
+  sky130_fd_pr__nfet_01v8_lvt__k2_diff_15=-0.0056244
+  sky130_fd_pr__nfet_01v8_lvt__pdits_diff_15=0.0
+  sky130_fd_pr__nfet_01v8_lvt__eta0_diff_15=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ua_diff_15=-2.2616e-12
+  sky130_fd_pr__nfet_01v8_lvt__ub_diff_15=9.0863e-20
+  sky130_fd_pr__nfet_01v8_lvt__a0_diff_15=-0.01554
+  sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_15=0.0
+  sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_15=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ags_diff_15=-0.05945
+  sky130_fd_pr__nfet_01v8_lvt__u0_diff_15=0.00070865
+  sky130_fd_pr__nfet_01v8_lvt__vsat_diff_15=0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 016, W = 5.0, L = 4.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_16=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ags_diff_16=-0.067693
+  sky130_fd_pr__nfet_01v8_lvt__u0_diff_16=0.00049371
+  sky130_fd_pr__nfet_01v8_lvt__vsat_diff_16=0.0
+  sky130_fd_pr__nfet_01v8_lvt__vth0_diff_16=-0.005429
+  sky130_fd_pr__nfet_01v8_lvt__kt1_diff_16=0.0
+  sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_16=0.18234
+  sky130_fd_pr__nfet_01v8_lvt__voff_diff_16=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b0_diff_16=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b1_diff_16=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_16=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pclm_diff_16=0.0
+  sky130_fd_pr__nfet_01v8_lvt__keta_diff_16=0.0
+  sky130_fd_pr__nfet_01v8_lvt__k2_diff_16=0.011012
+  sky130_fd_pr__nfet_01v8_lvt__pdits_diff_16=0.0
+  sky130_fd_pr__nfet_01v8_lvt__eta0_diff_16=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ua_diff_16=-4.1373e-13
+  sky130_fd_pr__nfet_01v8_lvt__ub_diff_16=9.5675e-20
+  sky130_fd_pr__nfet_01v8_lvt__a0_diff_16=0.011858
+  sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_16=0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 017, W = 5.0, L = 0.15
* ----------------------------------
+  sky130_fd_pr__nfet_01v8_lvt__a0_diff_17=0.0
+  sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_17=0.0
+  sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_17=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ags_diff_17=0.0
+  sky130_fd_pr__nfet_01v8_lvt__u0_diff_17=0.0021031
+  sky130_fd_pr__nfet_01v8_lvt__vsat_diff_17=30122.0
+  sky130_fd_pr__nfet_01v8_lvt__vth0_diff_17=0.029097
+  sky130_fd_pr__nfet_01v8_lvt__kt1_diff_17=0.0
+  sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_17=1.5408
+  sky130_fd_pr__nfet_01v8_lvt__voff_diff_17=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b0_diff_17=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b1_diff_17=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_17=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pclm_diff_17=0.0
+  sky130_fd_pr__nfet_01v8_lvt__keta_diff_17=0.0
+  sky130_fd_pr__nfet_01v8_lvt__k2_diff_17=-0.025776
+  sky130_fd_pr__nfet_01v8_lvt__pdits_diff_17=0.0
+  sky130_fd_pr__nfet_01v8_lvt__eta0_diff_17=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ua_diff_17=-2.1527e-11
+  sky130_fd_pr__nfet_01v8_lvt__ub_diff_17=2.4033e-19
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 018, W = 5.0, L = 0.18
* ----------------------------------
+  sky130_fd_pr__nfet_01v8_lvt__a0_diff_18=0.0
+  sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_18=0.0
+  sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_18=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ags_diff_18=0.0
+  sky130_fd_pr__nfet_01v8_lvt__u0_diff_18=0.00070574
+  sky130_fd_pr__nfet_01v8_lvt__vsat_diff_18=15222.0
+  sky130_fd_pr__nfet_01v8_lvt__vth0_diff_18=0.031285
+  sky130_fd_pr__nfet_01v8_lvt__kt1_diff_18=0.0
+  sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_18=1.357
+  sky130_fd_pr__nfet_01v8_lvt__voff_diff_18=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b0_diff_18=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b1_diff_18=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_18=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pclm_diff_18=0.0
+  sky130_fd_pr__nfet_01v8_lvt__keta_diff_18=0.0
+  sky130_fd_pr__nfet_01v8_lvt__k2_diff_18=-0.014864
+  sky130_fd_pr__nfet_01v8_lvt__pdits_diff_18=0.0
+  sky130_fd_pr__nfet_01v8_lvt__eta0_diff_18=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ua_diff_18=-9.7118e-12
+  sky130_fd_pr__nfet_01v8_lvt__ub_diff_18=1.1272e-19
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 019, W = 5.0, L = 0.25
* ----------------------------------
+  sky130_fd_pr__nfet_01v8_lvt__ub_diff_19=-1.1316e-19
+  sky130_fd_pr__nfet_01v8_lvt__a0_diff_19=0.0
+  sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_19=0.0
+  sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_19=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ags_diff_19=0.0
+  sky130_fd_pr__nfet_01v8_lvt__u0_diff_19=-0.0059387
+  sky130_fd_pr__nfet_01v8_lvt__vsat_diff_19=13387.0
+  sky130_fd_pr__nfet_01v8_lvt__vth0_diff_19=-0.0025422
+  sky130_fd_pr__nfet_01v8_lvt__kt1_diff_19=0.0
+  sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_19=1.3025
+  sky130_fd_pr__nfet_01v8_lvt__voff_diff_19=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b0_diff_19=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b1_diff_19=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_19=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pclm_diff_19=0.0
+  sky130_fd_pr__nfet_01v8_lvt__keta_diff_19=0.0
+  sky130_fd_pr__nfet_01v8_lvt__k2_diff_19=-0.00025623
+  sky130_fd_pr__nfet_01v8_lvt__pdits_diff_19=0.0
+  sky130_fd_pr__nfet_01v8_lvt__eta0_diff_19=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ua_diff_19=-6.7249e-11
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 020, W = 5.0, L = 0.5
* ---------------------------------
+  sky130_fd_pr__nfet_01v8_lvt__pdits_diff_20=0.0
+  sky130_fd_pr__nfet_01v8_lvt__eta0_diff_20=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ua_diff_20=-6.3489e-12
+  sky130_fd_pr__nfet_01v8_lvt__ub_diff_20=2.1234e-19
+  sky130_fd_pr__nfet_01v8_lvt__a0_diff_20=0.0
+  sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_20=0.0
+  sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_20=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ags_diff_20=0.0
+  sky130_fd_pr__nfet_01v8_lvt__u0_diff_20=0.0029292
+  sky130_fd_pr__nfet_01v8_lvt__vsat_diff_20=20921.0
+  sky130_fd_pr__nfet_01v8_lvt__vth0_diff_20=-0.0055971
+  sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_20=0.86492
+  sky130_fd_pr__nfet_01v8_lvt__kt1_diff_20=0.0
+  sky130_fd_pr__nfet_01v8_lvt__voff_diff_20=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b0_diff_20=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b1_diff_20=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_20=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pclm_diff_20=0.0
+  sky130_fd_pr__nfet_01v8_lvt__keta_diff_20=0.0
+  sky130_fd_pr__nfet_01v8_lvt__k2_diff_20=0.0045468
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 021, W = 7.0, L = 1.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8_lvt__pdits_diff_21=0.0
+  sky130_fd_pr__nfet_01v8_lvt__eta0_diff_21=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ua_diff_21=-2.7516e-12
+  sky130_fd_pr__nfet_01v8_lvt__ub_diff_21=1.2551e-19
+  sky130_fd_pr__nfet_01v8_lvt__a0_diff_21=-0.04154
+  sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_21=0.0
+  sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_21=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ags_diff_21=-0.057513
+  sky130_fd_pr__nfet_01v8_lvt__u0_diff_21=0.0014822
+  sky130_fd_pr__nfet_01v8_lvt__vsat_diff_21=0.0
+  sky130_fd_pr__nfet_01v8_lvt__vth0_diff_21=0.00081499
+  sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_21=0.74746
+  sky130_fd_pr__nfet_01v8_lvt__kt1_diff_21=0.0
+  sky130_fd_pr__nfet_01v8_lvt__voff_diff_21=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b0_diff_21=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b1_diff_21=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_21=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pclm_diff_21=0.0
+  sky130_fd_pr__nfet_01v8_lvt__keta_diff_21=0.0
+  sky130_fd_pr__nfet_01v8_lvt__k2_diff_21=-0.0021479
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 022, W = 7.0, L = 2.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8_lvt__keta_diff_22=0.0
+  sky130_fd_pr__nfet_01v8_lvt__k2_diff_22=0.0097484
+  sky130_fd_pr__nfet_01v8_lvt__pdits_diff_22=0.0
+  sky130_fd_pr__nfet_01v8_lvt__eta0_diff_22=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ua_diff_22=-9.3121e-13
+  sky130_fd_pr__nfet_01v8_lvt__ub_diff_22=9.5373e-20
+  sky130_fd_pr__nfet_01v8_lvt__a0_diff_22=-0.044389
+  sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_22=0.0
+  sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_22=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ags_diff_22=-0.11382
+  sky130_fd_pr__nfet_01v8_lvt__u0_diff_22=0.00081875
+  sky130_fd_pr__nfet_01v8_lvt__vsat_diff_22=0.0
+  sky130_fd_pr__nfet_01v8_lvt__vth0_diff_22=-0.0037978
+  sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_22=0.53425
+  sky130_fd_pr__nfet_01v8_lvt__kt1_diff_22=0.0
+  sky130_fd_pr__nfet_01v8_lvt__voff_diff_22=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b0_diff_22=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b1_diff_22=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_22=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pclm_diff_22=0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 023, W = 7.0, L = 8.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_23=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pclm_diff_23=0.0
+  sky130_fd_pr__nfet_01v8_lvt__keta_diff_23=0.0
+  sky130_fd_pr__nfet_01v8_lvt__k2_diff_23=0.0086791
+  sky130_fd_pr__nfet_01v8_lvt__pdits_diff_23=0.0
+  sky130_fd_pr__nfet_01v8_lvt__eta0_diff_23=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ua_diff_23=-2.7497e-12
+  sky130_fd_pr__nfet_01v8_lvt__ub_diff_23=1.6993e-19
+  sky130_fd_pr__nfet_01v8_lvt__a0_diff_23=0.0068567
+  sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_23=0.0
+  sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_23=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ags_diff_23=-0.0077843
+  sky130_fd_pr__nfet_01v8_lvt__u0_diff_23=0.00097538
+  sky130_fd_pr__nfet_01v8_lvt__vsat_diff_23=0.0
+  sky130_fd_pr__nfet_01v8_lvt__vth0_diff_23=-0.0037087
+  sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_23=0.44392
+  sky130_fd_pr__nfet_01v8_lvt__kt1_diff_23=0.0
+  sky130_fd_pr__nfet_01v8_lvt__voff_diff_23=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b0_diff_23=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b1_diff_23=0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 024, W = 7.0, L = 0.15
* ----------------------------------
+  sky130_fd_pr__nfet_01v8_lvt__b1_diff_24=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_24=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pclm_diff_24=0.0
+  sky130_fd_pr__nfet_01v8_lvt__keta_diff_24=0.0
+  sky130_fd_pr__nfet_01v8_lvt__k2_diff_24=-0.016515
+  sky130_fd_pr__nfet_01v8_lvt__pdits_diff_24=0.0
+  sky130_fd_pr__nfet_01v8_lvt__eta0_diff_24=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ua_diff_24=-6.0124e-14
+  sky130_fd_pr__nfet_01v8_lvt__ub_diff_24=-1.4258e-19
+  sky130_fd_pr__nfet_01v8_lvt__a0_diff_24=0.0
+  sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_24=0.0
+  sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_24=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ags_diff_24=0.0
+  sky130_fd_pr__nfet_01v8_lvt__u0_diff_24=-0.0016337
+  sky130_fd_pr__nfet_01v8_lvt__vsat_diff_24=21107.0
+  sky130_fd_pr__nfet_01v8_lvt__vth0_diff_24=0.011419
+  sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_24=1.5827
+  sky130_fd_pr__nfet_01v8_lvt__kt1_diff_24=0.0
+  sky130_fd_pr__nfet_01v8_lvt__voff_diff_24=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b0_diff_24=0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 025, W = 7.0, L = 0.18
* ----------------------------------
+  sky130_fd_pr__nfet_01v8_lvt__kt1_diff_25=0.0
+  sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_25=1.361
+  sky130_fd_pr__nfet_01v8_lvt__voff_diff_25=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b0_diff_25=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b1_diff_25=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_25=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pclm_diff_25=0.0
+  sky130_fd_pr__nfet_01v8_lvt__keta_diff_25=0.0
+  sky130_fd_pr__nfet_01v8_lvt__k2_diff_25=-0.0079681
+  sky130_fd_pr__nfet_01v8_lvt__pdits_diff_25=0.0
+  sky130_fd_pr__nfet_01v8_lvt__eta0_diff_25=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ua_diff_25=-1.2769e-12
+  sky130_fd_pr__nfet_01v8_lvt__ub_diff_25=2.4405e-19
+  sky130_fd_pr__nfet_01v8_lvt__a0_diff_25=0.0
+  sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_25=0.0
+  sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_25=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ags_diff_25=0.0
+  sky130_fd_pr__nfet_01v8_lvt__u0_diff_25=0.0021332
+  sky130_fd_pr__nfet_01v8_lvt__vsat_diff_25=22840.0
+  sky130_fd_pr__nfet_01v8_lvt__vth0_diff_25=0.0030577
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 026, W = 7.0, L = 0.25
* ----------------------------------
+  sky130_fd_pr__nfet_01v8_lvt__vth0_diff_26=-0.006733
+  sky130_fd_pr__nfet_01v8_lvt__kt1_diff_26=0.0
+  sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_26=1.3641
+  sky130_fd_pr__nfet_01v8_lvt__voff_diff_26=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b0_diff_26=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b1_diff_26=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_26=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pclm_diff_26=0.0
+  sky130_fd_pr__nfet_01v8_lvt__keta_diff_26=0.0
+  sky130_fd_pr__nfet_01v8_lvt__k2_diff_26=0.0013271
+  sky130_fd_pr__nfet_01v8_lvt__pdits_diff_26=0.0
+  sky130_fd_pr__nfet_01v8_lvt__eta0_diff_26=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ua_diff_26=2.3431e-12
+  sky130_fd_pr__nfet_01v8_lvt__ub_diff_26=6.2679e-20
+  sky130_fd_pr__nfet_01v8_lvt__a0_diff_26=0.0
+  sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_26=0.0
+  sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_26=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ags_diff_26=0.0
+  sky130_fd_pr__nfet_01v8_lvt__u0_diff_26=-0.003233
+  sky130_fd_pr__nfet_01v8_lvt__vsat_diff_26=30699.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 027, W = 7.0, L = 0.5
* ---------------------------------
+  sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_27=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ags_diff_27=0.0
+  sky130_fd_pr__nfet_01v8_lvt__u0_diff_27=0.0021917
+  sky130_fd_pr__nfet_01v8_lvt__vsat_diff_27=2182.4
+  sky130_fd_pr__nfet_01v8_lvt__vth0_diff_27=-0.00052024
+  sky130_fd_pr__nfet_01v8_lvt__kt1_diff_27=0.0
+  sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_27=1.1854
+  sky130_fd_pr__nfet_01v8_lvt__voff_diff_27=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b0_diff_27=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b1_diff_27=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_27=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pclm_diff_27=0.0
+  sky130_fd_pr__nfet_01v8_lvt__keta_diff_27=0.0
+  sky130_fd_pr__nfet_01v8_lvt__k2_diff_27=0.0042372
+  sky130_fd_pr__nfet_01v8_lvt__pdits_diff_27=0.0
+  sky130_fd_pr__nfet_01v8_lvt__eta0_diff_27=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ua_diff_27=-5.9962e-12
+  sky130_fd_pr__nfet_01v8_lvt__ub_diff_27=1.8543e-19
+  sky130_fd_pr__nfet_01v8_lvt__a0_diff_27=0.0
+  sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_27=0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 028, W = 0.42, L = 1.0
* ----------------------------------
+  sky130_fd_pr__nfet_01v8_lvt__a0_diff_28=0.0
+  sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_28=0.0
+  sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_28=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ags_diff_28=0.0
+  sky130_fd_pr__nfet_01v8_lvt__u0_diff_28=-0.0098936
+  sky130_fd_pr__nfet_01v8_lvt__vsat_diff_28=0.0
+  sky130_fd_pr__nfet_01v8_lvt__vth0_diff_28=-0.00673
+  sky130_fd_pr__nfet_01v8_lvt__kt1_diff_28=0.0
+  sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_28=0.78389
+  sky130_fd_pr__nfet_01v8_lvt__voff_diff_28=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b0_diff_28=5.58e-8
+  sky130_fd_pr__nfet_01v8_lvt__b1_diff_28=1.5703e-8
+  sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_28=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pclm_diff_28=0.0
+  sky130_fd_pr__nfet_01v8_lvt__keta_diff_28=0.0
+  sky130_fd_pr__nfet_01v8_lvt__k2_diff_28=0.0030676
+  sky130_fd_pr__nfet_01v8_lvt__pdits_diff_28=0.0
+  sky130_fd_pr__nfet_01v8_lvt__eta0_diff_28=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ua_diff_28=2.5848e-12
+  sky130_fd_pr__nfet_01v8_lvt__ub_diff_28=-4.1546e-19
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 029, W = 0.42, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8_lvt__a0_diff_29=0.0
+  sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_29=0.0
+  sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_29=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ags_diff_29=0.0
+  sky130_fd_pr__nfet_01v8_lvt__u0_diff_29=-0.00066428
+  sky130_fd_pr__nfet_01v8_lvt__vsat_diff_29=59754.0
+  sky130_fd_pr__nfet_01v8_lvt__vth0_diff_29=0.08747
+  sky130_fd_pr__nfet_01v8_lvt__kt1_diff_29=0.0
+  sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_29=1.6311
+  sky130_fd_pr__nfet_01v8_lvt__voff_diff_29=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b0_diff_29=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b1_diff_29=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_29=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pclm_diff_29=0.0
+  sky130_fd_pr__nfet_01v8_lvt__keta_diff_29=0.0
+  sky130_fd_pr__nfet_01v8_lvt__k2_diff_29=-0.020075
+  sky130_fd_pr__nfet_01v8_lvt__pdits_diff_29=0.0
+  sky130_fd_pr__nfet_01v8_lvt__eta0_diff_29=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ua_diff_29=-7.4884e-12
+  sky130_fd_pr__nfet_01v8_lvt__ub_diff_29=-2.6145e-19
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 030, W = 0.42, L = 0.18
* -----------------------------------
+  sky130_fd_pr__nfet_01v8_lvt__ub_diff_30=1.3839e-20
+  sky130_fd_pr__nfet_01v8_lvt__a0_diff_30=0.0
+  sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_30=0.0
+  sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_30=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ags_diff_30=0.0
+  sky130_fd_pr__nfet_01v8_lvt__u0_diff_30=0.0012542
+  sky130_fd_pr__nfet_01v8_lvt__vsat_diff_30=34097.0
+  sky130_fd_pr__nfet_01v8_lvt__vth0_diff_30=0.03095
+  sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_30=1.3955
+  sky130_fd_pr__nfet_01v8_lvt__kt1_diff_30=0.0
+  sky130_fd_pr__nfet_01v8_lvt__voff_diff_30=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b0_diff_30=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b1_diff_30=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_30=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pclm_diff_30=0.0
+  sky130_fd_pr__nfet_01v8_lvt__keta_diff_30=0.0
+  sky130_fd_pr__nfet_01v8_lvt__k2_diff_30=-0.0099934
+  sky130_fd_pr__nfet_01v8_lvt__ua_diff_30=-1.26e-11
+  sky130_fd_pr__nfet_01v8_lvt__pdits_diff_30=0.0
+  sky130_fd_pr__nfet_01v8_lvt__eta0_diff_30=0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 031, W = 0.55, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8_lvt__pdits_diff_31=0.0
+  sky130_fd_pr__nfet_01v8_lvt__eta0_diff_31=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ua_diff_31=-1.5783e-12
+  sky130_fd_pr__nfet_01v8_lvt__ub_diff_31=-1.6453e-19
+  sky130_fd_pr__nfet_01v8_lvt__a0_diff_31=0.0
+  sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_31=0.0
+  sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_31=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ags_diff_31=0.0
+  sky130_fd_pr__nfet_01v8_lvt__u0_diff_31=-0.00055666
+  sky130_fd_pr__nfet_01v8_lvt__vsat_diff_31=58025.0
+  sky130_fd_pr__nfet_01v8_lvt__vth0_diff_31=0.10909
+  sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_31=1.7747
+  sky130_fd_pr__nfet_01v8_lvt__kt1_diff_31=0.0
+  sky130_fd_pr__nfet_01v8_lvt__voff_diff_31=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b0_diff_31=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b1_diff_31=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_31=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pclm_diff_31=0.0
+  sky130_fd_pr__nfet_01v8_lvt__keta_diff_31=0.0
+  sky130_fd_pr__nfet_01v8_lvt__k2_diff_31=-0.014266
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 032, W = 0.64, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8_lvt__pdits_diff_32=0.0
+  sky130_fd_pr__nfet_01v8_lvt__eta0_diff_32=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ua_diff_32=-5.3029e-12
+  sky130_fd_pr__nfet_01v8_lvt__ub_diff_32=-4.4441e-19
+  sky130_fd_pr__nfet_01v8_lvt__a0_diff_32=0.0
+  sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_32=0.0
+  sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_32=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ags_diff_32=0.0
+  sky130_fd_pr__nfet_01v8_lvt__u0_diff_32=-0.0019696
+  sky130_fd_pr__nfet_01v8_lvt__vsat_diff_32=27382.0
+  sky130_fd_pr__nfet_01v8_lvt__vth0_diff_32=0.093609
+  sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_32=2.0551
+  sky130_fd_pr__nfet_01v8_lvt__kt1_diff_32=0.0
+  sky130_fd_pr__nfet_01v8_lvt__voff_diff_32=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b0_diff_32=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b1_diff_32=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_32=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pclm_diff_32=0.0
+  sky130_fd_pr__nfet_01v8_lvt__keta_diff_32=0.0
+  sky130_fd_pr__nfet_01v8_lvt__k2_diff_32=-0.016503
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 033, W = 0.84, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8_lvt__keta_diff_33=0.0
+  sky130_fd_pr__nfet_01v8_lvt__k2_diff_33=-0.017098
+  sky130_fd_pr__nfet_01v8_lvt__pdits_diff_33=0.0
+  sky130_fd_pr__nfet_01v8_lvt__eta0_diff_33=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ua_diff_33=-3.3781e-12
+  sky130_fd_pr__nfet_01v8_lvt__ub_diff_33=-3.1236e-19
+  sky130_fd_pr__nfet_01v8_lvt__a0_diff_33=0.0
+  sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_33=0.0
+  sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_33=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ags_diff_33=0.0
+  sky130_fd_pr__nfet_01v8_lvt__u0_diff_33=-0.0013071
+  sky130_fd_pr__nfet_01v8_lvt__vsat_diff_33=24130.0
+  sky130_fd_pr__nfet_01v8_lvt__vth0_diff_33=0.099
+  sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_33=2.0077
+  sky130_fd_pr__nfet_01v8_lvt__kt1_diff_33=0.0
+  sky130_fd_pr__nfet_01v8_lvt__voff_diff_33=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b0_diff_33=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b1_diff_33=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_33=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pclm_diff_33=0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 034, W = 1.65, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_34=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pclm_diff_34=0.0
+  sky130_fd_pr__nfet_01v8_lvt__keta_diff_34=0.0
+  sky130_fd_pr__nfet_01v8_lvt__k2_diff_34=-0.016502
+  sky130_fd_pr__nfet_01v8_lvt__pdits_diff_34=0.0
+  sky130_fd_pr__nfet_01v8_lvt__eta0_diff_34=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ua_diff_34=8.7643e-13
+  sky130_fd_pr__nfet_01v8_lvt__ub_diff_34=-1.3074e-19
+  sky130_fd_pr__nfet_01v8_lvt__a0_diff_34=0.0
+  sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_34=0.0
+  sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_34=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ags_diff_34=0.0
+  sky130_fd_pr__nfet_01v8_lvt__u0_diff_34=-0.0012865
+  sky130_fd_pr__nfet_01v8_lvt__vsat_diff_34=28542.0
+  sky130_fd_pr__nfet_01v8_lvt__vth0_diff_34=0.052168
+  sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_34=1.1539
+  sky130_fd_pr__nfet_01v8_lvt__kt1_diff_34=0.0
+  sky130_fd_pr__nfet_01v8_lvt__voff_diff_34=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b0_diff_34=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b1_diff_34=0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 035, W = 3.01, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8_lvt__b1_diff_35=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_35=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pclm_diff_35=0.0
+  sky130_fd_pr__nfet_01v8_lvt__keta_diff_35=0.0
+  sky130_fd_pr__nfet_01v8_lvt__k2_diff_35=-0.023286
+  sky130_fd_pr__nfet_01v8_lvt__pdits_diff_35=0.0
+  sky130_fd_pr__nfet_01v8_lvt__eta0_diff_35=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ua_diff_35=-2.8889e-14
+  sky130_fd_pr__nfet_01v8_lvt__ub_diff_35=-1.8324e-20
+  sky130_fd_pr__nfet_01v8_lvt__a0_diff_35=0.0
+  sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_35=0.0
+  sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_35=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ags_diff_35=0.0
+  sky130_fd_pr__nfet_01v8_lvt__u0_diff_35=-0.00053862
+  sky130_fd_pr__nfet_01v8_lvt__vsat_diff_35=23966.0
+  sky130_fd_pr__nfet_01v8_lvt__vth0_diff_35=0.01996
+  sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_35=1.5727
+  sky130_fd_pr__nfet_01v8_lvt__kt1_diff_35=0.0
+  sky130_fd_pr__nfet_01v8_lvt__voff_diff_35=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b0_diff_35=0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 036, W = 5.05, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8_lvt__kt1_diff_36=0.0
+  sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_36=1.7014
+  sky130_fd_pr__nfet_01v8_lvt__voff_diff_36=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b0_diff_36=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b1_diff_36=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_36=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pclm_diff_36=0.0
+  sky130_fd_pr__nfet_01v8_lvt__keta_diff_36=0.0
+  sky130_fd_pr__nfet_01v8_lvt__k2_diff_36=-0.025254
+  sky130_fd_pr__nfet_01v8_lvt__pdits_diff_36=0.0
+  sky130_fd_pr__nfet_01v8_lvt__eta0_diff_36=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ua_diff_36=-8.2455e-13
+  sky130_fd_pr__nfet_01v8_lvt__ub_diff_36=2.4661e-19
+  sky130_fd_pr__nfet_01v8_lvt__a0_diff_36=0.0
+  sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_36=0.0
+  sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_36=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ags_diff_36=0.0
+  sky130_fd_pr__nfet_01v8_lvt__u0_diff_36=0.0023035
+  sky130_fd_pr__nfet_01v8_lvt__vsat_diff_36=30390.0
+  sky130_fd_pr__nfet_01v8_lvt__vth0_diff_36=0.030922
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 037, W = 5.05, L = 0.25
* -----------------------------------
+  sky130_fd_pr__nfet_01v8_lvt__vth0_diff_37=0.0026675
+  sky130_fd_pr__nfet_01v8_lvt__kt1_diff_37=0.0
+  sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_37=1.43
+  sky130_fd_pr__nfet_01v8_lvt__voff_diff_37=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b0_diff_37=0.0
+  sky130_fd_pr__nfet_01v8_lvt__b1_diff_37=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_37=0.0
+  sky130_fd_pr__nfet_01v8_lvt__pclm_diff_37=0.0
+  sky130_fd_pr__nfet_01v8_lvt__keta_diff_37=0.0
+  sky130_fd_pr__nfet_01v8_lvt__k2_diff_37=-0.00064326
+  sky130_fd_pr__nfet_01v8_lvt__pdits_diff_37=0.0
+  sky130_fd_pr__nfet_01v8_lvt__eta0_diff_37=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ua_diff_37=2.8705e-11
+  sky130_fd_pr__nfet_01v8_lvt__ub_diff_37=-1.9627e-19
+  sky130_fd_pr__nfet_01v8_lvt__a0_diff_37=0.0
+  sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_37=0.0
+  sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_37=0.0
+  sky130_fd_pr__nfet_01v8_lvt__ags_diff_37=0.0
+  sky130_fd_pr__nfet_01v8_lvt__u0_diff_37=-0.005
+  sky130_fd_pr__nfet_01v8_lvt__vsat_diff_37=15849.0
.include "sky130_fd_pr__nfet_01v8_lvt.pm3.spice"
