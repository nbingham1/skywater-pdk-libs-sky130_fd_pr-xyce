* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 68
.param
+  sky130_fd_pr__pfet_01v8_hvt__toxe_mult=0.948
+  sky130_fd_pr__pfet_01v8_hvt__rshp_mult=1.0
+  sky130_fd_pr__pfet_01v8_hvt__overlap_mult=0.91064
+  sky130_fd_pr__pfet_01v8_hvt__lint_diff=1.7325e-8
+  sky130_fd_pr__pfet_01v8_hvt__wint_diff=-3.2175e-8
+  sky130_fd_pr__pfet_01v8_hvt__dlc_diff=1.7325e-8
+  sky130_fd_pr__pfet_01v8_hvt__dwc_diff=-3.2175e-8
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 000, W = 1.26, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_0=0.9411
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_0=-0.067047
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_0=0.00097522
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_0=6.9012e-20
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_0=0.00085309
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_0=-30001.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_0=-0.027673
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_0=-1.6478246e-9
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_0=1.8215e-10
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_0=-0.086124
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 001, W = 1.68, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_1=-0.30543
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_1=0.34808
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_1=-0.069196
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_1=-2.6856e-20
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_1=-0.0068783
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_1=0.00052304
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_1=-20000.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_1=-0.061598
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_1=1.9021e-10
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_1=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 002, W = 1.0, L = 1.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_2=3.9742
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_2=-0.16075
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_2=0.23459
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_2=-0.39733
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_2=1.7862e-19
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_2=-0.0030523
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_2=0.0021714
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_2=0.026641
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_2=6.0283e-10
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_2=2.0425e-10
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 003, W = 1.0, L = 2.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_3=-5.5786e-11
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_3=5.1747
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_3=-0.11369
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_3=0.13176
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_3=-0.42608
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_3=5.1865e-19
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_3=-0.0062951
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_3=0.0020189
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_3=0.036947
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_3=5.4208e-10
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 004, W = 1.0, L = 4.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_4=8.2752e-10
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_4=-6.1212e-11
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_4=6.2965
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_4=-0.12219
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_4=0.14139
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_4=-0.48038
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_4=4.5105e-19
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_4=-0.0087946
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_4=0.0016308
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_4=0.028938
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_4=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 005, W = 1.0, L = 8.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_5=9.6663e-8
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_5=3.4914e-11
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_5=6.8375
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_5=-0.051723
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_5=0.052671
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_5=-0.52626
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_5=4.024e-19
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_5=-0.010302
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_5=0.0021035
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_5=0.025158
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_5=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 006, W = 1.0, L = 0.15
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_6=4.112e-10
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_6=-0.098698
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_6=0.5161
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_6=-0.1228
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_6=-1.3862e-19
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_6=-0.013041
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_6=0.0015101
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_6=-28345.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_6=-0.047639
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 007, W = 1.0, L = 0.18
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_7=0.0010715
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_7=3.3792e-19
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_7=-16338.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_7=-0.058666
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_7=1.0152e-10
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_7=0.070503
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_7=1.2287
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_7=-0.15698
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_7=0.013182
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 008, W = 1.0, L = 0.25
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_8=0.0065099
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_8=0.0021339
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_8=3.4578e-19
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_8=-29942.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_8=0.037342
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_8=2.7913e-9
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_8=4.1649e-10
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_8=1.212
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_8=-0.18101
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 009, W = 1.0, L = 0.5
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_9=-0.32908
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_9=-0.012277
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_9=0.0045307
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_9=4.1908e-20
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_9=-10541.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_9=0.045269
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_9=7.9967e-10
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_9=7.7724e-10
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_9=2.5501
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 010, W = 3.0, L = 1.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_10=7.2706e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_10=-0.38496
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_10=-0.0051457
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_10=0.0060142
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_10=1.8584e-9
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_10=3.6422
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_10=0.0023343
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_10=0.019986
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_10=-0.010112
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_10=-1.437e-10
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 011, W = 3.0, L = 2.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_11=-1.3981e-10
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_11=9.452e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_11=-0.39579
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_11=0.01523
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_11=-0.020292
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_11=1.1978e-9
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_11=5.6703
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_11=0.0035032
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_11=0.013535
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_11=-0.011751
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 012, W = 3.0, L = 4.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_12=-0.010705
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_12=-1.7178e-10
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_12=1.079e-18
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_12=-0.44877
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_12=0.064952
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_12=-0.047067
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_12=8.0408e-10
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_12=6.5488
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_12=0.0041738
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_12=-0.017429
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 013, W = 3.0, L = 8.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_13=6.7444
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_13=0.0048333
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_13=0.0022365
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_13=-0.00843
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_13=-3.3818e-10
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_13=1.4661e-18
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_13=-0.47318
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_13=0.036319
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_13=-0.024161
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_13=1.0307e-10
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_13=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 014, W = 3.0, L = 0.15
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_14=-24769.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_14=0.34296
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_14=0.00040616
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_14=-0.047
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_14=-0.0042041
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_14=9.4745e-11
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_14=4.124e-20
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_14=-0.057777
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_14=-0.085891
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_14=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 015, W = 3.0, L = 0.18
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_15=-6222.8
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_15=1.4602
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_15=0.00089675
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_15=-0.071908
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_15=-8.1586e-5
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_15=1.6305e-10
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_15=1.0152e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_15=0.033077
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_15=-0.16802
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_15=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 016, W = 3.0, L = 0.25
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_16=-28762.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_16=1.3932
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_16=0.0012256
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_16=-0.0016827
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_16=0.0028259
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_16=1.3012e-10
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_16=2.539e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_16=-0.1887
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_16=4.3784e-10
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 017, W = 3.0, L = 0.5
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_17=1.382e-9
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_17=2.9409
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_17=0.0026197
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_17=13860.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_17=0.016554
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_17=-0.006883
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_17=1.1056e-10
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_17=5.0826e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_17=-0.33127
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_17=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 018, W = 5.0, L = 1.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_18=-0.0095271
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_18=0.01149
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_18=3.2771e-9
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_18=3.4979
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_18=0.0023182
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_18=0.016117
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_18=-0.011899
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_18=-1.6357e-10
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_18=7.6564e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_18=-0.35989
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 019, W = 5.0, L = 2.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_19=-0.36951
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_19=0.044883
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_19=-0.024452
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_19=2.107e-9
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_19=5.4335
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_19=0.0031152
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_19=0.0030947
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_19=-0.0081995
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_19=-2.5441e-10
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_19=1.0061e-18
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_19=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 020, W = 5.0, L = 4.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_20=-0.43329
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_20=0.018389
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_20=-0.0096878
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_20=1.2121e-6
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_20=6.4101
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_20=0.0046355
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_20=0.0015876
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_20=-0.0077373
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_20=-3.3629e-10
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_20=1.4023e-18
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 021, W = 5.0, L = 8.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_21=1.3543e-18
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_21=-0.43996
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_21=-0.013374
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_21=0.0048976
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_21=4.5994e-9
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_21=6.3549
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_21=0.0039766
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_21=0.017639
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_21=-0.0066951
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_21=-4.1477e-10
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 022, W = 5.0, L = 0.15
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_22=1.324e-10
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_22=-4.5976e-20
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_22=0.011771
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_22=-0.078894
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_22=-27102.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_22=0.43347
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_22=0.00041692
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_22=-0.069076
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_22=0.00045233
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 023, W = 5.0, L = 0.18
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_23=0.0076182
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_23=1.5074e-10
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_23=7.5942e-20
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_23=0.14242
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_23=-0.15688
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_23=-20000.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_23=1.51
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_23=0.00067272
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_23=-0.05202
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 024, W = 5.0, L = 0.25
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_24=1.4836
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_24=0.00084833
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_24=-0.0077155
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_24=0.001811
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_24=-2.852e-13
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_24=3.5019e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_24=-0.19151
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_24=8.1237e-10
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_24=-11017.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 025, W = 5.0, L = 0.5
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_25=-4202.8
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_25=2.6705
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_25=0.00033419
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_25=0.028862
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_25=-0.0086212
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_25=-1.3033e-11
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_25=1.7081e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_25=-0.29652
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_25=6.3262e-10
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_25=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 026, W = 7.0, L = 1.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_26=3.87
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_26=0.0033127
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_26=0.0066695
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_26=-0.0096254
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_26=-2.915e-10
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_26=1.086e-18
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_26=-0.38966
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_26=0.02118
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_26=-0.014087
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_26=4.7392e-10
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_26=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 027, W = 7.0, L = 2.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_27=5.2996
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_27=0.0045072
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_27=0.0031974
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_27=-0.010442
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_27=-3.7793e-10
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_27=1.4138e-18
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_27=-0.38823
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_27=0.053597
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_27=-0.02939
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_27=1.4678e-10
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 028, W = 7.0, L = 4.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_28=1.0671e-10
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_28=6.2257
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_28=0.0049774
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_28=0.017674
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_28=-0.0066393
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_28=-4.132e-10
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_28=1.5608e-18
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_28=-0.42989
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_28=-0.0077527
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_28=0.0041618
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 029, W = 7.0, L = 8.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_29=-0.0012317
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_29=0.0015529
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_29=5.8812e-10
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_29=6.4717
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_29=0.0092272
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_29=0.0087893
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_29=-0.011014
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_29=-5.3257e-11
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_29=1.8573e-18
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_29=-0.44129
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 030, W = 7.0, L = 0.15
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_30=-0.085522
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_30=-19295.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_30=0.30064
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_30=0.0008238
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_30=-0.070634
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_30=-0.019298
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_30=2.86e-10
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_30=-1.7396e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_30=0.0049521
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_30=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 031, W = 7.0, L = 0.18
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_31=0.15292
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_31=-0.17604
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_31=-3650.6
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_31=1.6642
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_31=0.00025649
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_31=-0.087564
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_31=0.0015551
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_31=-1.6895e-11
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_31=1.885e-19
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 032, W = 7.0, L = 0.25
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_32=2.5238e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_32=-0.19209
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_32=1.118e-9
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_32=-11755.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_32=1.4737
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_32=0.00068642
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_32=-0.003565
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_32=8.2421e-5
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_32=2.8428e-11
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 033, W = 7.0, L = 0.5
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_33=1.9174e-10
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_33=1.8e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_33=-0.33184
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_33=6.5698e-10
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_33=-20000.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_33=3.1038
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_33=0.0021414
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_33=0.0067101
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_33=-0.0091659
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 034, W = 0.42, L = 1.0
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_34=-0.011769
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_34=-1.0721e-10
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_34=1.3365e-18
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_34=-0.4505
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_34=3.0715e-9
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_34=7.9034e-8
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_34=1.0049e-7
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_34=5.6084
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_34=0.0050029
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_34=0.046227
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 035, W = 0.42, L = 20.0
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_35=9.8093
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_35=0.003451
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_35=-0.0087497
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_35=-0.017093
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_35=-1.9758e-10
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_35=9.821e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_35=-0.84741
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_35=-3.9839e-11
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_35=-1.023e-7
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_35=-6.4194e-11
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_35=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 036, W = 0.42, L = 2.0
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_36=5.6513
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_36=0.0062131
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_36=0.013867
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_36=-0.018297
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_36=6.1158e-11
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_36=1.2575e-18
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_36=-0.47411
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_36=3.8354e-10
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_36=5.5002e-8
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_36=8.3075e-10
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 037, W = 0.42, L = 4.0
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_37=2.1173e-9
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_37=6.5595
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_37=0.0031441
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_37=0.033858
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_37=-0.012048
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_37=1.0374e-10
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_37=4.574e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_37=-0.54958
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_37=9.1169e-10
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_37=9.5882e-8
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_37=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 038, W = 0.42, L = 8.0
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_38=4.3623e-8
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_38=-7.1004e-10
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_38=7.1302
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_38=0.0060424
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_38=0.0034632
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_38=-0.016469
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_38=7.736e-10
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_38=3.488e-20
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_38=-0.58662
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_38=4.2361e-10
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 039, W = 0.42, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_39=-4.1396435e-9
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_39=0.4363
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_39=0.0024706
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_39=-51583.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_39=0.050686
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_39=-0.0018016
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_39=5.933e-10
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_39=2.2929e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_39=-0.18611
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_39=-0.13359
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_39=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 040, W = 0.42, L = 0.18
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_40=-2.9262738e-9
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_40=-48473.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_40=-0.20707
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_40=0.0021211
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_40=0.014283
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_40=-0.0085993
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_40=5.5697e-10
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_40=6.3421e-20
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_40=-0.024675
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_40=-0.26698
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_40=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 041, W = 0.42, L = 0.5
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_41=-0.38089
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_41=2.9322e-9
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_41=-38888.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_41=2.8636
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_41=0.0057123
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_41=0.091478
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_41=-0.023719
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_41=4.3063e-10
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_41=8.5174e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_41=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 042, W = 0.55, L = 1.0
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_42=-0.41259
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_42=6.1243e-10
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_42=1.0526e-7
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_42=1.4625e-9
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_42=5.0565
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_42=0.0047
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_42=0.034667
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_42=-0.014806
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_42=7.2762e-10
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_42=-4.3961e-20
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 043, W = 0.55, L = 2.0
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_43=2.8498e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_43=-0.45547
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_43=6.0231e-10
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_43=1.1583e-7
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_43=5.7091e-9
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_43=5.3933
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_43=0.003296
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_43=0.041685
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_43=-0.0061916
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_43=2.8632e-10
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 044, W = 0.55, L = 4.0
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_44=-4.6452e-11
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_44=5.5996e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_44=-0.50649
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_44=7.8525e-10
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_44=9.7149e-8
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_44=1.657e-8
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_44=6.0133
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_44=0.0024625
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_44=0.03279
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_44=-0.0078584
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 045, W = 0.55, L = 8.0
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_45=-0.0088326
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_45=-1.474e-10
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_45=5.7719e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_45=-0.57582
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_45=2.6179e-10
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_45=7.7504e-8
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_45=1.7271e-9
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_45=7.1715
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_45=0.0019517
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_45=0.026282
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 046, W = 0.55, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_46=0.16148
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_46=0.0012053
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_46=-0.037017
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_46=-0.016442
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_46=2.1814e-10
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_46=1.5922e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_46=-0.25251
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_46=-0.033196
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_46=-40000.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 047, W = 0.55, L = 0.5
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_47=-56472.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_47=2.8779
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_47=0.015694
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_47=0.0785
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_47=-0.0080946
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_47=2.0e-9
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_47=1.1367e-18
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_47=-0.35542
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_47=9.3049e-10
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_47=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 048, W = 0.64, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_48=-25394.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_48=0.45527
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_48=0.0011827
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_48=-0.015914
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_48=-0.007354
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_48=2.5998e-10
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_48=1.7343e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_48=-0.18094
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_48=-0.10441
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_48=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 049, W = 0.84, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_49=-31462.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_49=0.4716
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_49=0.0017664
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_49=-0.0070482
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_49=-0.0068842
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_49=5.2165e-10
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_49=-1.2533e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_49=-0.14201
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_49=-0.10472
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_49=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 050, W = 0.64, L = 0.18
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_50=-30815.59945783
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_50=0.00121464
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_50=-0.35079954
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_50=-0.03395799
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_50=0.0010617
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_50=3.46701e-10
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_50=1.396e-20
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_50=-0.18093994
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_50=-0.01214901
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_50=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 051, W = 2.0, L = 0.15
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_51=-14515.01951136
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_51=1.88601e-5
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_51=0.05554018
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_51=-0.07252794
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_51=0.00703588
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_51=5.6917e-11
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_51=-2.9419e-20
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_51=-0.05777702
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_51=-0.044567
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_51=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 052, W = 1.12, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_52=-0.04196204
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_52=-7.6647e-8
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_52=-27284.97988195
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_52=0.0003019
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_52=-0.61499839
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_52=-0.04743662
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_52=0.012422
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_52=6.42999e-11
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_52=1.03621e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_52=-0.09869803
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_52=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 053, W = 1.65, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_53=-0.30542999
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_53=-0.03695201
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_53=-12573.194768
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_53=-0.00054436
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_53=-0.26048985
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_53=-0.07351899
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_53=0.00941368
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_53=-1.5565e-10
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_53=2.02164e-19
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 054, W = 0.84, L = 0.18
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_54=-2.0137e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_54=-0.14201002
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_54=-0.05571701
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_54=-25315.55791728
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_54=0.00157358
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_54=-0.94290034
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_54=-0.05520914
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_54=0.00330583
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_54=5.29585e-10
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 055, W = 1.68, L = 0.18
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_55=1.77615e-10
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_55=-1.065e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_55=0.033077
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_55=-0.11034
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_55=-39146.79616935
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_55=0.00036421
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_55=1.33405999
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_55=-0.0629978
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_55=0.01331141
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 056, W = 0.36, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_56=-0.017396
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_56=8.18463e-10
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_56=-0.00010861
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_56=1.24897e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_56=-0.12438
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_56=0.00033519
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_56=-0.14725461
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_56=0.00237543
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_56=-23579.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_56=-0.01242548
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_56=0.0027449
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_56=-1.1455
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_56=0.056312
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 057, W = 0.54, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_57=0.00036225
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_57=-2.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_57=-0.0060721
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_57=0.00032568
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_57=9.15401e-11
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_57=1.84959e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_57=-0.23683
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_57=-0.09313079
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_57=-0.00011339
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_57=-38643.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_57=0.0005931
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 058, W = 0.63, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_58=-28942.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_58=-0.00042217
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_58=0.0010525
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_58=-1.7696
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_58=-0.026898
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_58=-0.006093
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_58=3.1923e-10
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_58=3.08834e-20
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_58=-0.24292
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_58=0.00018846
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_58=-0.10216024
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_58=7.42226e-5
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_58=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 059, W = 0.7, L = 0.15
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_59=-27201.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_59=0.00143932
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_59=0.0013145
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_59=-2.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_59=-0.034552
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_59=-0.005647
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_59=4.11678e-10
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_59=-6.27298e-20
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_59=-0.19059
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_59=-0.00136297
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_59=-0.087752
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_59=-7.09239e-5
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_59=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 060, W = 0.75, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_60=-7.29796e-5
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_60=-25393.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_60=0.0012886
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_60=0.00148104
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_60=-2.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_60=-0.040648
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_60=-0.0047585
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_60=4.5847e-10
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_60=-1.17829e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_60=-0.14678
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_60=-0.084843
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_60=-0.00140248
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_60=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 061, W = 0.79, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_61=-4.9911e-5
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_61=-23783.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_61=0.00101288
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_61=0.0013326
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_61=-2.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_61=-0.043635
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_61=-0.0044981
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_61=4.91938e-10
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_61=-1.57174e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_61=-0.12427
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_61=-0.086691
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_61=-0.00095916
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_61=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 062, W = 0.82, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_62=-2.22611e-5
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_62=-21900.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_62=0.00045176
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_62=0.0013726
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_62=-2.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_62=-0.046029
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_62=-0.0029267
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_62=5.1504e-10
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_62=-1.84303e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_62=-0.11601
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_62=-0.090668
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_62=-0.0004278
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 063, W = 0.82, L = 0.18
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_63=-0.0004278
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_63=-0.10941523
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_63=-2.22613e-5
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_63=-23535.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_63=0.00045176
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_63=0.0015171
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_63=-1.9097
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_63=-0.026399
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_63=-0.013873
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_63=5.1504e-10
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_63=-1.84303e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_63=0.059877
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_63=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 064, W = 0.82, L = 0.25
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_64=0.31938
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_64=-434810.89830208
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_64=-0.00046359
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_64=0.00047433
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_64=-0.2004
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_64=3.46622e-5
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_64=-19223.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_64=0.0022188
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_64=2.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_64=0.011884
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_64=0.0049685
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_64=2.61701e-10
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_64=3.89042e-19
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 065, W = 0.82, L = 0.5
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_65=0.042562
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_65=-0.5
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_65=-15187.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_65=-0.00058999
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_65=1.4213
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_65=0.042493
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_65=-0.0016053
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_65=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 066, W = 0.86, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_66=4.61965e-10
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_66=-1.56897e-19
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_66=-0.13882
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_66=0.00031999
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_66=-0.10432908
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_66=1.91787e-6
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_66=-18965.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_66=2.59995e-5
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_66=0.0012435
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_66=-2.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_66=-0.054565
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_66=-0.0024326
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 067, W = 0.94, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_67=-0.0012624
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_67=2.20238e-10
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_67=1.67256e-21
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_67=-0.12553
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_67=0.00057533
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_67=-0.08465745
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_67=3.44709e-6
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_67=-17711.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_67=4.67463e-5
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_67=0.00053342
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_67=-1.6708
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_67=-0.038792
.include "sky130_fd_pr__pfet_01v8_hvt.pm3.spice"
