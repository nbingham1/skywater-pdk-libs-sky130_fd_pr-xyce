* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 11
.param
+  sky130_fd_pr__esd_nfet_g5v0d10v5__toxe_mult=1.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__rshn_mult=1.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__overlap_mult=0.89805
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ajunction_mult=9.9505e-1
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pjunction_mult=1.0144e+0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__lint_diff=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__wint_diff=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__dlc_diff=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__dwc_diff=0.0
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 000, W = 17.5, L = 0.55
* -----------------------------------
+  sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_0=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_0=0.23362
+  sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_0=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_0=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_0=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_0=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_0=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_0=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_0=0.010406
+  sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_0=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_0=0.001245
+  sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_0=0.012769
+  sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_0=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_0=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_0=-1672.2
+  sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_0=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_0=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_0=2.4153e-19
+  sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_0=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_0=-8.8395e-12
+  sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_0=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_0=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_0=0.0
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 001, W = 19.5, L = 0.55
* -----------------------------------
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_1=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_1=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_1=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_1=0.23014
+  sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_1=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_1=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_1=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_1=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_1=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_1=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_1=0.010327
+  sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_1=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_1=0.0029959
+  sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_1=0.014049
+  sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_1=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_1=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_1=-1443.7
+  sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_1=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_1=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_1=3.4221e-19
+  sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_1=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_1=-2.42e-11
+  sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_1=0.0
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 002, W = 21.5, L = 0.55
* -----------------------------------
+  sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_2=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_2=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_2=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_2=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_2=0.23391
+  sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_2=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_2=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_2=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_2=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_2=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_2=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_2=0.010304
+  sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_2=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_2=0.0012741
+  sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_2=0.013326
+  sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_2=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_2=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_2=-43.451
+  sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_2=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_2=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_2=3.291e-19
+  sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_2=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_2=-7.333e-12
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 003, W = 23.5, L = 0.55
* -----------------------------------
+  sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_3=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_3=-1.7201e-12
+  sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_3=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_3=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_3=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_3=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_3=0.23086
+  sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_3=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_3=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_3=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_3=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_3=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_3=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_3=0.010034
+  sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_3=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_3=0.0010628
+  sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_3=0.01319
+  sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_3=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_3=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_3=33.54
+  sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_3=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_3=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_3=3.183e-19
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 004, W = 26.5, L = 0.55
* -----------------------------------
+  sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_4=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_4=2.7249e-19
+  sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_4=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_4=-7.6527e-12
+  sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_4=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_4=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_4=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_4=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_4=0.22609
+  sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_4=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_4=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_4=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_4=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_4=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_4=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_4=0.0099796
+  sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_4=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_4=0.0013927
+  sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_4=0.011469
+  sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_4=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_4=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_4=-907.07
+  sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_4=0.0
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 005, W = 30.25, L = 1.0
* -----------------------------------
+  sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_5=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_5=-6.1783e-19
+  sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_5=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_5=8.2128e-11
+  sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_5=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_5=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_5=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_5=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_5=0.27056
+  sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_5=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_5=-0.021325
+  sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_5=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_5=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_5=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_5=-0.26694
+  sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_5=0.047533
+  sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_5=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_5=-0.0063931
+  sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_5=0.010431
+  sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_5=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_5=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_5=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_5=0.0
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 006, W = 30.25, L = 0.55
* ------------------------------------
+  sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_6=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_6=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_6=6.0666e-19
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_6=-7.0128e-12
+  sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_6=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_6=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_6=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_6=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_6=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_6=0.22669
+  sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_6=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_6=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_6=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_6=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_6=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_6=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_6=0.010019
+  sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_6=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_6=0.0016874
+  sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_6=0.011396
+  sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_6=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_6=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_6=1500.0
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 007, W = 40.31, L = 0.55
* ------------------------------------
+  sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_7=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_7=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_7=3019.2
+  sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_7=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_7=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_7=9.7977e-19
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_7=3.2228e-12
+  sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_7=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_7=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_7=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_7=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_7=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_7=0.19932
+  sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_7=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_7=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_7=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_7=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_7=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_7=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_7=0.010207
+  sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_7=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_7=0.0014468
+  sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_7=0.011899
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 008, W = 50.99, L = 1.0
* -----------------------------------
+  sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_8=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_8=-0.0088519
+  sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_8=-8.0124e-5
+  sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_8=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_8=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_8=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_8=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_8=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_8=-6.7671e-19
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_8=5.5348e-11
+  sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_8=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_8=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_8=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_8=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_8=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_8=0.25888
+  sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_8=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_8=0.0071088
+  sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_8=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_8=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_8=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_8=0.0024548
+  sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_8=0.010977
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 009, W = 50.99, L = 0.55
* ------------------------------------
+  sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_9=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_9=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_9=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_9=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_9=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_9=0.0014488
+  sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_9=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_9=0.0037985
+  sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_9=0.002943
+  sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_9=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_9=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_9=-191.5
+  sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_9=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_9=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_9=1.3051e-18
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_9=-1.3283e-11
+  sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_9=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_9=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_9=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_9=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_9=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_9=0.20721
+  sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_9=0.0
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 010, W = 5.4, L = 0.6
* ---------------------------------
+  sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_10=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_10=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_10=2.8803e-12
+  sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_10=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_10=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_10=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_10=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_10=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_10=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_10=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_10=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_10=-2502.2
+  sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_10=8.2506e-20
+  sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_10=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_10=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_10=0.0031768
+  sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_10=0.29591
+  sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_10=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_10=-0.00045045
+  sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_10=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_10=0.013543
+  sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_10=0.0
+  sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_10=0.0
.include "sky130_fd_pr__esd_nfet_g5v0d10v5.pm3.spice"
