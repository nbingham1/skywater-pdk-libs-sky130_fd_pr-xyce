* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 63
.param
+  sky130_fd_pr__nfet_01v8__toxe_mult=1.0
+  sky130_fd_pr__nfet_01v8__rshn_mult=1.0
+  sky130_fd_pr__nfet_01v8__overlap_mult=0.9642
+  sky130_fd_pr__nfet_01v8__lint_diff=0.0
+  sky130_fd_pr__nfet_01v8__wint_diff=0.0
+  sky130_fd_pr__nfet_01v8__dlc_diff=-.61491e-9
+  sky130_fd_pr__nfet_01v8__dwc_diff=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 000, W = 1.26, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__voff_diff_0=-0.064628
+  sky130_fd_pr__nfet_01v8__kt1_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_0=-1.1675e-19
+  sky130_fd_pr__nfet_01v8__pditsd_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_0=1.3935e-11
+  sky130_fd_pr__nfet_01v8__vsat_diff_0=2157.4
+  sky130_fd_pr__nfet_01v8__tvoff_diff_0=-0.0010664
+  sky130_fd_pr__nfet_01v8__ags_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_0=0.0013235
+  sky130_fd_pr__nfet_01v8__vth0_diff_0=-0.018052
+  sky130_fd_pr__nfet_01v8__nfactor_diff_0=0.5869
+  sky130_fd_pr__nfet_01v8__u0_diff_0=-0.0032648
+  sky130_fd_pr__nfet_01v8__eta0_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_0=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 001, W = 1.68, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__eta0_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_1=-0.062332
+  sky130_fd_pr__nfet_01v8__kt1_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_1=-1.6979e-19
+  sky130_fd_pr__nfet_01v8__pditsd_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_1=1.0381e-11
+  sky130_fd_pr__nfet_01v8__vsat_diff_1=1545.5
+  sky130_fd_pr__nfet_01v8__tvoff_diff_1=-0.0010597
+  sky130_fd_pr__nfet_01v8__ags_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_1=0.0030943
+  sky130_fd_pr__nfet_01v8__vth0_diff_1=0.012094
+  sky130_fd_pr__nfet_01v8__nfactor_diff_1=0.4994
+  sky130_fd_pr__nfet_01v8__u0_diff_1=-0.0025003
*
* sky130_fd_pr__nfet_01v8, Bin 002, W = 1.0, L = 1.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__nfactor_diff_2=0.79822
+  sky130_fd_pr__nfet_01v8__u0_diff_2=-1.4501e-5
+  sky130_fd_pr__nfet_01v8__vth0_diff_2=0.0093572
+  sky130_fd_pr__nfet_01v8__eta0_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_2=-0.097681
+  sky130_fd_pr__nfet_01v8__ub_diff_2=1.6548e-19
+  sky130_fd_pr__nfet_01v8__kt1_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_2=4.5462e-13
+  sky130_fd_pr__nfet_01v8__vsat_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_2=-0.0011898
+  sky130_fd_pr__nfet_01v8__ags_diff_2=-0.046289
+  sky130_fd_pr__nfet_01v8__a0_diff_2=0.20611
+  sky130_fd_pr__nfet_01v8__b0_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_2=-0.00724
*
* sky130_fd_pr__nfet_01v8, Bin 003, W = 1.0, L = 2.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__keta_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_3=-0.0072176
+  sky130_fd_pr__nfet_01v8__nfactor_diff_3=0.6874
+  sky130_fd_pr__nfet_01v8__u0_diff_3=-0.00018122
+  sky130_fd_pr__nfet_01v8__vth0_diff_3=0.0070337
+  sky130_fd_pr__nfet_01v8__eta0_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_3=-0.10233
+  sky130_fd_pr__nfet_01v8__ub_diff_3=9.8355e-20
+  sky130_fd_pr__nfet_01v8__kt1_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_3=5.2286e-13
+  sky130_fd_pr__nfet_01v8__vsat_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_3=-0.00088509
+  sky130_fd_pr__nfet_01v8__ags_diff_3=0.0089251
+  sky130_fd_pr__nfet_01v8__a0_diff_3=-0.0090083
+  sky130_fd_pr__nfet_01v8__b0_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_3=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 004, W = 1.0, L = 4.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__pdits_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_4=-0.0010891
+  sky130_fd_pr__nfet_01v8__nfactor_diff_4=0.78898
+  sky130_fd_pr__nfet_01v8__u0_diff_4=-0.0011684
+  sky130_fd_pr__nfet_01v8__vth0_diff_4=0.012209
+  sky130_fd_pr__nfet_01v8__eta0_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_4=-0.11872
+  sky130_fd_pr__nfet_01v8__ub_diff_4=-1.6247e-20
+  sky130_fd_pr__nfet_01v8__kt1_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_4=4.1897e-12
+  sky130_fd_pr__nfet_01v8__vsat_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_4=-0.00046714
+  sky130_fd_pr__nfet_01v8__ags_diff_4=0.017325
+  sky130_fd_pr__nfet_01v8__a0_diff_4=-0.021601
+  sky130_fd_pr__nfet_01v8__b0_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_4=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 005, W = 1.0, L = 8.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__pdits_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_5=0.0019485
+  sky130_fd_pr__nfet_01v8__nfactor_diff_5=0.81593
+  sky130_fd_pr__nfet_01v8__u0_diff_5=-0.0016431
+  sky130_fd_pr__nfet_01v8__vth0_diff_5=0.0075363
+  sky130_fd_pr__nfet_01v8__eta0_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_5=-0.1266
+  sky130_fd_pr__nfet_01v8__ub_diff_5=-2.1979e-20
+  sky130_fd_pr__nfet_01v8__kt1_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_5=5.0336e-12
+  sky130_fd_pr__nfet_01v8__vsat_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_5=0.00014598
+  sky130_fd_pr__nfet_01v8__ags_diff_5=0.0023677
+  sky130_fd_pr__nfet_01v8__a0_diff_5=0.0023303
+  sky130_fd_pr__nfet_01v8__b0_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_5=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 006, W = 1.0, L = 0.15
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__pclm_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_6=-0.0013648
+  sky130_fd_pr__nfet_01v8__nfactor_diff_6=0.60969
+  sky130_fd_pr__nfet_01v8__u0_diff_6=-0.0036763
+  sky130_fd_pr__nfet_01v8__vth0_diff_6=0.0053925
+  sky130_fd_pr__nfet_01v8__eta0_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_6=-0.07115
+  sky130_fd_pr__nfet_01v8__ub_diff_6=-3.443e-19
+  sky130_fd_pr__nfet_01v8__kt1_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_6=1.4919e-11
+  sky130_fd_pr__nfet_01v8__vsat_diff_6=-723.7
+  sky130_fd_pr__nfet_01v8__tvoff_diff_6=-0.0010051
+  sky130_fd_pr__nfet_01v8__ags_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_6=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 007, W = 1.0, L = 0.18
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__tvoff_diff_7=-0.0018088
+  sky130_fd_pr__nfet_01v8__b0_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_7=0.0020165
+  sky130_fd_pr__nfet_01v8__nfactor_diff_7=0.71326
+  sky130_fd_pr__nfet_01v8__u0_diff_7=-0.0036247
+  sky130_fd_pr__nfet_01v8__vth0_diff_7=-0.0087946
+  sky130_fd_pr__nfet_01v8__eta0_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_7=-0.072216
+  sky130_fd_pr__nfet_01v8__ub_diff_7=-2.5113e-19
+  sky130_fd_pr__nfet_01v8__kt1_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_7=1.4741e-11
+  sky130_fd_pr__nfet_01v8__vsat_diff_7=-4205.9
+  sky130_fd_pr__nfet_01v8__a0_diff_7=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 008, W = 1.0, L = 0.25
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__a0_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_8=1.9388e-11
+  sky130_fd_pr__nfet_01v8__tvoff_diff_8=-0.0017778
+  sky130_fd_pr__nfet_01v8__b0_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_8=-0.00090345
+  sky130_fd_pr__nfet_01v8__nfactor_diff_8=0.85238
+  sky130_fd_pr__nfet_01v8__u0_diff_8=-0.0050754
+  sky130_fd_pr__nfet_01v8__vth0_diff_8=-0.0056636
+  sky130_fd_pr__nfet_01v8__eta0_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_8=-0.085488
+  sky130_fd_pr__nfet_01v8__ub_diff_8=-7.5909e-20
+  sky130_fd_pr__nfet_01v8__kt1_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_8=-12323.0
*
* sky130_fd_pr__nfet_01v8, Bin 009, W = 1.0, L = 0.5
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__kt1_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_9=-1.1801e-19
+  sky130_fd_pr__nfet_01v8__vsat_diff_9=-3282.1
+  sky130_fd_pr__nfet_01v8__a0_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_9=6.0594e-12
+  sky130_fd_pr__nfet_01v8__tvoff_diff_9=-0.0011855
+  sky130_fd_pr__nfet_01v8__b0_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_9=0.0016142
+  sky130_fd_pr__nfet_01v8__nfactor_diff_9=0.71331
+  sky130_fd_pr__nfet_01v8__u0_diff_9=-0.0023313
+  sky130_fd_pr__nfet_01v8__vth0_diff_9=0.012758
+  sky130_fd_pr__nfet_01v8__eta0_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_9=-0.09488
*
* sky130_fd_pr__nfet_01v8, Bin 010, W = 2.0, L = 0.15
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__ags_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_10=0.0017497
+  sky130_fd_pr__nfet_01v8__ua_diff_10=6.5387e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_10=-1.6773e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_10=-0.0014711
+  sky130_fd_pr__nfet_01v8__a0_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_10=-1965.1
+  sky130_fd_pr__nfet_01v8__kt1_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_10=0.010515
+  sky130_fd_pr__nfet_01v8__pdits_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_10=-0.055251
+  sky130_fd_pr__nfet_01v8__b1_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_10=0.44391
+  sky130_fd_pr__nfet_01v8__u0_diff_10=-0.0015785
*
* sky130_fd_pr__nfet_01v8, Bin 011, W = 3.0, L = 1.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__pclm_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_11=0.54938
+  sky130_fd_pr__nfet_01v8__u0_diff_11=-0.00010243
+  sky130_fd_pr__nfet_01v8__ags_diff_11=0.032488
+  sky130_fd_pr__nfet_01v8__keta_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_11=-0.0047234
+  sky130_fd_pr__nfet_01v8__ua_diff_11=3.5948e-14
+  sky130_fd_pr__nfet_01v8__eta0_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_11=6.1194e-20
+  sky130_fd_pr__nfet_01v8__tvoff_diff_11=-0.0016212
+  sky130_fd_pr__nfet_01v8__a0_diff_11=0.0087374
+  sky130_fd_pr__nfet_01v8__rdsw_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_11=0.012888
+  sky130_fd_pr__nfet_01v8__pdits_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_11=-0.077584
+  sky130_fd_pr__nfet_01v8__b1_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_11=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 012, W = 3.0, L = 2.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__pditsd_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_12=0.63836
+  sky130_fd_pr__nfet_01v8__u0_diff_12=-0.0024136
+  sky130_fd_pr__nfet_01v8__ags_diff_12=0.022869
+  sky130_fd_pr__nfet_01v8__keta_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_12=-0.0028244
+  sky130_fd_pr__nfet_01v8__ua_diff_12=8.1792e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_12=-2.2603e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_12=-0.0018063
+  sky130_fd_pr__nfet_01v8__a0_diff_12=-0.014898
+  sky130_fd_pr__nfet_01v8__rdsw_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_12=0.013207
+  sky130_fd_pr__nfet_01v8__pdits_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_12=-0.089272
+  sky130_fd_pr__nfet_01v8__b1_diff_12=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 013, W = 3.0, L = 4.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__pdits_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_13=-0.098313
+  sky130_fd_pr__nfet_01v8__b1_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_13=0.66392
+  sky130_fd_pr__nfet_01v8__u0_diff_13=-0.0024877
+  sky130_fd_pr__nfet_01v8__ags_diff_13=0.030763
+  sky130_fd_pr__nfet_01v8__keta_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_13=-0.0023283
+  sky130_fd_pr__nfet_01v8__ua_diff_13=8.1683e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_13=-2.1077e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_13=-0.0012463
+  sky130_fd_pr__nfet_01v8__a0_diff_13=-0.040181
+  sky130_fd_pr__nfet_01v8__rdsw_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_13=0.013899
+  sky130_fd_pr__nfet_01v8__b0_diff_13=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 014, W = 3.0, L = 8.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__b0_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_14=-0.10972
+  sky130_fd_pr__nfet_01v8__b1_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_14=0.71135
+  sky130_fd_pr__nfet_01v8__u0_diff_14=-0.0018386
+  sky130_fd_pr__nfet_01v8__ags_diff_14=0.0025727
+  sky130_fd_pr__nfet_01v8__keta_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_14=-0.00010451
+  sky130_fd_pr__nfet_01v8__ua_diff_14=5.8682e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_14=-1.7238e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_14=-0.00052901
+  sky130_fd_pr__nfet_01v8__a0_diff_14=0.0015089
+  sky130_fd_pr__nfet_01v8__rdsw_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_14=0.010809
*
* sky130_fd_pr__nfet_01v8, Bin 015, W = 3.0, L = 0.15
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__kt1_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_15=2927.1
+  sky130_fd_pr__nfet_01v8__vth0_diff_15=-0.0010819
+  sky130_fd_pr__nfet_01v8__b0_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_15=-0.059619
+  sky130_fd_pr__nfet_01v8__b1_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_15=0.49831
+  sky130_fd_pr__nfet_01v8__u0_diff_15=-0.0033038
+  sky130_fd_pr__nfet_01v8__ags_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_15=0.0047759
+  sky130_fd_pr__nfet_01v8__ua_diff_15=1.3818e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_15=-3.6525e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_15=-0.0016275
+  sky130_fd_pr__nfet_01v8__a0_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_15=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 016, W = 3.0, L = 0.18
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__a0_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_16=435.25
+  sky130_fd_pr__nfet_01v8__vth0_diff_16=0.0053171
+  sky130_fd_pr__nfet_01v8__b0_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_16=-0.082621
+  sky130_fd_pr__nfet_01v8__b1_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_16=0.6968
+  sky130_fd_pr__nfet_01v8__u0_diff_16=-0.0016247
+  sky130_fd_pr__nfet_01v8__ags_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_16=0.0072238
+  sky130_fd_pr__nfet_01v8__ua_diff_16=7.4303e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_16=-3.9342e-20
+  sky130_fd_pr__nfet_01v8__tvoff_diff_16=-0.0015057
*
* sky130_fd_pr__nfet_01v8, Bin 017, W = 3.0, L = 0.25
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__tvoff_diff_17=-0.001088
+  sky130_fd_pr__nfet_01v8__a0_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_17=1659.5
+  sky130_fd_pr__nfet_01v8__vth0_diff_17=0.00057154
+  sky130_fd_pr__nfet_01v8__pdits_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_17=-0.10595
+  sky130_fd_pr__nfet_01v8__b0_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_17=0.86746
+  sky130_fd_pr__nfet_01v8__u0_diff_17=-0.00095171
+  sky130_fd_pr__nfet_01v8__ags_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_17=0.0026444
+  sky130_fd_pr__nfet_01v8__ua_diff_17=3.3377e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_17=8.1803e-20
*
* sky130_fd_pr__nfet_01v8, Bin 018, W = 3.0, L = 0.5
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__ub_diff_18=5.989e-20
+  sky130_fd_pr__nfet_01v8__tvoff_diff_18=-0.0016726
+  sky130_fd_pr__nfet_01v8__a0_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_18=5980.5
+  sky130_fd_pr__nfet_01v8__vth0_diff_18=0.0026655
+  sky130_fd_pr__nfet_01v8__pdits_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_18=-0.08199
+  sky130_fd_pr__nfet_01v8__b0_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_18=0.61703
+  sky130_fd_pr__nfet_01v8__u0_diff_18=-0.00076014
+  sky130_fd_pr__nfet_01v8__ags_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_18=0.00035836
+  sky130_fd_pr__nfet_01v8__ua_diff_18=2.2684e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_18=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 019, W = 5.0, L = 1.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__eta0_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_19=4.4209e-13
+  sky130_fd_pr__nfet_01v8__ub_diff_19=8.0805e-20
+  sky130_fd_pr__nfet_01v8__tvoff_diff_19=-0.002134
+  sky130_fd_pr__nfet_01v8__a0_diff_19=0.023621
+  sky130_fd_pr__nfet_01v8__rdsw_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_19=0.013467
+  sky130_fd_pr__nfet_01v8__pdits_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_19=-0.063774
+  sky130_fd_pr__nfet_01v8__b0_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_19=0.51452
+  sky130_fd_pr__nfet_01v8__u0_diff_19=-2.2775e-5
+  sky130_fd_pr__nfet_01v8__ags_diff_19=0.071639
+  sky130_fd_pr__nfet_01v8__keta_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_19=0.0026875
*
* sky130_fd_pr__nfet_01v8, Bin 020, W = 5.0, L = 2.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__ua_diff_20=1.2021e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_20=-3.4149e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_20=-0.0033097
+  sky130_fd_pr__nfet_01v8__a0_diff_20=-0.058498
+  sky130_fd_pr__nfet_01v8__rdsw_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_20=0.011105
+  sky130_fd_pr__nfet_01v8__pdits_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_20=-0.065636
+  sky130_fd_pr__nfet_01v8__b1_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_20=0.50805
+  sky130_fd_pr__nfet_01v8__u0_diff_20=-0.0035071
+  sky130_fd_pr__nfet_01v8__ags_diff_20=0.043441
+  sky130_fd_pr__nfet_01v8__keta_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_20=-0.0027139
*
* sky130_fd_pr__nfet_01v8, Bin 021, W = 5.0, L = 4.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__ags_diff_21=-0.013061
+  sky130_fd_pr__nfet_01v8__keta_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_21=-0.0019562
+  sky130_fd_pr__nfet_01v8__ua_diff_21=7.4952e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_21=-2.4257e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_21=-0.0014564
+  sky130_fd_pr__nfet_01v8__a0_diff_21=0.014722
+  sky130_fd_pr__nfet_01v8__rdsw_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_21=0.009246
+  sky130_fd_pr__nfet_01v8__pdits_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_21=-0.088517
+  sky130_fd_pr__nfet_01v8__b1_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_21=0.6428
+  sky130_fd_pr__nfet_01v8__u0_diff_21=-0.0022
*
* sky130_fd_pr__nfet_01v8, Bin 022, W = 5.0, L = 8.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__pclm_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_22=0.63922
+  sky130_fd_pr__nfet_01v8__u0_diff_22=-0.0010696
+  sky130_fd_pr__nfet_01v8__ags_diff_22=0.034141
+  sky130_fd_pr__nfet_01v8__keta_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_22=0.00030352
+  sky130_fd_pr__nfet_01v8__ua_diff_22=4.0804e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_22=-8.907e-20
+  sky130_fd_pr__nfet_01v8__tvoff_diff_22=-0.00092569
+  sky130_fd_pr__nfet_01v8__a0_diff_22=-0.032971
+  sky130_fd_pr__nfet_01v8__rdsw_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_22=0.015113
+  sky130_fd_pr__nfet_01v8__pdits_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_22=-0.10034
+  sky130_fd_pr__nfet_01v8__b1_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_22=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 023, W = 5.0, L = 0.15
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__pditsd_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_23=0.575
+  sky130_fd_pr__nfet_01v8__u0_diff_23=0.00044492
+  sky130_fd_pr__nfet_01v8__ags_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_23=-0.0027994
+  sky130_fd_pr__nfet_01v8__ua_diff_23=-6.8599e-13
+  sky130_fd_pr__nfet_01v8__eta0_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_23=5.4464e-20
+  sky130_fd_pr__nfet_01v8__tvoff_diff_23=-0.0018474
+  sky130_fd_pr__nfet_01v8__a0_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_23=9075.1
+  sky130_fd_pr__nfet_01v8__kt1_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_23=0.019052
+  sky130_fd_pr__nfet_01v8__pdits_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_23=-0.045722
+  sky130_fd_pr__nfet_01v8__b1_diff_23=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 024, W = 5.0, L = 0.18
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__pdits_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_24=-0.08713
+  sky130_fd_pr__nfet_01v8__b1_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_24=0.74684
+  sky130_fd_pr__nfet_01v8__u0_diff_24=-0.0062104
+  sky130_fd_pr__nfet_01v8__ags_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_24=-0.00046357
+  sky130_fd_pr__nfet_01v8__ua_diff_24=2.5229e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_24=-4.484e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_24=-0.0016383
+  sky130_fd_pr__nfet_01v8__a0_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_24=4959.2
+  sky130_fd_pr__nfet_01v8__kt1_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_24=0.011679
+  sky130_fd_pr__nfet_01v8__b0_diff_24=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 025, W = 5.0, L = 0.25
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__b0_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_25=-0.093762
+  sky130_fd_pr__nfet_01v8__b1_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_25=0.75331
+  sky130_fd_pr__nfet_01v8__u0_diff_25=-0.0006673
+  sky130_fd_pr__nfet_01v8__ags_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_25=0.0012241
+  sky130_fd_pr__nfet_01v8__ua_diff_25=2.7261e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_25=1.3675e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_25=-0.001606
+  sky130_fd_pr__nfet_01v8__a0_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_25=551.45
+  sky130_fd_pr__nfet_01v8__kt1_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_25=0.015315
*
* sky130_fd_pr__nfet_01v8, Bin 026, W = 5.0, L = 0.5
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__kt1_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_26=97.678
+  sky130_fd_pr__nfet_01v8__vth0_diff_26=0.0071389
+  sky130_fd_pr__nfet_01v8__b0_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_26=-0.078497
+  sky130_fd_pr__nfet_01v8__b1_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_26=0.59452
+  sky130_fd_pr__nfet_01v8__u0_diff_26=-5.6453e-5
+  sky130_fd_pr__nfet_01v8__ags_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_26=-0.00055127
+  sky130_fd_pr__nfet_01v8__ua_diff_26=-1.4727e-13
+  sky130_fd_pr__nfet_01v8__eta0_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_26=3.1599e-20
+  sky130_fd_pr__nfet_01v8__tvoff_diff_26=-0.001874
+  sky130_fd_pr__nfet_01v8__a0_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_26=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 027, W = 7.0, L = 1.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__a0_diff_27=-0.0096151
+  sky130_fd_pr__nfet_01v8__rdsw_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_27=4.6847e-5
+  sky130_fd_pr__nfet_01v8__b0_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_27=-0.053961
+  sky130_fd_pr__nfet_01v8__b1_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_27=0.42737
+  sky130_fd_pr__nfet_01v8__u0_diff_27=-0.0010941
+  sky130_fd_pr__nfet_01v8__ags_diff_27=0.01028
+  sky130_fd_pr__nfet_01v8__keta_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_27=-6.4543e-6
+  sky130_fd_pr__nfet_01v8__ua_diff_27=4.6745e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_27=-1.0031e-20
+  sky130_fd_pr__nfet_01v8__tvoff_diff_27=-0.0030825
*
* sky130_fd_pr__nfet_01v8, Bin 028, W = 7.0, L = 2.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__tvoff_diff_28=-0.0032098
+  sky130_fd_pr__nfet_01v8__a0_diff_28=-0.033895
+  sky130_fd_pr__nfet_01v8__rdsw_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_28=0.015331
+  sky130_fd_pr__nfet_01v8__pdits_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_28=-0.062388
+  sky130_fd_pr__nfet_01v8__b0_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_28=0.5083
+  sky130_fd_pr__nfet_01v8__u0_diff_28=-0.0010506
+  sky130_fd_pr__nfet_01v8__ags_diff_28=0.033476
+  sky130_fd_pr__nfet_01v8__keta_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_28=-0.0012416
+  sky130_fd_pr__nfet_01v8__ua_diff_28=4.7856e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_28=-7.3548e-20
*
* sky130_fd_pr__nfet_01v8, Bin 029, W = 7.0, L = 4.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__ub_diff_29=-4.1864e-20
+  sky130_fd_pr__nfet_01v8__tvoff_diff_29=-0.0025932
+  sky130_fd_pr__nfet_01v8__a0_diff_29=-0.075736
+  sky130_fd_pr__nfet_01v8__rdsw_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_29=0.010933
+  sky130_fd_pr__nfet_01v8__pdits_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_29=-0.070195
+  sky130_fd_pr__nfet_01v8__b0_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_29=0.52113
+  sky130_fd_pr__nfet_01v8__u0_diff_29=-0.00077386
+  sky130_fd_pr__nfet_01v8__ags_diff_29=0.056699
+  sky130_fd_pr__nfet_01v8__keta_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_29=-0.002407
+  sky130_fd_pr__nfet_01v8__ua_diff_29=3.7953e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_29=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 030, W = 7.0, L = 8.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__eta0_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_30=-6.3508e-20
+  sky130_fd_pr__nfet_01v8__tvoff_diff_30=-0.0020233
+  sky130_fd_pr__nfet_01v8__a0_diff_30=-0.022257
+  sky130_fd_pr__nfet_01v8__rdsw_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_30=0.014677
+  sky130_fd_pr__nfet_01v8__pdits_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_30=-0.076178
+  sky130_fd_pr__nfet_01v8__b1_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_30=0.50474
+  sky130_fd_pr__nfet_01v8__u0_diff_30=-0.00064091
+  sky130_fd_pr__nfet_01v8__ags_diff_30=0.025094
+  sky130_fd_pr__nfet_01v8__keta_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_30=0.00013166
+  sky130_fd_pr__nfet_01v8__ua_diff_30=2.9064e-12
*
* sky130_fd_pr__nfet_01v8, Bin 031, W = 7.0, L = 0.15
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__ua_diff_31=-6.1562e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_31=2.6424e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_31=-0.0015564
+  sky130_fd_pr__nfet_01v8__a0_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_31=6449.4
+  sky130_fd_pr__nfet_01v8__kt1_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_31=0.0077181
+  sky130_fd_pr__nfet_01v8__pdits_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_31=-0.040033
+  sky130_fd_pr__nfet_01v8__b1_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_31=0.32942
+  sky130_fd_pr__nfet_01v8__u0_diff_31=0.0021463
+  sky130_fd_pr__nfet_01v8__ags_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_31=-0.0028519
*
* sky130_fd_pr__nfet_01v8, Bin 032, W = 7.0, L = 0.18
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__ags_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_32=-0.00047936
+  sky130_fd_pr__nfet_01v8__ua_diff_32=2.0407e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_32=-3.0535e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_32=-0.00099185
+  sky130_fd_pr__nfet_01v8__a0_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_32=5345.4
+  sky130_fd_pr__nfet_01v8__kt1_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_32=0.0068981
+  sky130_fd_pr__nfet_01v8__pdits_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_32=-0.097013
+  sky130_fd_pr__nfet_01v8__b1_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_32=0.834
+  sky130_fd_pr__nfet_01v8__u0_diff_32=-0.0048436
*
* sky130_fd_pr__nfet_01v8, Bin 033, W = 7.0, L = 0.25
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__pclm_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_33=0.60689
+  sky130_fd_pr__nfet_01v8__u0_diff_33=-0.00085323
+  sky130_fd_pr__nfet_01v8__ags_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_33=0.0021179
+  sky130_fd_pr__nfet_01v8__ua_diff_33=3.6045e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_33=9.6789e-20
+  sky130_fd_pr__nfet_01v8__tvoff_diff_33=-0.0026528
+  sky130_fd_pr__nfet_01v8__a0_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_33=43.864
+  sky130_fd_pr__nfet_01v8__kt1_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_33=0.011424
+  sky130_fd_pr__nfet_01v8__pdits_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_33=-0.07207
+  sky130_fd_pr__nfet_01v8__b1_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_33=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 034, W = 7.0, L = 0.5
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__pditsd_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_34=0.48132
+  sky130_fd_pr__nfet_01v8__u0_diff_34=-3.0443e-5
+  sky130_fd_pr__nfet_01v8__ags_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_34=-0.001448
+  sky130_fd_pr__nfet_01v8__ua_diff_34=3.6306e-15
+  sky130_fd_pr__nfet_01v8__eta0_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_34=2.1029e-20
+  sky130_fd_pr__nfet_01v8__tvoff_diff_34=-0.0025929
+  sky130_fd_pr__nfet_01v8__a0_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_34=1751.1
+  sky130_fd_pr__nfet_01v8__kt1_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_34=0.0062944
+  sky130_fd_pr__nfet_01v8__pdits_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_34=-0.06035
+  sky130_fd_pr__nfet_01v8__b1_diff_34=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 035, W = 0.42, L = 1.0
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__pdits_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_35=-0.086838
+  sky130_fd_pr__nfet_01v8__b1_diff_35=1.326e-8
+  sky130_fd_pr__nfet_01v8__pditsd_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_35=0.64226
+  sky130_fd_pr__nfet_01v8__u0_diff_35=-0.0046136
+  sky130_fd_pr__nfet_01v8__ags_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_35=-0.0045356
+  sky130_fd_pr__nfet_01v8__ua_diff_35=1.4292e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_35=-1.067e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_35=-0.0018951
+  sky130_fd_pr__nfet_01v8__a0_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_35=0.0095294
+  sky130_fd_pr__nfet_01v8__b0_diff_35=-1.7482e-7
*
* sky130_fd_pr__nfet_01v8, Bin 036, W = 0.42, L = 20.0
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__b0_diff_36=6.6799e-10
+  sky130_fd_pr__nfet_01v8__pdits_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_36=-0.13837
+  sky130_fd_pr__nfet_01v8__b1_diff_36=2.9823e-8
+  sky130_fd_pr__nfet_01v8__pditsd_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_36=0.81197
+  sky130_fd_pr__nfet_01v8__u0_diff_36=-0.0031366
+  sky130_fd_pr__nfet_01v8__ags_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_36=7.0971e-5
+  sky130_fd_pr__nfet_01v8__ua_diff_36=7.4306e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_36=-1.172e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_36=0.00036145
+  sky130_fd_pr__nfet_01v8__a0_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_36=0.011079
*
* sky130_fd_pr__nfet_01v8, Bin 037, W = 0.42, L = 2.0
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__kt1_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_37=-0.016478
+  sky130_fd_pr__nfet_01v8__b0_diff_37=1.0042e-8
+  sky130_fd_pr__nfet_01v8__pdits_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_37=-0.076269
+  sky130_fd_pr__nfet_01v8__b1_diff_37=5.9759e-8
+  sky130_fd_pr__nfet_01v8__pditsd_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_37=0.56465
+  sky130_fd_pr__nfet_01v8__u0_diff_37=-0.0054879
+  sky130_fd_pr__nfet_01v8__ags_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_37=-0.0029444
+  sky130_fd_pr__nfet_01v8__ua_diff_37=1.7334e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_37=-2.4886e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_37=-0.0019302
+  sky130_fd_pr__nfet_01v8__a0_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_37=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 038, W = 0.42, L = 4.0
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__a0_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_38=-0.0064116
+  sky130_fd_pr__nfet_01v8__b0_diff_38=-2.365e-8
+  sky130_fd_pr__nfet_01v8__pdits_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_38=-0.1251
+  sky130_fd_pr__nfet_01v8__b1_diff_38=6.7905e-8
+  sky130_fd_pr__nfet_01v8__pditsd_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_38=0.76257
+  sky130_fd_pr__nfet_01v8__u0_diff_38=-0.0034069
+  sky130_fd_pr__nfet_01v8__ags_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_38=0.0027273
+  sky130_fd_pr__nfet_01v8__ua_diff_38=1.0335e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_38=-1.0155e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_38=-0.00013396
*
* sky130_fd_pr__nfet_01v8, Bin 039, W = 0.42, L = 8.0
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__tvoff_diff_39=0.00011651
+  sky130_fd_pr__nfet_01v8__a0_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_39=0.0094213
+  sky130_fd_pr__nfet_01v8__pdits_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_39=-0.12613
+  sky130_fd_pr__nfet_01v8__b0_diff_39=3.0127e-8
+  sky130_fd_pr__nfet_01v8__b1_diff_39=1.2883e-7
+  sky130_fd_pr__nfet_01v8__pditsd_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_39=0.71859
+  sky130_fd_pr__nfet_01v8__u0_diff_39=-0.0033995
+  sky130_fd_pr__nfet_01v8__ags_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_39=-0.0039806
+  sky130_fd_pr__nfet_01v8__ua_diff_39=8.7608e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_39=-1.6334e-19
*
* sky130_fd_pr__nfet_01v8, Bin 040, W = 0.42, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__tvoff_diff_40=-0.0013808
+  sky130_fd_pr__nfet_01v8__a0_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_40=1855.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_40=-0.014644
+  sky130_fd_pr__nfet_01v8__pdits_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_40=-0.087821
+  sky130_fd_pr__nfet_01v8__b1_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_40=0.73736
+  sky130_fd_pr__nfet_01v8__u0_diff_40=0.0022185
+  sky130_fd_pr__nfet_01v8__ags_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_40=7.3348e-5
+  sky130_fd_pr__nfet_01v8__ua_diff_40=-6.3825e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_40=6.55e-19
*
* sky130_fd_pr__nfet_01v8, Bin 041, W = 0.42, L = 0.18
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__eta0_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_41=-2.2736e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_41=-0.00076032
+  sky130_fd_pr__nfet_01v8__a0_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_41=-13158.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_41=-0.034921
+  sky130_fd_pr__nfet_01v8__pdits_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_41=-0.10707
+  sky130_fd_pr__nfet_01v8__b1_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_41=1.1282
+  sky130_fd_pr__nfet_01v8__u0_diff_41=-0.0065285
+  sky130_fd_pr__nfet_01v8__ags_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_41=-0.0041958
+  sky130_fd_pr__nfet_01v8__ua_diff_41=2.7564e-11
*
* sky130_fd_pr__nfet_01v8, Bin 042, W = 0.42, L = 0.5
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__ua_diff_42=1.5471e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_42=-1.3038e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_42=-0.0020275
+  sky130_fd_pr__nfet_01v8__a0_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_42=-3055.8
+  sky130_fd_pr__nfet_01v8__kt1_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_42=0.0079242
+  sky130_fd_pr__nfet_01v8__pdits_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_42=-0.085417
+  sky130_fd_pr__nfet_01v8__b1_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_42=0.67583
+  sky130_fd_pr__nfet_01v8__u0_diff_42=-0.0046047
+  sky130_fd_pr__nfet_01v8__ags_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_42=0.0039683
*
* sky130_fd_pr__nfet_01v8, Bin 043, W = 0.55, L = 1.0
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__ags_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_43=0.0032814
+  sky130_fd_pr__nfet_01v8__ua_diff_43=5.5055e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_43=5.3284e-20
+  sky130_fd_pr__nfet_01v8__tvoff_diff_43=-0.0012175
+  sky130_fd_pr__nfet_01v8__a0_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_43=0.013261
+  sky130_fd_pr__nfet_01v8__pdits_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_43=8.6965e-8
+  sky130_fd_pr__nfet_01v8__voff_diff_43=-0.09315
+  sky130_fd_pr__nfet_01v8__b1_diff_43=6.9528e-9
+  sky130_fd_pr__nfet_01v8__pditsd_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_43=0.66652
+  sky130_fd_pr__nfet_01v8__u0_diff_43=-0.0020805
*
* sky130_fd_pr__nfet_01v8, Bin 044, W = 0.55, L = 2.0
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__pclm_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_44=0.75122
+  sky130_fd_pr__nfet_01v8__u0_diff_44=-0.006668
+  sky130_fd_pr__nfet_01v8__ags_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_44=-0.004111
+  sky130_fd_pr__nfet_01v8__ua_diff_44=2.0025e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_44=-4.8209e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_44=-0.0016217
+  sky130_fd_pr__nfet_01v8__a0_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_44=0.010156
+  sky130_fd_pr__nfet_01v8__pdits_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_44=7.0112e-9
+  sky130_fd_pr__nfet_01v8__voff_diff_44=-0.10091
+  sky130_fd_pr__nfet_01v8__b1_diff_44=9.8129e-8
+  sky130_fd_pr__nfet_01v8__pditsd_diff_44=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 045, W = 0.55, L = 4.0
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__pditsd_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_45=0.68645
+  sky130_fd_pr__nfet_01v8__u0_diff_45=-0.003889
+  sky130_fd_pr__nfet_01v8__ags_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_45=-0.0012654
+  sky130_fd_pr__nfet_01v8__ua_diff_45=1.1458e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_45=-1.9509e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_45=-0.00059293
+  sky130_fd_pr__nfet_01v8__a0_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_45=0.0051537
+  sky130_fd_pr__nfet_01v8__pdits_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_45=9.5011e-9
+  sky130_fd_pr__nfet_01v8__voff_diff_45=-0.10091
+  sky130_fd_pr__nfet_01v8__b1_diff_45=4.309e-8
*
* sky130_fd_pr__nfet_01v8, Bin 046, W = 0.55, L = 8.0
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__pdits_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_46=-0.11715
+  sky130_fd_pr__nfet_01v8__b1_diff_46=7.9566e-8
+  sky130_fd_pr__nfet_01v8__pditsd_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_46=0.83192
+  sky130_fd_pr__nfet_01v8__u0_diff_46=-0.0022816
+  sky130_fd_pr__nfet_01v8__ags_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_46=0.00031106
+  sky130_fd_pr__nfet_01v8__ua_diff_46=6.4629e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_46=-7.4503e-22
+  sky130_fd_pr__nfet_01v8__tvoff_diff_46=9.173e-5
+  sky130_fd_pr__nfet_01v8__a0_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_46=0.010481
+  sky130_fd_pr__nfet_01v8__b0_diff_46=1.5128e-10
*
* sky130_fd_pr__nfet_01v8, Bin 047, W = 0.55, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__b0_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_47=-0.070588
+  sky130_fd_pr__nfet_01v8__b1_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_47=0.648
+  sky130_fd_pr__nfet_01v8__u0_diff_47=-0.0038493
+  sky130_fd_pr__nfet_01v8__ags_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_47=-0.00088012
+  sky130_fd_pr__nfet_01v8__ua_diff_47=1.6315e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_47=-6.6985e-20
+  sky130_fd_pr__nfet_01v8__tvoff_diff_47=-0.0012742
+  sky130_fd_pr__nfet_01v8__a0_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_47=649.63
+  sky130_fd_pr__nfet_01v8__kt1_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_47=-0.014637
*
* sky130_fd_pr__nfet_01v8, Bin 048, W = 0.55, L = 0.5
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__kt1_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_48=-6915.2
+  sky130_fd_pr__nfet_01v8__vth0_diff_48=-0.00021304
+  sky130_fd_pr__nfet_01v8__b0_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_48=-0.082997
+  sky130_fd_pr__nfet_01v8__b1_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_48=0.66798
+  sky130_fd_pr__nfet_01v8__u0_diff_48=-0.0018701
+  sky130_fd_pr__nfet_01v8__ags_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_48=-0.00087423
+  sky130_fd_pr__nfet_01v8__ua_diff_48=3.9332e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_48=-3.7598e-21
+  sky130_fd_pr__nfet_01v8__tvoff_diff_48=-0.0022201
+  sky130_fd_pr__nfet_01v8__a0_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_48=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 049, W = 0.64, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__a0_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_49=4130.2
+  sky130_fd_pr__nfet_01v8__vth0_diff_49=0.017766
+  sky130_fd_pr__nfet_01v8__b0_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_49=-0.073864
+  sky130_fd_pr__nfet_01v8__b1_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_49=0.59343
+  sky130_fd_pr__nfet_01v8__u0_diff_49=-0.0026796
+  sky130_fd_pr__nfet_01v8__ags_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_49=0.0021621
+  sky130_fd_pr__nfet_01v8__ua_diff_49=1.1487e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_49=-1.3093e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_49=-0.0012604
*
* sky130_fd_pr__nfet_01v8, Bin 050, W = 0.84, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__tvoff_diff_50=-0.0020453
+  sky130_fd_pr__nfet_01v8__a0_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_50=7078.7
+  sky130_fd_pr__nfet_01v8__kt1_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_50=-0.012537
+  sky130_fd_pr__nfet_01v8__pdits_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_50=-0.046951
+  sky130_fd_pr__nfet_01v8__b1_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_50=0.41011
+  sky130_fd_pr__nfet_01v8__u0_diff_50=-0.0025461
+  sky130_fd_pr__nfet_01v8__ags_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_50=-0.00063737
+  sky130_fd_pr__nfet_01v8__ua_diff_50=1.0629e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_50=-4.8113e-21
*
* sky130_fd_pr__nfet_01v8, Bin 051, W = 0.74, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__nfactor_diff_51=0.10603823
+  sky130_fd_pr__nfet_01v8__keta_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_51=-3.00003e-14
+  sky130_fd_pr__nfet_01v8__pclm_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_51=-0.00170921
+  sky130_fd_pr__nfet_01v8__ags_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_51=0.00019725
+  sky130_fd_pr__nfet_01v8__voff_diff_51=-0.05847488
+  sky130_fd_pr__nfet_01v8__k2_diff_51=-0.00162947
+  sky130_fd_pr__nfet_01v8__kt1_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_51=1388.60586357
+  sky130_fd_pr__nfet_01v8__vth0_diff_51=0.00556959
*
* sky130_fd_pr__nfet_01v8, Bin 052, W = 0.36, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__ub_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_52=2522.7
+  sky130_fd_pr__nfet_01v8__kt1_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_52=0.042691
+  sky130_fd_pr__nfet_01v8__pdits_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_52=0.0031326
+  sky130_fd_pr__nfet_01v8__nfactor_diff_52=0.93967
+  sky130_fd_pr__nfet_01v8__keta_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_52=-0.011632
+  sky130_fd_pr__nfet_01v8__ua_diff_52=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 053, W = 0.39, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__ua_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_53=1928.2
+  sky130_fd_pr__nfet_01v8__kt1_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_53=0.032658
+  sky130_fd_pr__nfet_01v8__pdits_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_53=0.0029052
+  sky130_fd_pr__nfet_01v8__nfactor_diff_53=0.83163
+  sky130_fd_pr__nfet_01v8__keta_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_53=-0.009063
*
* sky130_fd_pr__nfet_01v8, Bin 054, W = 0.52, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__keta_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_54=-0.00038398
+  sky130_fd_pr__nfet_01v8__ua_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_54=2675.4
+  sky130_fd_pr__nfet_01v8__kt1_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_54=0.00010821
+  sky130_fd_pr__nfet_01v8__pdits_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_54=0.0028323
+  sky130_fd_pr__nfet_01v8__nfactor_diff_54=0.44435
*
* sky130_fd_pr__nfet_01v8, Bin 055, W = 0.54, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__pclm_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_55=0.0032327
+  sky130_fd_pr__nfet_01v8__nfactor_diff_55=0.33971
+  sky130_fd_pr__nfet_01v8__keta_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_55=-0.00049375
+  sky130_fd_pr__nfet_01v8__ua_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_55=2857.4
+  sky130_fd_pr__nfet_01v8__kt1_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_55=0.00055169
+  sky130_fd_pr__nfet_01v8__pdits_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_55=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 056, W = 0.58, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__pditsd_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_56=0.0013065
+  sky130_fd_pr__nfet_01v8__nfactor_diff_56=0.36133
+  sky130_fd_pr__nfet_01v8__keta_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_56=-0.0010528
+  sky130_fd_pr__nfet_01v8__ua_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_56=5027.9
+  sky130_fd_pr__nfet_01v8__kt1_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_56=-7.693e-5
+  sky130_fd_pr__nfet_01v8__pdits_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_56=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 057, W = 0.6, L = 0.15
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__pdits_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_57=-0.00098689
+  sky130_fd_pr__nfet_01v8__nfactor_diff_57=0.51825
+  sky130_fd_pr__nfet_01v8__keta_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_57=0.00092631
+  sky130_fd_pr__nfet_01v8__ua_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_57=7175.7
+  sky130_fd_pr__nfet_01v8__kt1_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_57=-0.0014905
+  sky130_fd_pr__nfet_01v8__b0_diff_57=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 058, W = 0.61, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__b0_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_58=-0.00046704
+  sky130_fd_pr__nfet_01v8__nfactor_diff_58=0.48571
+  sky130_fd_pr__nfet_01v8__keta_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_58=0.00058075
+  sky130_fd_pr__nfet_01v8__ua_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_58=8409.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_58=-0.0011114
*
* sky130_fd_pr__nfet_01v8, Bin 059, W = 0.65, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__kt1_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_59=5838.2
+  sky130_fd_pr__nfet_01v8__vth0_diff_59=-0.00066578
+  sky130_fd_pr__nfet_01v8__b0_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_59=0.0010877
+  sky130_fd_pr__nfet_01v8__nfactor_diff_59=0.55642
+  sky130_fd_pr__nfet_01v8__keta_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_59=0.00023346
+  sky130_fd_pr__nfet_01v8__ua_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_59=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 060, W = 0.65, L = 0.18
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__vsat_diff_60=12193.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_60=0.00035634
+  sky130_fd_pr__nfet_01v8__pdits_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_60=0.0018309
+  sky130_fd_pr__nfet_01v8__nfactor_diff_60=0.54191
+  sky130_fd_pr__nfet_01v8__keta_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_60=-0.0037472
+  sky130_fd_pr__nfet_01v8__ua_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_60=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 061, W = 0.65, L = 0.25
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__tvoff_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_61=16254.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_61=-0.002334
+  sky130_fd_pr__nfet_01v8__pdits_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_61=0.0015766
+  sky130_fd_pr__nfet_01v8__nfactor_diff_61=0.92024
+  sky130_fd_pr__nfet_01v8__keta_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_61=-0.0013286
+  sky130_fd_pr__nfet_01v8__ua_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_61=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 062, W = 0.65, L = 0.5
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__tvoff_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_62=14599.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_62=-0.0023875
+  sky130_fd_pr__nfet_01v8__pdits_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_62=0.0015543
+  sky130_fd_pr__nfet_01v8__nfactor_diff_62=0.35686
+  sky130_fd_pr__nfet_01v8__keta_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_62=-0.0015962
+  sky130_fd_pr__nfet_01v8__ua_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_62=0.0
.include "sky130_fd_pr__nfet_01v8.pm3.spice"
