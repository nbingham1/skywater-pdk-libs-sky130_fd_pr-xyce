* Bipolar transistor I-V characteristic

* Include SkyWater sky130 device models
.include "../../../models/corners/tt/nonfet.spice"
.include "../sky130_fd_pr__npn_05v5__wafer.corner.spice"

* Base bias
Rb 1 2 680
X1 3 2 0 0 sky130_fd_pr__npn_05v5_W1p00L2p00 M=1
Rc 3 4 100

* DC source for current measure
Vic 4 5 DC 0V
Vbb 1 0 DC 0V
Vce 5 0 DC 0V

.control
* Sweep Vce from 0 to 1.8V
dc Vce 0 1.8 0.01 vbb 0 1.2 0.01
wrdata sky130_fd_pr__npn_05v5_W1p00L2p00__iv.data -Vic#branch V ( 1 ) V ( 3 )

* Sweep Vce from 0 to 3.3V, Vbb from 0 to 2.0V
dc Vce 0 3.3 0.02 Vbb 0.6 0.9 0.01
let beta=Vic#branch / Vbb#branch
wrdata sky130_fd_pr__npn_05v5_W1p00L2p00__beta.data beta V ( 2 ) V ( 3 )
echo maximum beta
print maximum ( beta )
quit
.endc
.end
