* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 63
.param
+  sky130_fd_pr__nfet_01v8__toxe_mult=0.948
+  sky130_fd_pr__nfet_01v8__rshn_mult=1.0
+  sky130_fd_pr__nfet_01v8__overlap_mult=0.94816
+  sky130_fd_pr__nfet_01v8__lint_diff=1.7325e-8
+  sky130_fd_pr__nfet_01v8__wint_diff=-3.2175e-8
+  sky130_fd_pr__nfet_01v8__dlc_diff=12.773e-9
+  sky130_fd_pr__nfet_01v8__dwc_diff=-3.2175e-8
*
* sky130_fd_pr__nfet_01v8, Bin 000, W = 1.26, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__voff_diff_0=-0.092208
+  sky130_fd_pr__nfet_01v8__kt1_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_0=-1.7055e-19
+  sky130_fd_pr__nfet_01v8__pditsd_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_0=9.7995e-11
+  sky130_fd_pr__nfet_01v8__vsat_diff_0=-45772.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_0=0.00062266
+  sky130_fd_pr__nfet_01v8__ags_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_0=0.064071
+  sky130_fd_pr__nfet_01v8__vth0_diff_0=-0.13212
+  sky130_fd_pr__nfet_01v8__nfactor_diff_0=0.3527
+  sky130_fd_pr__nfet_01v8__u0_diff_0=-0.0078344
+  sky130_fd_pr__nfet_01v8__eta0_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_0=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 001, W = 1.68, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__eta0_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_1=-0.070854
+  sky130_fd_pr__nfet_01v8__kt1_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_1=-2.3753e-19
+  sky130_fd_pr__nfet_01v8__pditsd_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_1=2.9323e-10
+  sky130_fd_pr__nfet_01v8__vsat_diff_1=-38447.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_1=0.00067814
+  sky130_fd_pr__nfet_01v8__ags_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_1=0.061447
+  sky130_fd_pr__nfet_01v8__vth0_diff_1=-0.10045
+  sky130_fd_pr__nfet_01v8__nfactor_diff_1=0.55865
+  sky130_fd_pr__nfet_01v8__u0_diff_1=-0.0051543
*
* sky130_fd_pr__nfet_01v8, Bin 002, W = 1.0, L = 1.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__nfactor_diff_2=1.3489
+  sky130_fd_pr__nfet_01v8__u0_diff_2=0.00076854
+  sky130_fd_pr__nfet_01v8__vth0_diff_2=-0.0029124
+  sky130_fd_pr__nfet_01v8__eta0_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_2=-0.16449
+  sky130_fd_pr__nfet_01v8__ub_diff_2=2.7741e-19
+  sky130_fd_pr__nfet_01v8__kt1_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_2=2.9297e-12
+  sky130_fd_pr__nfet_01v8__vsat_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_2=0.00090563
+  sky130_fd_pr__nfet_01v8__ags_diff_2=-0.15706
+  sky130_fd_pr__nfet_01v8__a0_diff_2=0.4
+  sky130_fd_pr__nfet_01v8__b0_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_2=-0.00537
*
* sky130_fd_pr__nfet_01v8, Bin 003, W = 1.0, L = 2.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__keta_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_3=-0.0067371
+  sky130_fd_pr__nfet_01v8__nfactor_diff_3=1.0669
+  sky130_fd_pr__nfet_01v8__u0_diff_3=0.00036601
+  sky130_fd_pr__nfet_01v8__vth0_diff_3=-0.0019543
+  sky130_fd_pr__nfet_01v8__eta0_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_3=-0.17244
+  sky130_fd_pr__nfet_01v8__ub_diff_3=2.4903e-19
+  sky130_fd_pr__nfet_01v8__kt1_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_3=1.4357e-12
+  sky130_fd_pr__nfet_01v8__vsat_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_3=0.001068
+  sky130_fd_pr__nfet_01v8__ags_diff_3=-0.050995
+  sky130_fd_pr__nfet_01v8__a0_diff_3=0.090682
+  sky130_fd_pr__nfet_01v8__b0_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_3=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 004, W = 1.0, L = 4.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__pdits_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_4=-0.0019298
+  sky130_fd_pr__nfet_01v8__nfactor_diff_4=0.93949
+  sky130_fd_pr__nfet_01v8__u0_diff_4=-0.0010157
+  sky130_fd_pr__nfet_01v8__vth0_diff_4=0.0071716
+  sky130_fd_pr__nfet_01v8__eta0_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_4=-0.21377
+  sky130_fd_pr__nfet_01v8__ub_diff_4=1.1623e-19
+  sky130_fd_pr__nfet_01v8__kt1_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_4=6.0814e-12
+  sky130_fd_pr__nfet_01v8__vsat_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_4=0.0019039
+  sky130_fd_pr__nfet_01v8__ags_diff_4=0.0029314
+  sky130_fd_pr__nfet_01v8__a0_diff_4=0.0018101
+  sky130_fd_pr__nfet_01v8__b0_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_4=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 005, W = 1.0, L = 8.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__pdits_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_5=0.0015842
+  sky130_fd_pr__nfet_01v8__nfactor_diff_5=0.89143
+  sky130_fd_pr__nfet_01v8__u0_diff_5=-0.0012539
+  sky130_fd_pr__nfet_01v8__vth0_diff_5=0.0047277
+  sky130_fd_pr__nfet_01v8__eta0_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_5=-0.21387
+  sky130_fd_pr__nfet_01v8__ub_diff_5=1.1829e-19
+  sky130_fd_pr__nfet_01v8__kt1_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_5=6.317e-12
+  sky130_fd_pr__nfet_01v8__vsat_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_5=0.0025066
+  sky130_fd_pr__nfet_01v8__ags_diff_5=-0.015678
+  sky130_fd_pr__nfet_01v8__a0_diff_5=0.017921
+  sky130_fd_pr__nfet_01v8__b0_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_5=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 006, W = 1.0, L = 0.15
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__pclm_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_6=0.060131
+  sky130_fd_pr__nfet_01v8__nfactor_diff_6=0.64009
+  sky130_fd_pr__nfet_01v8__u0_diff_6=-0.0079755
+  sky130_fd_pr__nfet_01v8__vth0_diff_6=-0.11261
+  sky130_fd_pr__nfet_01v8__eta0_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_6=-0.10887
+  sky130_fd_pr__nfet_01v8__ub_diff_6=-2.3042e-19
+  sky130_fd_pr__nfet_01v8__kt1_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_6=8.7967e-11
+  sky130_fd_pr__nfet_01v8__vsat_diff_6=-47470.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_6=0.00095785
+  sky130_fd_pr__nfet_01v8__ags_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_6=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 007, W = 1.0, L = 0.18
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__tvoff_diff_7=0.00023658
+  sky130_fd_pr__nfet_01v8__b0_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_7=0.032569
+  sky130_fd_pr__nfet_01v8__nfactor_diff_7=0.80109
+  sky130_fd_pr__nfet_01v8__u0_diff_7=-0.0048082
+  sky130_fd_pr__nfet_01v8__vth0_diff_7=-0.08417
+  sky130_fd_pr__nfet_01v8__eta0_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_7=-0.10775
+  sky130_fd_pr__nfet_01v8__ub_diff_7=5.3746e-20
+  sky130_fd_pr__nfet_01v8__kt1_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_7=7.3291e-11
+  sky130_fd_pr__nfet_01v8__vsat_diff_7=-42109.0
+  sky130_fd_pr__nfet_01v8__a0_diff_7=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 008, W = 1.0, L = 0.25
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__a0_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_8=3.4905e-11
+  sky130_fd_pr__nfet_01v8__tvoff_diff_8=0.00054176
+  sky130_fd_pr__nfet_01v8__b0_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_8=0.0090206
+  sky130_fd_pr__nfet_01v8__nfactor_diff_8=0.92698
+  sky130_fd_pr__nfet_01v8__u0_diff_8=-0.0023881
+  sky130_fd_pr__nfet_01v8__vth0_diff_8=-0.045052
+  sky130_fd_pr__nfet_01v8__eta0_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_8=-0.14541
+  sky130_fd_pr__nfet_01v8__ub_diff_8=3.627e-19
+  sky130_fd_pr__nfet_01v8__kt1_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_8=-38315.0
*
* sky130_fd_pr__nfet_01v8, Bin 009, W = 1.0, L = 0.5
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__kt1_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_9=1.0588e-20
+  sky130_fd_pr__nfet_01v8__vsat_diff_9=-20000.0
+  sky130_fd_pr__nfet_01v8__a0_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_9=1.1384e-11
+  sky130_fd_pr__nfet_01v8__tvoff_diff_9=0.0013235
+  sky130_fd_pr__nfet_01v8__b0_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_9=0.0016241
+  sky130_fd_pr__nfet_01v8__nfactor_diff_9=1.0743
+  sky130_fd_pr__nfet_01v8__u0_diff_9=-0.002489
+  sky130_fd_pr__nfet_01v8__vth0_diff_9=0.0024268
+  sky130_fd_pr__nfet_01v8__eta0_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_9=-0.16654
*
* sky130_fd_pr__nfet_01v8, Bin 010, W = 2.0, L = 0.15
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__ags_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_10=0.065173
+  sky130_fd_pr__nfet_01v8__ua_diff_10=1.6099e-10
+  sky130_fd_pr__nfet_01v8__eta0_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_10=-1.7509e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_10=0.00056884
+  sky130_fd_pr__nfet_01v8__a0_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_10=-41913.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_10=-0.091578
+  sky130_fd_pr__nfet_01v8__pdits_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_10=-0.086335
+  sky130_fd_pr__nfet_01v8__b1_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_10=0.63287
+  sky130_fd_pr__nfet_01v8__u0_diff_10=-0.0056082
*
* sky130_fd_pr__nfet_01v8, Bin 011, W = 3.0, L = 1.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__pclm_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_11=1.1484
+  sky130_fd_pr__nfet_01v8__u0_diff_11=-8.0462e-5
+  sky130_fd_pr__nfet_01v8__ags_diff_11=-0.0856
+  sky130_fd_pr__nfet_01v8__keta_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_11=-0.0030943
+  sky130_fd_pr__nfet_01v8__ua_diff_11=3.8253e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_11=1.3598e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_11=0.00090432
+  sky130_fd_pr__nfet_01v8__a0_diff_11=0.0042624
+  sky130_fd_pr__nfet_01v8__rdsw_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_11=0.010196
+  sky130_fd_pr__nfet_01v8__pdits_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_11=-0.15799
+  sky130_fd_pr__nfet_01v8__b1_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_11=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 012, W = 3.0, L = 2.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__pditsd_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_12=1.5376
+  sky130_fd_pr__nfet_01v8__u0_diff_12=-0.0020612
+  sky130_fd_pr__nfet_01v8__ags_diff_12=0.053123
+  sky130_fd_pr__nfet_01v8__keta_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_12=-0.0043376
+  sky130_fd_pr__nfet_01v8__ua_diff_12=9.7365e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_12=-8.334e-20
+  sky130_fd_pr__nfet_01v8__tvoff_diff_12=0.00070107
+  sky130_fd_pr__nfet_01v8__a0_diff_12=-0.043697
+  sky130_fd_pr__nfet_01v8__rdsw_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_12=0.017497
+  sky130_fd_pr__nfet_01v8__pdits_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_12=-0.14715
+  sky130_fd_pr__nfet_01v8__b1_diff_12=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 013, W = 3.0, L = 4.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__pdits_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_13=-0.17609
+  sky130_fd_pr__nfet_01v8__b1_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_13=0.94848
+  sky130_fd_pr__nfet_01v8__u0_diff_13=-0.0031539
+  sky130_fd_pr__nfet_01v8__ags_diff_13=0.057876
+  sky130_fd_pr__nfet_01v8__keta_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_13=-0.0034486
+  sky130_fd_pr__nfet_01v8__ua_diff_13=2.3484e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_13=-2.0159e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_13=0.00097957
+  sky130_fd_pr__nfet_01v8__a0_diff_13=-0.075963
+  sky130_fd_pr__nfet_01v8__rdsw_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_13=0.015153
+  sky130_fd_pr__nfet_01v8__b0_diff_13=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 014, W = 3.0, L = 8.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__b0_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_14=-0.19876
+  sky130_fd_pr__nfet_01v8__b1_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_14=0.93044
+  sky130_fd_pr__nfet_01v8__u0_diff_14=-0.0022485
+  sky130_fd_pr__nfet_01v8__ags_diff_14=0.02164
+  sky130_fd_pr__nfet_01v8__keta_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_14=8.7155e-6
+  sky130_fd_pr__nfet_01v8__ua_diff_14=8.8314e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_14=-1.3143e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_14=0.0017711
+  sky130_fd_pr__nfet_01v8__a0_diff_14=-0.02545
+  sky130_fd_pr__nfet_01v8__rdsw_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_14=0.014266
*
* sky130_fd_pr__nfet_01v8, Bin 015, W = 3.0, L = 0.15
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__kt1_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_15=-35036.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_15=-0.097639
+  sky130_fd_pr__nfet_01v8__b0_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_15=-0.092395
+  sky130_fd_pr__nfet_01v8__b1_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_15=0.36426
+  sky130_fd_pr__nfet_01v8__u0_diff_15=-0.0079323
+  sky130_fd_pr__nfet_01v8__ags_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_15=0.066641
+  sky130_fd_pr__nfet_01v8__ua_diff_15=2.0806e-10
+  sky130_fd_pr__nfet_01v8__eta0_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_15=-6.6411e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_15=0.00031221
+  sky130_fd_pr__nfet_01v8__a0_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_15=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 016, W = 3.0, L = 0.18
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__a0_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_16=-29294.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_16=-0.052668
+  sky130_fd_pr__nfet_01v8__b0_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_16=-0.12792
+  sky130_fd_pr__nfet_01v8__b1_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_16=0.82563
+  sky130_fd_pr__nfet_01v8__u0_diff_16=-0.004604
+  sky130_fd_pr__nfet_01v8__ags_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_16=0.042932
+  sky130_fd_pr__nfet_01v8__ua_diff_16=5.0291e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_16=1.0238e-20
+  sky130_fd_pr__nfet_01v8__tvoff_diff_16=0.0004294
*
* sky130_fd_pr__nfet_01v8, Bin 017, W = 3.0, L = 0.25
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__tvoff_diff_17=0.0015274
+  sky130_fd_pr__nfet_01v8__a0_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_17=-20000.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_17=-0.017108
+  sky130_fd_pr__nfet_01v8__pdits_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_17=-0.11831
+  sky130_fd_pr__nfet_01v8__b0_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_17=2.162
+  sky130_fd_pr__nfet_01v8__u0_diff_17=-0.00086326
+  sky130_fd_pr__nfet_01v8__ags_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_17=0.013739
+  sky130_fd_pr__nfet_01v8__ua_diff_17=1.6132e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_17=1.5827e-19
*
* sky130_fd_pr__nfet_01v8, Bin 018, W = 3.0, L = 0.5
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__ub_diff_18=1.0693e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_18=0.0015145
+  sky130_fd_pr__nfet_01v8__a0_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_18=-6267.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_18=-0.003475
+  sky130_fd_pr__nfet_01v8__pdits_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_18=-0.12451
+  sky130_fd_pr__nfet_01v8__b0_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_18=1.8738
+  sky130_fd_pr__nfet_01v8__u0_diff_18=-0.0014893
+  sky130_fd_pr__nfet_01v8__ags_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_18=0.0015584
+  sky130_fd_pr__nfet_01v8__ua_diff_18=7.5866e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_18=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 019, W = 5.0, L = 1.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__eta0_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_19=2.7522e-12
+  sky130_fd_pr__nfet_01v8__ub_diff_19=1.1735e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_19=0.00055238
+  sky130_fd_pr__nfet_01v8__a0_diff_19=0.030186
+  sky130_fd_pr__nfet_01v8__rdsw_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_19=0.015834
+  sky130_fd_pr__nfet_01v8__pdits_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_19=-0.15099
+  sky130_fd_pr__nfet_01v8__b0_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_19=0.91418
+  sky130_fd_pr__nfet_01v8__u0_diff_19=-0.00032054
+  sky130_fd_pr__nfet_01v8__ags_diff_19=0.080308
+  sky130_fd_pr__nfet_01v8__keta_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_19=0.0021661
*
* sky130_fd_pr__nfet_01v8, Bin 020, W = 5.0, L = 2.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__ua_diff_20=1.3722e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_20=-2.3913e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_20=0.00055775
+  sky130_fd_pr__nfet_01v8__a0_diff_20=-0.096915
+  sky130_fd_pr__nfet_01v8__rdsw_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_20=0.014112
+  sky130_fd_pr__nfet_01v8__pdits_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_20=-0.14025
+  sky130_fd_pr__nfet_01v8__b1_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_20=1.4934
+  sky130_fd_pr__nfet_01v8__u0_diff_20=-0.0032532
+  sky130_fd_pr__nfet_01v8__ags_diff_20=0.065381
+  sky130_fd_pr__nfet_01v8__keta_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_20=-0.00469
*
* sky130_fd_pr__nfet_01v8, Bin 021, W = 5.0, L = 4.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__ags_diff_21=0.0057722
+  sky130_fd_pr__nfet_01v8__keta_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_21=-0.00328
+  sky130_fd_pr__nfet_01v8__ua_diff_21=8.6809e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_21=-1.4951e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_21=0.00086952
+  sky130_fd_pr__nfet_01v8__a0_diff_21=-0.0107
+  sky130_fd_pr__nfet_01v8__rdsw_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_21=0.011791
+  sky130_fd_pr__nfet_01v8__pdits_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_21=-0.15594
+  sky130_fd_pr__nfet_01v8__b1_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_21=1.1013
+  sky130_fd_pr__nfet_01v8__u0_diff_21=-0.0019909
*
* sky130_fd_pr__nfet_01v8, Bin 022, W = 5.0, L = 8.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__pclm_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_22=2.0594
+  sky130_fd_pr__nfet_01v8__u0_diff_22=-0.0013364
+  sky130_fd_pr__nfet_01v8__ags_diff_22=0.051684
+  sky130_fd_pr__nfet_01v8__keta_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_22=0.00021745
+  sky130_fd_pr__nfet_01v8__ua_diff_22=6.6072e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_22=-5.991e-20
+  sky130_fd_pr__nfet_01v8__tvoff_diff_22=0.0018135
+  sky130_fd_pr__nfet_01v8__a0_diff_22=-0.069442
+  sky130_fd_pr__nfet_01v8__rdsw_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_22=0.019187
+  sky130_fd_pr__nfet_01v8__pdits_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_22=-0.14785
+  sky130_fd_pr__nfet_01v8__b1_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_22=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 023, W = 5.0, L = 0.15
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__pditsd_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_23=0.41231
+  sky130_fd_pr__nfet_01v8__u0_diff_23=-0.0031868
+  sky130_fd_pr__nfet_01v8__ags_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_23=0.057387
+  sky130_fd_pr__nfet_01v8__ua_diff_23=3.2545e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_23=-1.2193e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_23=0.00043062
+  sky130_fd_pr__nfet_01v8__a0_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_23=-27396.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_23=-0.070621
+  sky130_fd_pr__nfet_01v8__pdits_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_23=-0.06684
+  sky130_fd_pr__nfet_01v8__b1_diff_23=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 024, W = 5.0, L = 0.18
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__pdits_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_24=-0.10801
+  sky130_fd_pr__nfet_01v8__b1_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_24=0.73977
+  sky130_fd_pr__nfet_01v8__u0_diff_24=-0.01
+  sky130_fd_pr__nfet_01v8__ags_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_24=0.030058
+  sky130_fd_pr__nfet_01v8__ua_diff_24=1.0018e-10
+  sky130_fd_pr__nfet_01v8__eta0_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_24=-5.7461e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_24=0.00052686
+  sky130_fd_pr__nfet_01v8__a0_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_24=-19422.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_24=-0.036205
+  sky130_fd_pr__nfet_01v8__b0_diff_24=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 025, W = 5.0, L = 0.25
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__b0_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_25=-0.12568
+  sky130_fd_pr__nfet_01v8__b1_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_25=0.89736
+  sky130_fd_pr__nfet_01v8__u0_diff_25=-0.00076282
+  sky130_fd_pr__nfet_01v8__ags_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_25=0.013522
+  sky130_fd_pr__nfet_01v8__ua_diff_25=1.4882e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_25=1.7745e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_25=0.00039839
+  sky130_fd_pr__nfet_01v8__a0_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_25=-20000.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_25=-0.00416
*
* sky130_fd_pr__nfet_01v8, Bin 026, W = 5.0, L = 0.5
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__kt1_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_26=-8424.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_26=2.1783e-5
+  sky130_fd_pr__nfet_01v8__b0_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_26=-0.12329
+  sky130_fd_pr__nfet_01v8__b1_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_26=1.9195
+  sky130_fd_pr__nfet_01v8__u0_diff_26=-0.001181
+  sky130_fd_pr__nfet_01v8__ags_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_26=-0.0008125
+  sky130_fd_pr__nfet_01v8__ua_diff_26=5.7866e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_26=2.944e-20
+  sky130_fd_pr__nfet_01v8__tvoff_diff_26=0.0014635
+  sky130_fd_pr__nfet_01v8__a0_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_26=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 027, W = 7.0, L = 1.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__a0_diff_27=-0.0099235
+  sky130_fd_pr__nfet_01v8__rdsw_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_27=0.0036866
+  sky130_fd_pr__nfet_01v8__b0_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_27=-0.15275
+  sky130_fd_pr__nfet_01v8__b1_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_27=1.1725
+  sky130_fd_pr__nfet_01v8__u0_diff_27=-0.001336
+  sky130_fd_pr__nfet_01v8__ags_diff_27=0.012567
+  sky130_fd_pr__nfet_01v8__keta_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_27=-6.8657e-5
+  sky130_fd_pr__nfet_01v8__ua_diff_27=7.5127e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_27=3.0668e-20
+  sky130_fd_pr__nfet_01v8__tvoff_diff_27=0.0007405
*
* sky130_fd_pr__nfet_01v8, Bin 028, W = 7.0, L = 2.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__tvoff_diff_28=0.00053354
+  sky130_fd_pr__nfet_01v8__a0_diff_28=-0.08158
+  sky130_fd_pr__nfet_01v8__rdsw_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_28=0.020447
+  sky130_fd_pr__nfet_01v8__pdits_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_28=-0.16256
+  sky130_fd_pr__nfet_01v8__b0_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_28=1.0041
+  sky130_fd_pr__nfet_01v8__u0_diff_28=-0.0008184
+  sky130_fd_pr__nfet_01v8__ags_diff_28=0.085346
+  sky130_fd_pr__nfet_01v8__keta_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_28=-0.0022986
+  sky130_fd_pr__nfet_01v8__ua_diff_28=5.9578e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_28=1.497e-20
*
* sky130_fd_pr__nfet_01v8, Bin 029, W = 7.0, L = 4.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__ub_diff_29=5.7665e-20
+  sky130_fd_pr__nfet_01v8__tvoff_diff_29=0.00079835
+  sky130_fd_pr__nfet_01v8__a0_diff_29=-0.089992
+  sky130_fd_pr__nfet_01v8__rdsw_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_29=0.014426
+  sky130_fd_pr__nfet_01v8__pdits_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_29=-0.16243
+  sky130_fd_pr__nfet_01v8__b0_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_29=0.88549
+  sky130_fd_pr__nfet_01v8__u0_diff_29=-0.00041967
+  sky130_fd_pr__nfet_01v8__ags_diff_29=0.073911
+  sky130_fd_pr__nfet_01v8__keta_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_29=-0.0036846
+  sky130_fd_pr__nfet_01v8__ua_diff_29=4.5264e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_29=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 030, W = 7.0, L = 8.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__eta0_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_30=-2.1952e-21
+  sky130_fd_pr__nfet_01v8__tvoff_diff_30=0.00096922
+  sky130_fd_pr__nfet_01v8__a0_diff_30=-0.041769
+  sky130_fd_pr__nfet_01v8__rdsw_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_30=0.018988
+  sky130_fd_pr__nfet_01v8__pdits_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_30=-0.15568
+  sky130_fd_pr__nfet_01v8__b1_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_30=0.88119
+  sky130_fd_pr__nfet_01v8__u0_diff_30=-0.0004775
+  sky130_fd_pr__nfet_01v8__ags_diff_30=0.050012
+  sky130_fd_pr__nfet_01v8__keta_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_30=-0.00027712
+  sky130_fd_pr__nfet_01v8__ua_diff_30=3.5649e-12
*
* sky130_fd_pr__nfet_01v8, Bin 031, W = 7.0, L = 0.15
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__ua_diff_31=2.1889e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_31=1.9277e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_31=-8.2467e-6
+  sky130_fd_pr__nfet_01v8__a0_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_31=-26014.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_31=-0.074679
+  sky130_fd_pr__nfet_01v8__pdits_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_31=-0.072443
+  sky130_fd_pr__nfet_01v8__b1_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_31=0.62721
+  sky130_fd_pr__nfet_01v8__u0_diff_31=-0.00067706
+  sky130_fd_pr__nfet_01v8__ags_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_31=0.058993
*
* sky130_fd_pr__nfet_01v8, Bin 032, W = 7.0, L = 0.18
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__ags_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_32=0.033554
+  sky130_fd_pr__nfet_01v8__ua_diff_32=8.9417e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_32=-4.4851e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_32=0.0010243
+  sky130_fd_pr__nfet_01v8__a0_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_32=-18748.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_32=-0.03961
+  sky130_fd_pr__nfet_01v8__pdits_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_32=-0.12432
+  sky130_fd_pr__nfet_01v8__b1_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_32=0.97595
+  sky130_fd_pr__nfet_01v8__u0_diff_32=-0.009415
*
* sky130_fd_pr__nfet_01v8, Bin 033, W = 7.0, L = 0.25
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__pclm_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_33=1.1882
+  sky130_fd_pr__nfet_01v8__u0_diff_33=-0.0009389
+  sky130_fd_pr__nfet_01v8__ags_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_33=0.015406
+  sky130_fd_pr__nfet_01v8__ua_diff_33=1.539e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_33=1.2331e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_33=0.00022332
+  sky130_fd_pr__nfet_01v8__a0_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_33=-20000.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_33=-0.0036613
+  sky130_fd_pr__nfet_01v8__pdits_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_33=-0.10283
+  sky130_fd_pr__nfet_01v8__b1_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_33=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 034, W = 7.0, L = 0.5
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__pditsd_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_34=1.0447
+  sky130_fd_pr__nfet_01v8__u0_diff_34=-0.0011518
+  sky130_fd_pr__nfet_01v8__ags_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_34=-0.001068
+  sky130_fd_pr__nfet_01v8__ua_diff_34=5.7302e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_34=2.5808e-20
+  sky130_fd_pr__nfet_01v8__tvoff_diff_34=0.0010508
+  sky130_fd_pr__nfet_01v8__a0_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_34=-6076.5
+  sky130_fd_pr__nfet_01v8__kt1_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_34=-0.0010719
+  sky130_fd_pr__nfet_01v8__pdits_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_34=-0.14874
+  sky130_fd_pr__nfet_01v8__b1_diff_34=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 035, W = 0.42, L = 1.0
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__pdits_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_35=-0.16063
+  sky130_fd_pr__nfet_01v8__b1_diff_35=2.1916e-8
+  sky130_fd_pr__nfet_01v8__pditsd_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_35=0.70032
+  sky130_fd_pr__nfet_01v8__u0_diff_35=-0.0032529
+  sky130_fd_pr__nfet_01v8__ags_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_35=-0.0073494
+  sky130_fd_pr__nfet_01v8__ua_diff_35=1.4141e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_35=9.0986e-20
+  sky130_fd_pr__nfet_01v8__tvoff_diff_35=0.00056884
+  sky130_fd_pr__nfet_01v8__a0_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_35=-0.015841
+  sky130_fd_pr__nfet_01v8__b0_diff_35=-3.0074e-8
*
* sky130_fd_pr__nfet_01v8, Bin 036, W = 0.42, L = 20.0
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__b0_diff_36=7.2143e-8
+  sky130_fd_pr__nfet_01v8__pdits_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_36=-0.21983
+  sky130_fd_pr__nfet_01v8__b1_diff_36=2.555e-8
+  sky130_fd_pr__nfet_01v8__pditsd_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_36=0.94441
+  sky130_fd_pr__nfet_01v8__u0_diff_36=-0.001827
+  sky130_fd_pr__nfet_01v8__ags_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_36=-0.00255
+  sky130_fd_pr__nfet_01v8__ua_diff_36=7.1952e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_36=1.1903e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_36=0.0025941
+  sky130_fd_pr__nfet_01v8__a0_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_36=0.010103
*
* sky130_fd_pr__nfet_01v8, Bin 037, W = 0.42, L = 2.0
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__kt1_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_37=-0.034629
+  sky130_fd_pr__nfet_01v8__b0_diff_37=1.5084e-7
+  sky130_fd_pr__nfet_01v8__pdits_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_37=-0.16551
+  sky130_fd_pr__nfet_01v8__b1_diff_37=4.3624e-8
+  sky130_fd_pr__nfet_01v8__pditsd_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_37=0.5737
+  sky130_fd_pr__nfet_01v8__u0_diff_37=-0.0043599
+  sky130_fd_pr__nfet_01v8__ags_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_37=-0.0049843
+  sky130_fd_pr__nfet_01v8__ua_diff_37=1.8074e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_37=-2.5396e-20
+  sky130_fd_pr__nfet_01v8__tvoff_diff_37=0.00089228
+  sky130_fd_pr__nfet_01v8__a0_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_37=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 038, W = 0.42, L = 4.0
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__a0_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_38=-0.018148
+  sky130_fd_pr__nfet_01v8__b0_diff_38=7.6522e-8
+  sky130_fd_pr__nfet_01v8__pdits_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_38=-0.19475
+  sky130_fd_pr__nfet_01v8__b1_diff_38=6.8599e-8
+  sky130_fd_pr__nfet_01v8__pditsd_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_38=0.60373
+  sky130_fd_pr__nfet_01v8__u0_diff_38=-0.0030142
+  sky130_fd_pr__nfet_01v8__ags_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_38=0.0028015
+  sky130_fd_pr__nfet_01v8__ua_diff_38=1.2381e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_38=1.0995e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_38=0.0016718
*
* sky130_fd_pr__nfet_01v8, Bin 039, W = 0.42, L = 8.0
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__tvoff_diff_39=0.0030764
+  sky130_fd_pr__nfet_01v8__a0_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_39=0.0047978
+  sky130_fd_pr__nfet_01v8__pdits_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_39=-0.20634
+  sky130_fd_pr__nfet_01v8__b0_diff_39=1.0347e-7
+  sky130_fd_pr__nfet_01v8__b1_diff_39=5.4285e-8
+  sky130_fd_pr__nfet_01v8__pditsd_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_39=0.90339
+  sky130_fd_pr__nfet_01v8__u0_diff_39=-0.0024064
+  sky130_fd_pr__nfet_01v8__ags_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_39=-0.0049858
+  sky130_fd_pr__nfet_01v8__ua_diff_39=9.289e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_39=7.14e-20
*
* sky130_fd_pr__nfet_01v8, Bin 040, W = 0.42, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__tvoff_diff_40=0.00092338
+  sky130_fd_pr__nfet_01v8__a0_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_40=-65000.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_40=-0.19319
+  sky130_fd_pr__nfet_01v8__pdits_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_40=-2.5003e-7
+  sky130_fd_pr__nfet_01v8__voff_diff_40=-0.070484
+  sky130_fd_pr__nfet_01v8__b1_diff_40=2.2838e-8
+  sky130_fd_pr__nfet_01v8__pditsd_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_40=1.3186
+  sky130_fd_pr__nfet_01v8__u0_diff_40=-0.0035405
+  sky130_fd_pr__nfet_01v8__ags_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_40=0.050198
+  sky130_fd_pr__nfet_01v8__ua_diff_40=2.6203e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_40=8.2092e-19
*
* sky130_fd_pr__nfet_01v8, Bin 041, W = 0.42, L = 0.18
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__eta0_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_41=2.8701e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_41=0.0015429
+  sky130_fd_pr__nfet_01v8__a0_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_41=-20000.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_41=-0.15
+  sky130_fd_pr__nfet_01v8__pdits_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_41=1.0704e-6
+  sky130_fd_pr__nfet_01v8__voff_diff_41=-0.058942
+  sky130_fd_pr__nfet_01v8__b1_diff_41=1.6377e-8
+  sky130_fd_pr__nfet_01v8__pditsd_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_41=2.3606
+  sky130_fd_pr__nfet_01v8__u0_diff_41=-0.007813
+  sky130_fd_pr__nfet_01v8__ags_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_41=0.023244
+  sky130_fd_pr__nfet_01v8__ua_diff_41=3.3007e-11
*
* sky130_fd_pr__nfet_01v8, Bin 042, W = 0.42, L = 0.5
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__ua_diff_42=1.0402e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_42=1.7881e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_42=0.0010375
+  sky130_fd_pr__nfet_01v8__a0_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_42=12469.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_42=-0.025797
+  sky130_fd_pr__nfet_01v8__pdits_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_42=3.4771e-7
+  sky130_fd_pr__nfet_01v8__voff_diff_42=-0.16534
+  sky130_fd_pr__nfet_01v8__b1_diff_42=5.442e-9
+  sky130_fd_pr__nfet_01v8__pditsd_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_42=0.59804
+  sky130_fd_pr__nfet_01v8__u0_diff_42=-0.0033999
+  sky130_fd_pr__nfet_01v8__ags_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_42=0.0031941
*
* sky130_fd_pr__nfet_01v8, Bin 043, W = 0.55, L = 1.0
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__ags_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_43=0.0060878
+  sky130_fd_pr__nfet_01v8__ua_diff_43=4.7217e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_43=2.7907e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_43=0.0008979
+  sky130_fd_pr__nfet_01v8__a0_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_43=-0.0084492
+  sky130_fd_pr__nfet_01v8__pdits_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_43=2.5069e-7
+  sky130_fd_pr__nfet_01v8__voff_diff_43=-0.16319
+  sky130_fd_pr__nfet_01v8__b1_diff_43=1.5641e-8
+  sky130_fd_pr__nfet_01v8__pditsd_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_43=0.89794
+  sky130_fd_pr__nfet_01v8__u0_diff_43=-0.00060264
*
* sky130_fd_pr__nfet_01v8, Bin 044, W = 0.55, L = 2.0
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__pclm_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_44=0.94421
+  sky130_fd_pr__nfet_01v8__u0_diff_44=-0.0055055
+  sky130_fd_pr__nfet_01v8__ags_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_44=-0.0069084
+  sky130_fd_pr__nfet_01v8__ua_diff_44=2.0545e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_44=-2.3455e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_44=0.00088634
+  sky130_fd_pr__nfet_01v8__a0_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_44=-0.0029039
+  sky130_fd_pr__nfet_01v8__pdits_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_44=1.322e-7
+  sky130_fd_pr__nfet_01v8__voff_diff_44=-0.18813
+  sky130_fd_pr__nfet_01v8__b1_diff_44=3.4191e-8
+  sky130_fd_pr__nfet_01v8__pditsd_diff_44=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 045, W = 0.55, L = 4.0
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__pditsd_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_45=0.76721
+  sky130_fd_pr__nfet_01v8__u0_diff_45=-0.0034722
+  sky130_fd_pr__nfet_01v8__ags_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_45=-0.00094003
+  sky130_fd_pr__nfet_01v8__ua_diff_45=1.2951e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_45=-3.0424e-20
+  sky130_fd_pr__nfet_01v8__tvoff_diff_45=0.0021067
+  sky130_fd_pr__nfet_01v8__a0_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_45=-0.0029546
+  sky130_fd_pr__nfet_01v8__pdits_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_45=1.1102e-7
+  sky130_fd_pr__nfet_01v8__voff_diff_45=-0.20011
+  sky130_fd_pr__nfet_01v8__b1_diff_45=4.3136e-8
*
* sky130_fd_pr__nfet_01v8, Bin 046, W = 0.55, L = 8.0
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__pdits_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_46=-0.21928
+  sky130_fd_pr__nfet_01v8__b1_diff_46=2.1477e-8
+  sky130_fd_pr__nfet_01v8__pditsd_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_46=0.93312
+  sky130_fd_pr__nfet_01v8__u0_diff_46=-0.0014405
+  sky130_fd_pr__nfet_01v8__ags_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_46=-0.00060464
+  sky130_fd_pr__nfet_01v8__ua_diff_46=6.9653e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_46=1.879e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_46=0.0039673
+  sky130_fd_pr__nfet_01v8__a0_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_46=0.0050482
+  sky130_fd_pr__nfet_01v8__b0_diff_46=7.4684e-8
*
* sky130_fd_pr__nfet_01v8, Bin 047, W = 0.55, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__b0_diff_47=4.5808e-7
+  sky130_fd_pr__nfet_01v8__pdits_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_47=-0.096863
+  sky130_fd_pr__nfet_01v8__b1_diff_47=1.6807e-8
+  sky130_fd_pr__nfet_01v8__pditsd_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_47=-0.18196
+  sky130_fd_pr__nfet_01v8__u0_diff_47=-0.0077831
+  sky130_fd_pr__nfet_01v8__ags_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_47=0.055331
+  sky130_fd_pr__nfet_01v8__ua_diff_47=2.0e-10
+  sky130_fd_pr__nfet_01v8__eta0_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_47=-2.8249e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_47=0.00042973
+  sky130_fd_pr__nfet_01v8__a0_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_47=-59771.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_47=-0.19041
*
* sky130_fd_pr__nfet_01v8, Bin 048, W = 0.55, L = 0.5
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__kt1_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_48=-51400.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_48=-0.029427
+  sky130_fd_pr__nfet_01v8__b0_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_48=-0.17394
+  sky130_fd_pr__nfet_01v8__b1_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_48=0.90238
+  sky130_fd_pr__nfet_01v8__u0_diff_48=-0.00080565
+  sky130_fd_pr__nfet_01v8__ags_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_48=-0.0017978
+  sky130_fd_pr__nfet_01v8__ua_diff_48=1.7994e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_48=2.3756e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_48=0.0012794
+  sky130_fd_pr__nfet_01v8__a0_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_48=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 049, W = 0.64, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__a0_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_49=-47316.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_49=-0.12544
+  sky130_fd_pr__nfet_01v8__b0_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_49=-0.10895
+  sky130_fd_pr__nfet_01v8__b1_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_49=0.34841
+  sky130_fd_pr__nfet_01v8__u0_diff_49=-0.0059627
+  sky130_fd_pr__nfet_01v8__ags_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_49=0.061234
+  sky130_fd_pr__nfet_01v8__ua_diff_49=7.3072e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_49=1.5828e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_49=0.00071499
*
* sky130_fd_pr__nfet_01v8, Bin 050, W = 0.84, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__tvoff_diff_50=0.00051568
+  sky130_fd_pr__nfet_01v8__a0_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_50=-43976.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_50=-0.15083
+  sky130_fd_pr__nfet_01v8__pdits_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_50=5.7064e-7
+  sky130_fd_pr__nfet_01v8__voff_diff_50=-0.09516
+  sky130_fd_pr__nfet_01v8__b1_diff_50=-8.1551e-10
+  sky130_fd_pr__nfet_01v8__pditsd_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_50=0.13758
+  sky130_fd_pr__nfet_01v8__u0_diff_50=-0.0075524
+  sky130_fd_pr__nfet_01v8__ags_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_50=0.058891
+  sky130_fd_pr__nfet_01v8__ua_diff_50=3.0207e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_50=1.4434e-20
*
* sky130_fd_pr__nfet_01v8, Bin 051, W = 0.74, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__tvoff_diff_51=0.00060223
+  sky130_fd_pr__nfet_01v8__rdsw_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_51=-49908.81969071
+  sky130_fd_pr__nfet_01v8__kt1_diff_51=6.07518e-5
+  sky130_fd_pr__nfet_01v8__vth0_diff_51=-0.13485178
+  sky130_fd_pr__nfet_01v8__pdits_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_51=3.22831e-7
+  sky130_fd_pr__nfet_01v8__b1_diff_51=-4.61362e-10
+  sky130_fd_pr__nfet_01v8__voff_diff_51=-0.10114852
+  sky130_fd_pr__nfet_01v8__pditsd_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_51=0.00033347
+  sky130_fd_pr__nfet_01v8__u0_diff_51=-0.00405443
+  sky130_fd_pr__nfet_01v8__nfactor_diff_51=-0.15343144
+  sky130_fd_pr__nfet_01v8__keta_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_51=0.05766859
+  sky130_fd_pr__nfet_01v8__ua_diff_51=3.78254e-11
+  sky130_fd_pr__nfet_01v8__ub_diff_51=1.35715e-19
+  sky130_fd_pr__nfet_01v8__eta0_diff_51=-3.00454e-14
*
* sky130_fd_pr__nfet_01v8, Bin 052, W = 0.36, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__ub_diff_52=4.16095e-19
+  sky130_fd_pr__nfet_01v8__eta0_diff_52=3.2537e-5
+  sky130_fd_pr__nfet_01v8__tvoff_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_52=-65067.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_52=-0.045241
+  sky130_fd_pr__nfet_01v8__vth0_diff_52=-0.19181
+  sky130_fd_pr__nfet_01v8__pdits_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_52=-7.39989e-7
+  sky130_fd_pr__nfet_01v8__b1_diff_52=2.7011e-8
+  sky130_fd_pr__nfet_01v8__voff_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_52=0.00091873
+  sky130_fd_pr__nfet_01v8__u0_diff_52=-0.0083504
+  sky130_fd_pr__nfet_01v8__nfactor_diff_52=0.27572
+  sky130_fd_pr__nfet_01v8__keta_diff_52=0.00306555
+  sky130_fd_pr__nfet_01v8__ags_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_52=0.020341
+  sky130_fd_pr__nfet_01v8__ua_diff_52=-4.02468e-11
*
* sky130_fd_pr__nfet_01v8, Bin 053, W = 0.39, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__ua_diff_53=-4.99625e-12
+  sky130_fd_pr__nfet_01v8__ub_diff_53=3.05799e-19
+  sky130_fd_pr__nfet_01v8__eta0_diff_53=1.15988e-5
+  sky130_fd_pr__nfet_01v8__tvoff_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_53=-59191.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_53=-0.053893
+  sky130_fd_pr__nfet_01v8__vth0_diff_53=-0.19305
+  sky130_fd_pr__nfet_01v8__pdits_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_53=-4.77112e-7
+  sky130_fd_pr__nfet_01v8__b1_diff_53=2.47721e-8
+  sky130_fd_pr__nfet_01v8__voff_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_53=0.00032751
+  sky130_fd_pr__nfet_01v8__u0_diff_53=-0.0072906
+  sky130_fd_pr__nfet_01v8__nfactor_diff_53=0.36174
+  sky130_fd_pr__nfet_01v8__keta_diff_53=0.0010928
+  sky130_fd_pr__nfet_01v8__ags_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_53=0.022274
*
* sky130_fd_pr__nfet_01v8, Bin 054, W = 0.52, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__keta_diff_54=-0.00037717
+  sky130_fd_pr__nfet_01v8__ags_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_54=0.029985
+  sky130_fd_pr__nfet_01v8__ua_diff_54=1.04128e-10
+  sky130_fd_pr__nfet_01v8__ub_diff_54=-6.43431e-20
+  sky130_fd_pr__nfet_01v8__eta0_diff_54=-4.00316e-6
+  sky130_fd_pr__nfet_01v8__tvoff_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_54=-49054.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_54=-0.081672
+  sky130_fd_pr__nfet_01v8__vth0_diff_54=-0.20111
+  sky130_fd_pr__nfet_01v8__pdits_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_54=3.24896e-7
+  sky130_fd_pr__nfet_01v8__b1_diff_54=1.79413e-8
+  sky130_fd_pr__nfet_01v8__voff_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_54=-0.00011304
+  sky130_fd_pr__nfet_01v8__u0_diff_54=-0.00048232
+  sky130_fd_pr__nfet_01v8__nfactor_diff_54=0.35204
*
* sky130_fd_pr__nfet_01v8, Bin 055, W = 0.54, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__pclm_diff_55=-4.18441e-5
+  sky130_fd_pr__nfet_01v8__u0_diff_55=-0.00096228
+  sky130_fd_pr__nfet_01v8__nfactor_diff_55=0.18786
+  sky130_fd_pr__nfet_01v8__keta_diff_55=-0.00013962
+  sky130_fd_pr__nfet_01v8__ags_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_55=0.031175
+  sky130_fd_pr__nfet_01v8__ua_diff_55=1.16564e-10
+  sky130_fd_pr__nfet_01v8__ub_diff_55=-1.09034e-19
+  sky130_fd_pr__nfet_01v8__eta0_diff_55=-1.48189e-6
+  sky130_fd_pr__nfet_01v8__tvoff_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_55=-47873.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_55=-0.12696
+  sky130_fd_pr__nfet_01v8__vth0_diff_55=-0.19431
+  sky130_fd_pr__nfet_01v8__pdits_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_55=4.15269e-7
+  sky130_fd_pr__nfet_01v8__b1_diff_55=1.71716e-8
+  sky130_fd_pr__nfet_01v8__voff_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_55=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 056, W = 0.58, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__pditsd_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_56=-7.83128e-5
+  sky130_fd_pr__nfet_01v8__u0_diff_56=0.00065384
+  sky130_fd_pr__nfet_01v8__nfactor_diff_56=0.20262
+  sky130_fd_pr__nfet_01v8__keta_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_56=0.030661
+  sky130_fd_pr__nfet_01v8__ua_diff_56=8.51462e-11
+  sky130_fd_pr__nfet_01v8__ub_diff_56=4.16055e-20
+  sky130_fd_pr__nfet_01v8__eta0_diff_56=2.77352e-6
+  sky130_fd_pr__nfet_01v8__tvoff_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_56=-48118.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_56=-0.13565
+  sky130_fd_pr__nfet_01v8__vth0_diff_56=-0.18869
+  sky130_fd_pr__nfet_01v8__pdits_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_56=2.90133e-7
+  sky130_fd_pr__nfet_01v8__b1_diff_56=1.0645e-8
+  sky130_fd_pr__nfet_01v8__voff_diff_56=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 057, W = 0.6, L = 0.15
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__pdits_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_57=6.86799e-9
+  sky130_fd_pr__nfet_01v8__voff_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_57=-8.11826e-5
+  sky130_fd_pr__nfet_01v8__u0_diff_57=0.001579
+  sky130_fd_pr__nfet_01v8__nfactor_diff_57=0.10358
+  sky130_fd_pr__nfet_01v8__keta_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_57=0.030486
+  sky130_fd_pr__nfet_01v8__ua_diff_57=6.22602e-11
+  sky130_fd_pr__nfet_01v8__ub_diff_57=1.46466e-19
+  sky130_fd_pr__nfet_01v8__eta0_diff_57=2.87515e-6
+  sky130_fd_pr__nfet_01v8__tvoff_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_57=-49294.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_57=-0.17672
+  sky130_fd_pr__nfet_01v8__vth0_diff_57=-0.18333
+  sky130_fd_pr__nfet_01v8__b0_diff_57=1.87189e-7
*
* sky130_fd_pr__nfet_01v8, Bin 058, W = 0.61, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__b0_diff_58=1.38166e-7
+  sky130_fd_pr__nfet_01v8__pdits_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_58=5.06931e-9
+  sky130_fd_pr__nfet_01v8__voff_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_58=-7.0636e-5
+  sky130_fd_pr__nfet_01v8__u0_diff_58=0.0016663
+  sky130_fd_pr__nfet_01v8__nfactor_diff_58=0.14442
+  sky130_fd_pr__nfet_01v8__keta_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_58=0.03038
+  sky130_fd_pr__nfet_01v8__ua_diff_58=5.13586e-11
+  sky130_fd_pr__nfet_01v8__ub_diff_58=1.96251e-19
+  sky130_fd_pr__nfet_01v8__eta0_diff_58=2.50164e-6
+  sky130_fd_pr__nfet_01v8__tvoff_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_58=-49772.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_58=-0.1688
+  sky130_fd_pr__nfet_01v8__vth0_diff_58=-0.18189
*
* sky130_fd_pr__nfet_01v8, Bin 059, W = 0.65, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__kt1_diff_59=-0.17526
+  sky130_fd_pr__nfet_01v8__vsat_diff_59=-42486.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_59=-0.17876
+  sky130_fd_pr__nfet_01v8__b0_diff_59=3.66155e-8
+  sky130_fd_pr__nfet_01v8__pdits_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_59=-5.23278e-11
+  sky130_fd_pr__nfet_01v8__voff_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_59=8.25295e-5
+  sky130_fd_pr__nfet_01v8__u0_diff_59=0.0016984
+  sky130_fd_pr__nfet_01v8__nfactor_diff_59=0.14425
+  sky130_fd_pr__nfet_01v8__keta_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_59=0.0299
+  sky130_fd_pr__nfet_01v8__ua_diff_59=2.10287e-11
+  sky130_fd_pr__nfet_01v8__ub_diff_59=3.16657e-19
+  sky130_fd_pr__nfet_01v8__eta0_diff_59=-4.84694e-17
+  sky130_fd_pr__nfet_01v8__tvoff_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_59=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 060, W = 0.65, L = 0.18
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__vsat_diff_60=-41425.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_60=-0.18935
+  sky130_fd_pr__nfet_01v8__vth0_diff_60=-0.11919
+  sky130_fd_pr__nfet_01v8__pdits_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_60=3.66155e-8
+  sky130_fd_pr__nfet_01v8__voff_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_60=-5.23278e-11
+  sky130_fd_pr__nfet_01v8__pditsd_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_60=8.25291e-5
+  sky130_fd_pr__nfet_01v8__u0_diff_60=0.00078095
+  sky130_fd_pr__nfet_01v8__nfactor_diff_60=0.74631
+  sky130_fd_pr__nfet_01v8__keta_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_60=0.012547
+  sky130_fd_pr__nfet_01v8__ua_diff_60=2.10287e-11
+  sky130_fd_pr__nfet_01v8__ub_diff_60=3.16657e-19
+  sky130_fd_pr__nfet_01v8__eta0_diff_60=-2.39546e-11
+  sky130_fd_pr__nfet_01v8__tvoff_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_60=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 061, W = 0.65, L = 0.25
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__tvoff_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_61=-37582.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_61=-0.16559
+  sky130_fd_pr__nfet_01v8__vth0_diff_61=-0.065342
+  sky130_fd_pr__nfet_01v8__pdits_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_61=0.0030431
+  sky130_fd_pr__nfet_01v8__nfactor_diff_61=1.9071
+  sky130_fd_pr__nfet_01v8__keta_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_61=0.0058357
+  sky130_fd_pr__nfet_01v8__ua_diff_61=-9.108e-12
+  sky130_fd_pr__nfet_01v8__ub_diff_61=4.60449e-19
+  sky130_fd_pr__nfet_01v8__eta0_diff_61=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 062, W = 0.65, L = 0.5
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__tvoff_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_62=-49521.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_62=-0.37856
+  sky130_fd_pr__nfet_01v8__vth0_diff_62=-0.059145
+  sky130_fd_pr__nfet_01v8__pdits_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_62=5.45502e-17
+  sky130_fd_pr__nfet_01v8__b1_diff_62=-2.18149e-18
+  sky130_fd_pr__nfet_01v8__voff_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_62=0.0014459
+  sky130_fd_pr__nfet_01v8__nfactor_diff_62=1.928
+  sky130_fd_pr__nfet_01v8__keta_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_62=-0.0023861
+  sky130_fd_pr__nfet_01v8__ua_diff_62=2.9602e-12
+  sky130_fd_pr__nfet_01v8__ub_diff_62=2.5142e-19
+  sky130_fd_pr__nfet_01v8__eta0_diff_62=0.0
.include "sky130_fd_pr__nfet_01v8.pm3.spice"
