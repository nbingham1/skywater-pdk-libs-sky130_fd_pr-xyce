* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param sky130_fd_pr__special_nfet_pass__tox_slope_spectre=0.0
.param sky130_fd_pr__special_nfet_pass__vth0_slope_spectre=0.0
.param sky130_fd_pr__special_nfet_pass__voff_slope_spectre=0.0
.param sky130_fd_pr__special_nfet_pass__nfactor_slope_spectre=0.0
* statistics {
*   process {
*   }
*   mismatch {
*     vary sky130_fd_pr__special_nfet_pass__tox_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__special_nfet_pass__vth0_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__special_nfet_pass__voff_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__special_nfet_pass__nfactor_slope_spectre dist=gauss std = 1.0
*   }
* }
.subckt sky130_fd_pr__special_nfet_pass d g s b
.param l=1 w=1 ad=0 as=0 pd=0 ps=0 nrd=0 nrs=0 mult=1 sa=0 sb=0 sd=0.0
msky130_fd_pr__special_nfet_pass d g s b sky130_fd_pr__special_nfet_pass__model l={l} w={w} ad={ad} as={as} pd={pd} ps={ps} nrd={nrd} nrs={nrs}
.model sky130_fd_pr__special_nfet_pass__model.0 nmos
+  lmin=7.5e-08 lmax=1.505e-007 wmin=1.395e-007 wmax=1.405e-7
+  level=49.0
+  tnom=30.0
+  version=3.2
+  tox={4.148e-009*sky130_fd_pr__special_nfet_pass__tox_mult+sky130_fd_pr__special_nfet_pass__tox_slope_spectre*(4.148e-009*sky130_fd_pr__special_nfet_pass__tox_mult*(sky130_fd_pr__special_nfet_pass__tox_slope/sqrt(l*w*mult)))}
+  toxm=4.148e-9
+  xj=1.2e-7
+  nch=1.12471e+18
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint={0+sky130_fd_pr__special_nfet_pass__lint_diff}
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint={0+sky130_fd_pr__special_nfet_pass__wint_diff}
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  mobmod=1.0
+  binunit=2.0
+  dwg=0.0
+  dwb=0.0
* Diode Parameters
+  ldif=0.0
+  hdif=0.0
+  rd=0.0
+  rs=0.0
+  rsc=0.0
+  rdc=0.0
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.65009+sky130_fd_pr__special_nfet_pass__vth0_diff_0+sky130_fd_pr__special_nfet_pass__vth0_slope_spectre*(sky130_fd_pr__special_nfet_pass__vth0_slope/sqrt(w*l*mult))}
+  k1=0.53066
+  k2={-0.12745+sky130_fd_pr__special_nfet_pass__k2_diff_0}
+  k3={0+sky130_fd_pr__special_nfet_pass__k3_diff}
+  dvt0={0+sky130_fd_pr__special_nfet_pass__dvt0_diff}
+  dvt1=0.53
+  dvt2=0.0
+  dvt0w=0.0
+  dvt1w=10100.0
+  dvt2w=0.0
+  nlx=0.0
+  w0=1.0e-6
+  k3b=0.0
+  ngate=1.0e+23
+  vfb=-0.9693
* Mobility Parameters
+  vsat={101250+sky130_fd_pr__special_nfet_pass__vsat_diff_0}
+  ua=-1.9925e-9
+  ub=1.9307e-18
+  uc=4.5872e-11
+  rdsw={103.2113+sky130_fd_pr__special_nfet_pass__rdsw_diff_0}
+  prwb=0.3
+  prwg=0.2
+  wr=1.0
+  u0={0.01592+sky130_fd_pr__special_nfet_pass__u0_diff_0}
+  a0=1.0
+  keta=-0.061906
+  a1=0.0
+  a2=1.0
+  ags=0.5115
+  b0=0.0
+  b1=0.0
* Subthreshold Current Parameters
+  voff={-0.15507+sky130_fd_pr__special_nfet_pass__voff_diff_0+sky130_fd_pr__special_nfet_pass__voff_slope_spectre*(sky130_fd_pr__special_nfet_pass__voff_slope/sqrt(w*l*mult))}
+  nfactor={1.7935+sky130_fd_pr__special_nfet_pass__nfactor_diff_0+sky130_fd_pr__special_nfet_pass__nfactor_slope_spectre*(sky130_fd_pr__special_nfet_pass__nfactor_slope/sqrt(w*l*mult))}
+  cit={0+sky130_fd_pr__special_nfet_pass__cit_diff}
+  cdsc={0+sky130_fd_pr__special_nfet_pass__cdsc_diff}
+  cdscb={0+sky130_fd_pr__special_nfet_pass__cdscb_diff}
+  cdscd={0+sky130_fd_pr__special_nfet_pass__cdscd_diff}
+  eta0=0.1168
+  etab=0.00804
+  dsub=0.5
* Rout Parameters
+  pclm=0.93451
+  pdiblc1=0.0
+  pdiblc2=0.035291
+  pdiblcb=-0.15462
+  drout=0.5
+  pscbe1=7.8166e+8
+  pscbe2=1.0e-20
+  pvag=0.0
+  delta=0.0104
+  alpha0=0.00064059
+  alpha1=0.0
+  beta0=26.6
* Temperature Effects Parameters
+  kt1={-0.245+sky130_fd_pr__special_nfet_pass__kt1_diff_0}
+  kt2={-0.01458+sky130_fd_pr__special_nfet_pass__kt2_diff}
+  at=25430.0
+  ute=-1.1259
+  ua1=3.7209e-10
+  ub1=-1.3557e-19
+  uc1=-2.31e-12
+  kt1l={0+sky130_fd_pr__special_nfet_pass__kt1l_diff}
+  prt=0.0
* Capacitance Parameters
+  cj={0.0013459*sky130_fd_pr__special_nfet_pass__ajunction_mult}
+  mj=0.44
+  pb=0.729
+  cjsw={3.6001e-011*sky130_fd_pr__special_nfet_pass__pjunction_mult}
+  mjsw=0.0009
+  pbsw=0.2
+  cjswg={2.3347e-010*sky130_fd_pr__special_nfet_pass__pjunction_mult}
+  mjswg=0.8000
+  pbswg=0.95578
+  tpb=0.0012287
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.000792
+  tcjsw=1.0e-5
+  tcjswg=0.0
+  js=0.0027500000000000003
+  jsw=6.0e-10
+  nj=1.2928
+  xti=2.0
+  cgdo={3.2e-010*sky130_fd_pr__special_nfet_pass__overlap_mult}
+  cgso={3.2e-010*sky130_fd_pr__special_nfet_pass__overlap_mult}
+  cgbo=1.0e-13
+  capmod=3.0
+  nqsmod=0.0
+  elm=0.0
+  xpart=0.0
+  cgsl={0*sky130_fd_pr__special_nfet_pass__overlap_mult}
+  cgdl={0*sky130_fd_pr__special_nfet_pass__overlap_mult}
+  ckappa=0.6
+  cf=1.4067e-12
+  clc=1.0e-7
+  cle=0.6
+  dlc={1.8739e-008+sky130_fd_pr__special_nfet_pass__dlc_diff+sky130_fd_pr__special_nfet_pass__dlc_rotweak}
+  dwc={0+sky130_fd_pr__special_nfet_pass__dwc_diff}
+  vfbcv=-1.0
+  acde=0.4
+  moin=6.9
+  noff=3.621
+  voffcv=-0.1372
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
+  noimod=2.0
+  noia={1.1737146E+41*1.6e-21}
+  noib={3.2036721E+25*1.6e-21}
+  noic={-3.7339643E+08*1.6e-21}
+  em=4.1000000e+7
+  ef=0.8439365
.ends sky130_fd_pr__special_nfet_pass
