* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 52
.param
+  sky130_fd_pr__pfet_01v8__toxe_mult=0.948
+  sky130_fd_pr__pfet_01v8__rshp_mult=1.0
+  sky130_fd_pr__pfet_01v8__overlap_mult=0.95436
+  sky130_fd_pr__pfet_01v8__ajunction_mult=0.90161
+  sky130_fd_pr__pfet_01v8__pjunction_mult=0.90587
+  sky130_fd_pr__pfet_01v8__lint_diff=1.7325e-8
+  sky130_fd_pr__pfet_01v8__wint_diff=-3.2175e-8
+  sky130_fd_pr__pfet_01v8__dlc_diff=1.7325e-8
+  sky130_fd_pr__pfet_01v8__dwc_diff=-3.2175e-8
*
* sky130_fd_pr__pfet_01v8, Bin 000, W = 1.26, L = 0.15
* -----------------------------------
+  sky130_fd_pr__pfet_01v8__agidl_diff_0=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_0=3.9271
+  sky130_fd_pr__pfet_01v8__vsat_diff_0=-12590.0
+  sky130_fd_pr__pfet_01v8__a0_diff_0=0.0
+  sky130_fd_pr__pfet_01v8__pdits_diff_0=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_0=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_0=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_0=-0.046667
+  sky130_fd_pr__pfet_01v8__eta0_diff_0=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_0=-2.3326e-12
+  sky130_fd_pr__pfet_01v8__keta_diff_0=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_0=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_0=0.0045512
+  sky130_fd_pr__pfet_01v8__vth0_diff_0=-0.060116
+  sky130_fd_pr__pfet_01v8__pditsd_diff_0=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_0=0.00066699
+  sky130_fd_pr__pfet_01v8__b1_diff_0=0.0
+  sky130_fd_pr__pfet_01v8__cgidl_diff_0=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_0=0.00014246
+  sky130_fd_pr__pfet_01v8__voff_diff_0=-0.20341
+  sky130_fd_pr__pfet_01v8__ags_diff_0=0.0
+  sky130_fd_pr__pfet_01v8__bgidl_diff_0=0.0
+  sky130_fd_pr__pfet_01v8__ub_diff_0=4.1498e-19
*
* sky130_fd_pr__pfet_01v8, Bin 001, W = 1.68, L = 0.15
* -----------------------------------
+  sky130_fd_pr__pfet_01v8__bgidl_diff_1=0.0
+  sky130_fd_pr__pfet_01v8__ub_diff_1=3.0525e-19
+  sky130_fd_pr__pfet_01v8__agidl_diff_1=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_1=1.747
+  sky130_fd_pr__pfet_01v8__vsat_diff_1=-16150.0
+  sky130_fd_pr__pfet_01v8__a0_diff_1=0.0
+  sky130_fd_pr__pfet_01v8__pdits_diff_1=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_1=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_1=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_1=0.26882
+  sky130_fd_pr__pfet_01v8__eta0_diff_1=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_1=-3.8211e-11
+  sky130_fd_pr__pfet_01v8__keta_diff_1=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_1=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_1=4.4689e-5
+  sky130_fd_pr__pfet_01v8__vth0_diff_1=-0.12401
+  sky130_fd_pr__pfet_01v8__pditsd_diff_1=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_1=0.0003403
+  sky130_fd_pr__pfet_01v8__b1_diff_1=0.0
+  sky130_fd_pr__pfet_01v8__cgidl_diff_1=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_1=0.00016892
+  sky130_fd_pr__pfet_01v8__voff_diff_1=-0.20951
+  sky130_fd_pr__pfet_01v8__ags_diff_1=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 002, W = 1.0, L = 1.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__cgidl_diff_2=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_2=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_2=-0.38202
+  sky130_fd_pr__pfet_01v8__ags_diff_2=0.090628
+  sky130_fd_pr__pfet_01v8__bgidl_diff_2=0.0
+  sky130_fd_pr__pfet_01v8__ub_diff_2=5.467e-19
+  sky130_fd_pr__pfet_01v8__agidl_diff_2=3.5884e-10
+  sky130_fd_pr__pfet_01v8__nfactor_diff_2=2.341
+  sky130_fd_pr__pfet_01v8__vsat_diff_2=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_2=-0.080923
+  sky130_fd_pr__pfet_01v8__pdits_diff_2=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_2=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_2=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_2=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_2=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_2=3.5075e-12
+  sky130_fd_pr__pfet_01v8__keta_diff_2=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_2=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_2=-0.0075788
+  sky130_fd_pr__pfet_01v8__vth0_diff_2=0.0086043
+  sky130_fd_pr__pfet_01v8__pditsd_diff_2=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_2=0.0024412
+  sky130_fd_pr__pfet_01v8__b1_diff_2=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 003, W = 1.0, L = 2.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__b1_diff_3=0.0
+  sky130_fd_pr__pfet_01v8__cgidl_diff_3=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_3=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_3=-0.49539
+  sky130_fd_pr__pfet_01v8__ags_diff_3=0.031106
+  sky130_fd_pr__pfet_01v8__bgidl_diff_3=0.0
+  sky130_fd_pr__pfet_01v8__ub_diff_3=6.3506e-19
+  sky130_fd_pr__pfet_01v8__nfactor_diff_3=3.1461
+  sky130_fd_pr__pfet_01v8__vsat_diff_3=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_3=3.3327e-11
+  sky130_fd_pr__pfet_01v8__a0_diff_3=-0.033883
+  sky130_fd_pr__pfet_01v8__pdits_diff_3=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_3=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_3=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_3=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_3=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_3=-2.4052e-12
+  sky130_fd_pr__pfet_01v8__keta_diff_3=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_3=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_3=-0.012185
+  sky130_fd_pr__pfet_01v8__vth0_diff_3=0.012973
+  sky130_fd_pr__pfet_01v8__pditsd_diff_3=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_3=0.0029724
*
* sky130_fd_pr__pfet_01v8, Bin 004, W = 1.0, L = 4.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__pditsd_diff_4=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_4=0.0030608
+  sky130_fd_pr__pfet_01v8__vth0_diff_4=-0.0038108
+  sky130_fd_pr__pfet_01v8__b1_diff_4=0.0
+  sky130_fd_pr__pfet_01v8__cgidl_diff_4=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_4=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_4=-0.5
+  sky130_fd_pr__pfet_01v8__ags_diff_4=0.045074
+  sky130_fd_pr__pfet_01v8__ub_diff_4=6.1783e-19
+  sky130_fd_pr__pfet_01v8__bgidl_diff_4=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_4=3.8259
+  sky130_fd_pr__pfet_01v8__vsat_diff_4=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_4=4.5377e-10
+  sky130_fd_pr__pfet_01v8__a0_diff_4=-0.044369
+  sky130_fd_pr__pfet_01v8__pdits_diff_4=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_4=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_4=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_4=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_4=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_4=3.5061e-13
+  sky130_fd_pr__pfet_01v8__keta_diff_4=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_4=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_4=-0.013265
*
* sky130_fd_pr__pfet_01v8, Bin 005, W = 1.0, L = 8.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__keta_diff_5=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_5=-0.015073
+  sky130_fd_pr__pfet_01v8__pditsd_diff_5=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_5=0.0025277
+  sky130_fd_pr__pfet_01v8__vth0_diff_5=-0.019932
+  sky130_fd_pr__pfet_01v8__b1_diff_5=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_5=-0.51622
+  sky130_fd_pr__pfet_01v8__cgidl_diff_5=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_5=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_5=0.085945
+  sky130_fd_pr__pfet_01v8__ub_diff_5=5.1769e-19
+  sky130_fd_pr__pfet_01v8__bgidl_diff_5=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_5=4.4585
+  sky130_fd_pr__pfet_01v8__vsat_diff_5=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_5=2.8514e-10
+  sky130_fd_pr__pfet_01v8__a0_diff_5=-0.079147
+  sky130_fd_pr__pfet_01v8__pdits_diff_5=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_5=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_5=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_5=-0.25
+  sky130_fd_pr__pfet_01v8__eta0_diff_5=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_5=-6.2498e-12
+  sky130_fd_pr__pfet_01v8__rdsw_diff_5=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 006, W = 1.0, L = 0.15
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__rdsw_diff_6=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_6=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_6=0.025127
+  sky130_fd_pr__pfet_01v8__pditsd_diff_6=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_6=-0.00052537
+  sky130_fd_pr__pfet_01v8__vth0_diff_6=-0.10378
+  sky130_fd_pr__pfet_01v8__b1_diff_6=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_6=-0.057734
+  sky130_fd_pr__pfet_01v8__cgidl_diff_6=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_6=-2.2501e-5
+  sky130_fd_pr__pfet_01v8__ags_diff_6=0.0
+  sky130_fd_pr__pfet_01v8__ub_diff_6=7.825e-19
+  sky130_fd_pr__pfet_01v8__bgidl_diff_6=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_6=1.4849
+  sky130_fd_pr__pfet_01v8__vsat_diff_6=-20000.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_6=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_6=0.0
+  sky130_fd_pr__pfet_01v8__pdits_diff_6=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_6=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_6=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_6=0.024244
+  sky130_fd_pr__pfet_01v8__eta0_diff_6=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_6=-5.0e-10
*
* sky130_fd_pr__pfet_01v8, Bin 007, W = 1.0, L = 0.18
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__kt1_diff_7=0.055183
+  sky130_fd_pr__pfet_01v8__eta0_diff_7=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_7=1.2857e-10
+  sky130_fd_pr__pfet_01v8__rdsw_diff_7=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_7=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_7=-0.00076543
+  sky130_fd_pr__pfet_01v8__pditsd_diff_7=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_7=0.00070488
+  sky130_fd_pr__pfet_01v8__vth0_diff_7=-0.081389
+  sky130_fd_pr__pfet_01v8__b1_diff_7=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_7=-0.045269
+  sky130_fd_pr__pfet_01v8__cgidl_diff_7=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_7=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_7=0.0
+  sky130_fd_pr__pfet_01v8__ub_diff_7=2.2283e-19
+  sky130_fd_pr__pfet_01v8__bgidl_diff_7=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_7=-0.011494
+  sky130_fd_pr__pfet_01v8__vsat_diff_7=-20000.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_7=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_7=0.0
+  sky130_fd_pr__pfet_01v8__pdits_diff_7=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_7=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_7=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 008, W = 1.0, L = 0.25
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__pclm_diff_8=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_8=0.14284
+  sky130_fd_pr__pfet_01v8__eta0_diff_8=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_8=2.7416e-11
+  sky130_fd_pr__pfet_01v8__rdsw_diff_8=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_8=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_8=-0.0021971
+  sky130_fd_pr__pfet_01v8__pditsd_diff_8=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_8=0.00017366
+  sky130_fd_pr__pfet_01v8__vth0_diff_8=-0.00087253
+  sky130_fd_pr__pfet_01v8__b1_diff_8=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_8=-0.20736
+  sky130_fd_pr__pfet_01v8__cgidl_diff_8=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_8=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_8=0.0
+  sky130_fd_pr__pfet_01v8__ub_diff_8=2.9171e-19
+  sky130_fd_pr__pfet_01v8__bgidl_diff_8=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_8=1.1224
+  sky130_fd_pr__pfet_01v8__vsat_diff_8=100000.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_8=-2.1595e-10
+  sky130_fd_pr__pfet_01v8__a0_diff_8=0.0
+  sky130_fd_pr__pfet_01v8__pdits_diff_8=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_8=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 009, W = 1.0, L = 0.5
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__pdits_diff_9=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_9=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_9=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_9=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_9=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_9=1.0972e-12
+  sky130_fd_pr__pfet_01v8__rdsw_diff_9=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_9=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_9=-0.0087514
+  sky130_fd_pr__pfet_01v8__pditsd_diff_9=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_9=0.0011707
+  sky130_fd_pr__pfet_01v8__vth0_diff_9=0.044728
+  sky130_fd_pr__pfet_01v8__b1_diff_9=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_9=-1.0025
+  sky130_fd_pr__pfet_01v8__cgidl_diff_9=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_9=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_9=0.0
+  sky130_fd_pr__pfet_01v8__ub_diff_9=4.4605e-19
+  sky130_fd_pr__pfet_01v8__bgidl_diff_9=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_9=0.41724
+  sky130_fd_pr__pfet_01v8__vsat_diff_9=-3032.7
+  sky130_fd_pr__pfet_01v8__agidl_diff_9=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_9=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 010, W = 2.0, L = 0.15
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__pditsd_diff_10=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_10=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_10=-20000.0
+  sky130_fd_pr__pfet_01v8__u0_diff_10=-0.00070501
+  sky130_fd_pr__pfet_01v8__vth0_diff_10=-0.08634
+  sky130_fd_pr__pfet_01v8__cgidl_diff_10=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_10=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_10=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_10=0.20358
+  sky130_fd_pr__pfet_01v8__pclm_diff_10=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_10=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_10=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_10=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_10=-2.9668e-10
+  sky130_fd_pr__pfet_01v8__bgidl_diff_10=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_10=1.0176
+  sky130_fd_pr__pfet_01v8__ub_diff_10=3.3082e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_10=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_10=-0.00010189
+  sky130_fd_pr__pfet_01v8__ags_diff_10=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_10=0.039771
+  sky130_fd_pr__pfet_01v8__voff_diff_10=-0.10358
+  sky130_fd_pr__pfet_01v8__a0_diff_10=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 011, W = 3.0, L = 1.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__voff_diff_11=-0.37512
+  sky130_fd_pr__pfet_01v8__a0_diff_11=-0.12119
+  sky130_fd_pr__pfet_01v8__pditsd_diff_11=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_11=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_11=27194.0
+  sky130_fd_pr__pfet_01v8__u0_diff_11=0.0018883
+  sky130_fd_pr__pfet_01v8__vth0_diff_11=-0.0031631
+  sky130_fd_pr__pfet_01v8__cgidl_diff_11=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_11=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_11=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_11=3.9344e-6
+  sky130_fd_pr__pfet_01v8__pclm_diff_11=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_11=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_11=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_11=9.2899e-10
+  sky130_fd_pr__pfet_01v8__ua_diff_11=-3.8915e-11
+  sky130_fd_pr__pfet_01v8__bgidl_diff_11=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_11=2.5816
+  sky130_fd_pr__pfet_01v8__ub_diff_11=4.9719e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_11=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_11=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_11=0.098819
+  sky130_fd_pr__pfet_01v8__k2_diff_11=-0.014591
*
* sky130_fd_pr__pfet_01v8, Bin 012, W = 3.0, L = 2.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__pdits_diff_12=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_12=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_12=0.091497
+  sky130_fd_pr__pfet_01v8__k2_diff_12=-0.0081409
+  sky130_fd_pr__pfet_01v8__voff_diff_12=-0.39425
+  sky130_fd_pr__pfet_01v8__a0_diff_12=-0.1016
+  sky130_fd_pr__pfet_01v8__pditsd_diff_12=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_12=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_12=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_12=0.002524
+  sky130_fd_pr__pfet_01v8__vth0_diff_12=-0.0034613
+  sky130_fd_pr__pfet_01v8__cgidl_diff_12=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_12=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_12=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_12=-5.9055e-6
+  sky130_fd_pr__pfet_01v8__pclm_diff_12=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_12=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_12=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_12=8.6561e-11
+  sky130_fd_pr__pfet_01v8__ua_diff_12=-4.5581e-12
+  sky130_fd_pr__pfet_01v8__bgidl_diff_12=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_12=2.7379
+  sky130_fd_pr__pfet_01v8__ub_diff_12=5.4069e-19
*
* sky130_fd_pr__pfet_01v8, Bin 013, W = 3.0, L = 4.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__bgidl_diff_13=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_13=4.0
+  sky130_fd_pr__pfet_01v8__ub_diff_13=5.6615e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_13=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_13=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_13=0.066928
+  sky130_fd_pr__pfet_01v8__k2_diff_13=-0.0062466
+  sky130_fd_pr__pfet_01v8__voff_diff_13=-0.4
+  sky130_fd_pr__pfet_01v8__a0_diff_13=-0.073723
+  sky130_fd_pr__pfet_01v8__eta0_diff_13=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_13=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_13=0.0027737
+  sky130_fd_pr__pfet_01v8__vsat_diff_13=0.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_13=0.001697
+  sky130_fd_pr__pfet_01v8__cgidl_diff_13=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_13=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_13=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_13=-0.12264
+  sky130_fd_pr__pfet_01v8__pclm_diff_13=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_13=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_13=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_13=1.6289e-10
+  sky130_fd_pr__pfet_01v8__ua_diff_13=-3.3779e-12
*
* sky130_fd_pr__pfet_01v8, Bin 014, W = 3.0, L = 8.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__agidl_diff_14=3.1829e-9
+  sky130_fd_pr__pfet_01v8__b1_diff_14=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_14=-3.0908e-12
+  sky130_fd_pr__pfet_01v8__bgidl_diff_14=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_14=4.0
+  sky130_fd_pr__pfet_01v8__ub_diff_14=6.5948e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_14=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_14=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_14=0.048267
+  sky130_fd_pr__pfet_01v8__k2_diff_14=-0.0063904
+  sky130_fd_pr__pfet_01v8__voff_diff_14=-0.4
+  sky130_fd_pr__pfet_01v8__eta0_diff_14=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_14=-0.05886
+  sky130_fd_pr__pfet_01v8__pditsd_diff_14=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_14=0.003279
+  sky130_fd_pr__pfet_01v8__vsat_diff_14=0.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_14=0.0041156
+  sky130_fd_pr__pfet_01v8__cgidl_diff_14=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_14=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_14=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_14=-0.45471
+  sky130_fd_pr__pfet_01v8__pclm_diff_14=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_14=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 015, W = 3.0, L = 0.15
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__b0_diff_15=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_15=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_15=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_15=2.9356e-10
+  sky130_fd_pr__pfet_01v8__bgidl_diff_15=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_15=0.45655
+  sky130_fd_pr__pfet_01v8__ub_diff_15=-5.5818e-20
+  sky130_fd_pr__pfet_01v8__tvoff_diff_15=0.007
+  sky130_fd_pr__pfet_01v8__ags_diff_15=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_15=0.00079783
+  sky130_fd_pr__pfet_01v8__pdits_diff_15=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_15=-0.082195
+  sky130_fd_pr__pfet_01v8__eta0_diff_15=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_15=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_15=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_15=0.0010674
+  sky130_fd_pr__pfet_01v8__vsat_diff_15=-20000.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_15=-0.15768
+  sky130_fd_pr__pfet_01v8__cgidl_diff_15=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_15=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_15=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_15=0.36152
+  sky130_fd_pr__pfet_01v8__pclm_diff_15=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 016, W = 3.0, L = 0.18
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__pclm_diff_16=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_16=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_16=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_16=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_16=2.0851e-11
+  sky130_fd_pr__pfet_01v8__bgidl_diff_16=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_16=0.2935
+  sky130_fd_pr__pfet_01v8__tvoff_diff_16=1.1012e-5
+  sky130_fd_pr__pfet_01v8__ags_diff_16=0.0
+  sky130_fd_pr__pfet_01v8__ub_diff_16=1.946e-19
+  sky130_fd_pr__pfet_01v8__k2_diff_16=0.0030068
+  sky130_fd_pr__pfet_01v8__pdits_diff_16=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_16=-0.10254
+  sky130_fd_pr__pfet_01v8__eta0_diff_16=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_16=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_16=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_16=0.00041253
+  sky130_fd_pr__pfet_01v8__vsat_diff_16=-17517.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_16=-0.07292
+  sky130_fd_pr__pfet_01v8__cgidl_diff_16=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_16=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_16=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_16=-0.0010807
*
* sky130_fd_pr__pfet_01v8, Bin 017, W = 3.0, L = 0.25
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__kt1_diff_17=0.53407
+  sky130_fd_pr__pfet_01v8__pclm_diff_17=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_17=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_17=1.0001e-10
+  sky130_fd_pr__pfet_01v8__b1_diff_17=0.0
+  sky130_fd_pr__pfet_01v8__bgidl_diff_17=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_17=0.83987
+  sky130_fd_pr__pfet_01v8__ua_diff_17=-1.804e-11
+  sky130_fd_pr__pfet_01v8__tvoff_diff_17=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_17=0.0
+  sky130_fd_pr__pfet_01v8__ub_diff_17=2.52e-19
+  sky130_fd_pr__pfet_01v8__k2_diff_17=0.001971
+  sky130_fd_pr__pfet_01v8__pdits_diff_17=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_17=-0.21242
+  sky130_fd_pr__pfet_01v8__eta0_diff_17=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_17=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_17=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_17=-4.6213e-5
+  sky130_fd_pr__pfet_01v8__vsat_diff_17=-17319.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_17=0.04076
+  sky130_fd_pr__pfet_01v8__cgidl_diff_17=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_17=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_17=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 018, W = 3.0, L = 0.5
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__rdsw_diff_18=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_18=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_18=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_18=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_18=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_18=0.0
+  sky130_fd_pr__pfet_01v8__bgidl_diff_18=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_18=0.63675
+  sky130_fd_pr__pfet_01v8__ua_diff_18=1.4339e-11
+  sky130_fd_pr__pfet_01v8__tvoff_diff_18=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_18=0.0
+  sky130_fd_pr__pfet_01v8__ub_diff_18=3.5515e-19
+  sky130_fd_pr__pfet_01v8__k2_diff_18=-0.012538
+  sky130_fd_pr__pfet_01v8__pdits_diff_18=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_18=-1.3476
+  sky130_fd_pr__pfet_01v8__eta0_diff_18=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_18=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_18=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_18=0.0013831
+  sky130_fd_pr__pfet_01v8__vsat_diff_18=15158.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_18=0.01865
+  sky130_fd_pr__pfet_01v8__cgidl_diff_18=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_18=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 019, W = 5.0, L = 1.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__cgidl_diff_19=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_19=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_19=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_19=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_19=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_19=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_19=6.0145e-10
+  sky130_fd_pr__pfet_01v8__b1_diff_19=0.0
+  sky130_fd_pr__pfet_01v8__bgidl_diff_19=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_19=2.3221
+  sky130_fd_pr__pfet_01v8__ua_diff_19=-9.2578e-12
+  sky130_fd_pr__pfet_01v8__tvoff_diff_19=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_19=0.17047
+  sky130_fd_pr__pfet_01v8__ub_diff_19=3.6396e-19
+  sky130_fd_pr__pfet_01v8__k2_diff_19=-0.009739
+  sky130_fd_pr__pfet_01v8__pdits_diff_19=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_19=-0.34631
+  sky130_fd_pr__pfet_01v8__eta0_diff_19=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_19=-0.16939
+  sky130_fd_pr__pfet_01v8__pditsd_diff_19=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_19=0.0015601
+  sky130_fd_pr__pfet_01v8__vsat_diff_19=0.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_19=0.01352
*
* sky130_fd_pr__pfet_01v8, Bin 020, W = 5.0, L = 2.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__u0_diff_20=0.0017436
+  sky130_fd_pr__pfet_01v8__vth0_diff_20=0.0098523
+  sky130_fd_pr__pfet_01v8__cgidl_diff_20=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_20=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_20=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_20=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_20=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_20=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_20=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_20=1.9618e-9
+  sky130_fd_pr__pfet_01v8__ua_diff_20=-2.3869e-12
+  sky130_fd_pr__pfet_01v8__bgidl_diff_20=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_20=2.794
+  sky130_fd_pr__pfet_01v8__ub_diff_20=3.5988e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_20=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_20=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_20=0.040922
+  sky130_fd_pr__pfet_01v8__k2_diff_20=-0.0091133
+  sky130_fd_pr__pfet_01v8__voff_diff_20=-0.38844
+  sky130_fd_pr__pfet_01v8__a0_diff_20=-0.044531
+  sky130_fd_pr__pfet_01v8__pditsd_diff_20=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_20=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_20=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 021, W = 5.0, L = 4.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__pditsd_diff_21=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_21=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_21=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_21=0.0024494
+  sky130_fd_pr__pfet_01v8__vth0_diff_21=0.0088283
+  sky130_fd_pr__pfet_01v8__cgidl_diff_21=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_21=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_21=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_21=-0.073293
+  sky130_fd_pr__pfet_01v8__pclm_diff_21=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_21=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_21=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_21=4.6058e-9
+  sky130_fd_pr__pfet_01v8__ua_diff_21=-4.1623e-12
+  sky130_fd_pr__pfet_01v8__bgidl_diff_21=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_21=4.0
+  sky130_fd_pr__pfet_01v8__ub_diff_21=4.7009e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_21=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_21=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_21=0.049075
+  sky130_fd_pr__pfet_01v8__k2_diff_21=-0.0096588
+  sky130_fd_pr__pfet_01v8__voff_diff_21=-0.4
+  sky130_fd_pr__pfet_01v8__a0_diff_21=-0.059424
*
* sky130_fd_pr__pfet_01v8, Bin 022, W = 5.0, L = 8.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__voff_diff_22=-0.4
+  sky130_fd_pr__pfet_01v8__a0_diff_22=-0.064689
+  sky130_fd_pr__pfet_01v8__pditsd_diff_22=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_22=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_22=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_22=0.0026485
+  sky130_fd_pr__pfet_01v8__vth0_diff_22=0.0030374
+  sky130_fd_pr__pfet_01v8__cgidl_diff_22=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_22=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_22=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_22=-0.42913
+  sky130_fd_pr__pfet_01v8__pclm_diff_22=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_22=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_22=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_22=7.6144e-9
+  sky130_fd_pr__pfet_01v8__ua_diff_22=-2.2073e-12
+  sky130_fd_pr__pfet_01v8__bgidl_diff_22=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_22=4.0
+  sky130_fd_pr__pfet_01v8__ub_diff_22=5.0422e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_22=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_22=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_22=0.039071
+  sky130_fd_pr__pfet_01v8__k2_diff_22=-0.009782
*
* sky130_fd_pr__pfet_01v8, Bin 023, W = 5.0, L = 0.15
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__pdits_diff_23=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_23=0.00061853
+  sky130_fd_pr__pfet_01v8__ags_diff_23=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_23=0.040345
+  sky130_fd_pr__pfet_01v8__voff_diff_23=-0.12462
+  sky130_fd_pr__pfet_01v8__a0_diff_23=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_23=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_23=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_23=-20000.0
+  sky130_fd_pr__pfet_01v8__u0_diff_23=-0.0012
+  sky130_fd_pr__pfet_01v8__vth0_diff_23=-0.096011
+  sky130_fd_pr__pfet_01v8__cgidl_diff_23=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_23=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_23=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_23=0.25038
+  sky130_fd_pr__pfet_01v8__pclm_diff_23=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_23=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_23=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_23=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_23=-4.5385e-10
+  sky130_fd_pr__pfet_01v8__bgidl_diff_23=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_23=0.65407
+  sky130_fd_pr__pfet_01v8__ub_diff_23=4.7501e-19
*
* sky130_fd_pr__pfet_01v8, Bin 024, W = 5.0, L = 0.18
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__bgidl_diff_24=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_24=0.32687
+  sky130_fd_pr__pfet_01v8__ub_diff_24=1.4305e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_24=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_24=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_24=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_24=0.0052883
+  sky130_fd_pr__pfet_01v8__voff_diff_24=-0.11464
+  sky130_fd_pr__pfet_01v8__a0_diff_24=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_24=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_24=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_24=8.3631e-5
+  sky130_fd_pr__pfet_01v8__vsat_diff_24=-4518.1
+  sky130_fd_pr__pfet_01v8__vth0_diff_24=-0.086527
+  sky130_fd_pr__pfet_01v8__cgidl_diff_24=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_24=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_24=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_24=-0.013482
+  sky130_fd_pr__pfet_01v8__pclm_diff_24=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_24=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_24=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_24=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_24=-5.787e-12
*
* sky130_fd_pr__pfet_01v8, Bin 025, W = 5.0, L = 0.25
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__agidl_diff_25=4.1688e-9
+  sky130_fd_pr__pfet_01v8__b1_diff_25=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_25=1.5952e-12
+  sky130_fd_pr__pfet_01v8__bgidl_diff_25=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_25=0.56131
+  sky130_fd_pr__pfet_01v8__ub_diff_25=2.0125e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_25=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_25=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_25=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_25=-0.00017766
+  sky130_fd_pr__pfet_01v8__voff_diff_25=-0.20387
+  sky130_fd_pr__pfet_01v8__eta0_diff_25=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_25=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_25=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_25=0.00043723
+  sky130_fd_pr__pfet_01v8__vsat_diff_25=4287.1
+  sky130_fd_pr__pfet_01v8__vth0_diff_25=-0.046289
+  sky130_fd_pr__pfet_01v8__cgidl_diff_25=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_25=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_25=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_25=-0.018093
+  sky130_fd_pr__pfet_01v8__pclm_diff_25=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_25=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 026, W = 5.0, L = 0.5
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__b0_diff_26=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_26=7.6855e-10
+  sky130_fd_pr__pfet_01v8__b1_diff_26=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_26=2.4056e-11
+  sky130_fd_pr__pfet_01v8__bgidl_diff_26=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_26=0.30254
+  sky130_fd_pr__pfet_01v8__ub_diff_26=3.3049e-19
+  sky130_fd_pr__pfet_01v8__tvoff_diff_26=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_26=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_26=-0.011709
+  sky130_fd_pr__pfet_01v8__pdits_diff_26=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_26=-0.63249
+  sky130_fd_pr__pfet_01v8__eta0_diff_26=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_26=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_26=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_26=0.0015274
+  sky130_fd_pr__pfet_01v8__vsat_diff_26=-7322.9
+  sky130_fd_pr__pfet_01v8__vth0_diff_26=0.01124
+  sky130_fd_pr__pfet_01v8__cgidl_diff_26=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_26=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_26=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_26=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_26=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 027, W = 7.0, L = 1.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__pclm_diff_27=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_27=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_27=2.1179e-9
+  sky130_fd_pr__pfet_01v8__b1_diff_27=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_27=6.4042e-12
+  sky130_fd_pr__pfet_01v8__bgidl_diff_27=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_27=2.3627
+  sky130_fd_pr__pfet_01v8__tvoff_diff_27=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_27=0.12022
+  sky130_fd_pr__pfet_01v8__ub_diff_27=3.8976e-19
+  sky130_fd_pr__pfet_01v8__k2_diff_27=-0.0083062
+  sky130_fd_pr__pfet_01v8__pdits_diff_27=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_27=-0.34838
+  sky130_fd_pr__pfet_01v8__eta0_diff_27=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_27=-0.16849
+  sky130_fd_pr__pfet_01v8__pditsd_diff_27=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_27=0.0018165
+  sky130_fd_pr__pfet_01v8__vsat_diff_27=0.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_27=0.0033973
+  sky130_fd_pr__pfet_01v8__cgidl_diff_27=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_27=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_27=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_27=1.3861e-6
*
* sky130_fd_pr__pfet_01v8, Bin 028, W = 7.0, L = 2.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__kt1_diff_28=1.2233e-5
+  sky130_fd_pr__pfet_01v8__pclm_diff_28=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_28=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_28=2.6754e-10
+  sky130_fd_pr__pfet_01v8__b1_diff_28=0.0
+  sky130_fd_pr__pfet_01v8__bgidl_diff_28=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_28=2.9273
+  sky130_fd_pr__pfet_01v8__ua_diff_28=-3.7462e-12
+  sky130_fd_pr__pfet_01v8__tvoff_diff_28=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_28=0.093518
+  sky130_fd_pr__pfet_01v8__ub_diff_28=3.9115e-19
+  sky130_fd_pr__pfet_01v8__k2_diff_28=-0.010797
+  sky130_fd_pr__pfet_01v8__pdits_diff_28=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_28=-0.4
+  sky130_fd_pr__pfet_01v8__eta0_diff_28=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_28=-0.10184
+  sky130_fd_pr__pfet_01v8__pditsd_diff_28=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_28=0.0019362
+  sky130_fd_pr__pfet_01v8__vsat_diff_28=0.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_28=0.010296
+  sky130_fd_pr__pfet_01v8__cgidl_diff_28=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_28=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_28=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 029, W = 7.0, L = 4.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__rdsw_diff_29=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_29=-0.065705
+  sky130_fd_pr__pfet_01v8__pclm_diff_29=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_29=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_29=9.9946e-11
+  sky130_fd_pr__pfet_01v8__b1_diff_29=0.0
+  sky130_fd_pr__pfet_01v8__bgidl_diff_29=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_29=4.0
+  sky130_fd_pr__pfet_01v8__ua_diff_29=-1.9042e-12
+  sky130_fd_pr__pfet_01v8__tvoff_diff_29=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_29=0.058081
+  sky130_fd_pr__pfet_01v8__ub_diff_29=5.042e-19
+  sky130_fd_pr__pfet_01v8__k2_diff_29=-0.010381
+  sky130_fd_pr__pfet_01v8__pdits_diff_29=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_29=-0.4
+  sky130_fd_pr__pfet_01v8__eta0_diff_29=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_29=-0.066757
+  sky130_fd_pr__pfet_01v8__pditsd_diff_29=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_29=0.002706
+  sky130_fd_pr__pfet_01v8__vsat_diff_29=0.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_29=0.0027207
+  sky130_fd_pr__pfet_01v8__cgidl_diff_29=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_29=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 030, W = 7.0, L = 8.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__cgidl_diff_30=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_30=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_30=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_30=-0.4903
+  sky130_fd_pr__pfet_01v8__pclm_diff_30=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_30=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_30=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_30=6.6323e-10
+  sky130_fd_pr__pfet_01v8__ua_diff_30=-5.5272e-12
+  sky130_fd_pr__pfet_01v8__bgidl_diff_30=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_30=4.0
+  sky130_fd_pr__pfet_01v8__ub_diff_30=5.2353e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_30=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_30=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_30=0.057548
+  sky130_fd_pr__pfet_01v8__k2_diff_30=-0.010828
+  sky130_fd_pr__pfet_01v8__voff_diff_30=-0.4
+  sky130_fd_pr__pfet_01v8__a0_diff_30=-0.061742
+  sky130_fd_pr__pfet_01v8__pditsd_diff_30=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_30=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_30=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_30=0.002801
+  sky130_fd_pr__pfet_01v8__vth0_diff_30=0.0014165
*
* sky130_fd_pr__pfet_01v8, Bin 031, W = 7.0, L = 0.15
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__u0_diff_31=2.2779e-5
+  sky130_fd_pr__pfet_01v8__vth0_diff_31=-0.15393
+  sky130_fd_pr__pfet_01v8__cgidl_diff_31=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_31=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_31=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_31=0.37435
+  sky130_fd_pr__pfet_01v8__pclm_diff_31=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_31=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_31=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_31=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_31=-2.4799e-11
+  sky130_fd_pr__pfet_01v8__bgidl_diff_31=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_31=0.070567
+  sky130_fd_pr__pfet_01v8__ub_diff_31=1.2123e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_31=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_31=0.007
+  sky130_fd_pr__pfet_01v8__ags_diff_31=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_31=0.0033879
+  sky130_fd_pr__pfet_01v8__voff_diff_31=-0.090975
+  sky130_fd_pr__pfet_01v8__a0_diff_31=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_31=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_31=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_31=-16980.0
*
* sky130_fd_pr__pfet_01v8, Bin 032, W = 7.0, L = 0.18
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__pditsd_diff_32=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_32=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_32=-9382.4
+  sky130_fd_pr__pfet_01v8__u0_diff_32=0.00018292
+  sky130_fd_pr__pfet_01v8__vth0_diff_32=-0.089235
+  sky130_fd_pr__pfet_01v8__cgidl_diff_32=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_32=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_32=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_32=0.013313
+  sky130_fd_pr__pfet_01v8__pclm_diff_32=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_32=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_32=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_32=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_32=1.8792e-11
+  sky130_fd_pr__pfet_01v8__bgidl_diff_32=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_32=0.21464
+  sky130_fd_pr__pfet_01v8__ub_diff_32=1.0728e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_32=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_32=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_32=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_32=0.0012343
+  sky130_fd_pr__pfet_01v8__voff_diff_32=-0.076584
+  sky130_fd_pr__pfet_01v8__a0_diff_32=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 033, W = 7.0, L = 0.25
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__voff_diff_33=-0.13694
+  sky130_fd_pr__pfet_01v8__a0_diff_33=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_33=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_33=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_33=8184.4
+  sky130_fd_pr__pfet_01v8__u0_diff_33=0.00037451
+  sky130_fd_pr__pfet_01v8__vth0_diff_33=-0.043301
+  sky130_fd_pr__pfet_01v8__cgidl_diff_33=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_33=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_33=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_33=-0.053103
+  sky130_fd_pr__pfet_01v8__pclm_diff_33=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_33=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_33=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_33=2.1747e-9
+  sky130_fd_pr__pfet_01v8__ua_diff_33=3.1868e-12
+  sky130_fd_pr__pfet_01v8__bgidl_diff_33=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_33=0.32299
+  sky130_fd_pr__pfet_01v8__ub_diff_33=1.7315e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_33=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_33=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_33=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_33=-0.0032062
*
* sky130_fd_pr__pfet_01v8, Bin 034, W = 7.0, L = 0.5
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__pdits_diff_34=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_34=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_34=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_34=-0.014635
+  sky130_fd_pr__pfet_01v8__voff_diff_34=-0.94104
+  sky130_fd_pr__pfet_01v8__a0_diff_34=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_34=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_34=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_34=18609.0
+  sky130_fd_pr__pfet_01v8__u0_diff_34=0.0015571
+  sky130_fd_pr__pfet_01v8__vth0_diff_34=-0.0010985
+  sky130_fd_pr__pfet_01v8__cgidl_diff_34=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_34=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_34=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_34=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_34=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_34=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_34=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_34=1.4168e-10
+  sky130_fd_pr__pfet_01v8__ua_diff_34=3.2727e-12
+  sky130_fd_pr__pfet_01v8__bgidl_diff_34=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_34=0.48298
+  sky130_fd_pr__pfet_01v8__ub_diff_34=3.9575e-19
*
* sky130_fd_pr__pfet_01v8, Bin 035, W = 0.42, L = 1.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__bgidl_diff_35=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_35=2.7859
+  sky130_fd_pr__pfet_01v8__ub_diff_35=6.0253e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_35=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_35=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_35=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_35=-0.0086286
+  sky130_fd_pr__pfet_01v8__voff_diff_35=-0.39652
+  sky130_fd_pr__pfet_01v8__a0_diff_35=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_35=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_35=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_35=0.0027005
+  sky130_fd_pr__pfet_01v8__vsat_diff_35=0.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_35=0.012947
+  sky130_fd_pr__pfet_01v8__cgidl_diff_35=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_35=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_35=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_35=-5.8416e-6
+  sky130_fd_pr__pfet_01v8__pclm_diff_35=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_35=1.0933e-8
+  sky130_fd_pr__pfet_01v8__b1_diff_35=2.1687e-11
+  sky130_fd_pr__pfet_01v8__agidl_diff_35=-8.4706e-10
+  sky130_fd_pr__pfet_01v8__ua_diff_35=1.3766e-12
*
* sky130_fd_pr__pfet_01v8, Bin 036, W = 0.42, L = 20.0
* -----------------------------------
+  sky130_fd_pr__pfet_01v8__agidl_diff_36=1.9928e-8
+  sky130_fd_pr__pfet_01v8__b1_diff_36=3.5968e-11
+  sky130_fd_pr__pfet_01v8__ua_diff_36=-3.2012e-11
+  sky130_fd_pr__pfet_01v8__bgidl_diff_36=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_36=4.0
+  sky130_fd_pr__pfet_01v8__ub_diff_36=2.0645e-20
+  sky130_fd_pr__pfet_01v8__pdits_diff_36=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_36=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_36=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_36=-0.0021702
+  sky130_fd_pr__pfet_01v8__voff_diff_36=-0.4
+  sky130_fd_pr__pfet_01v8__eta0_diff_36=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_36=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_36=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_36=-0.00031963
+  sky130_fd_pr__pfet_01v8__vsat_diff_36=20006.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_36=0.043888
+  sky130_fd_pr__pfet_01v8__cgidl_diff_36=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_36=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_36=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_36=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_36=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_36=-7.6937e-9
*
* sky130_fd_pr__pfet_01v8, Bin 037, W = 0.42, L = 2.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__b0_diff_37=-2.3635e-8
+  sky130_fd_pr__pfet_01v8__agidl_diff_37=-1.9945e-10
+  sky130_fd_pr__pfet_01v8__b1_diff_37=-3.9942e-10
+  sky130_fd_pr__pfet_01v8__ua_diff_37=-7.2077e-12
+  sky130_fd_pr__pfet_01v8__bgidl_diff_37=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_37=3.7892
+  sky130_fd_pr__pfet_01v8__ub_diff_37=7.308e-19
+  sky130_fd_pr__pfet_01v8__tvoff_diff_37=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_37=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_37=-0.0068908
+  sky130_fd_pr__pfet_01v8__pdits_diff_37=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_37=-0.39966
+  sky130_fd_pr__pfet_01v8__eta0_diff_37=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_37=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_37=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_37=0.0032114
+  sky130_fd_pr__pfet_01v8__vsat_diff_37=0.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_37=0.032454
+  sky130_fd_pr__pfet_01v8__cgidl_diff_37=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_37=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_37=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_37=1.6838e-5
+  sky130_fd_pr__pfet_01v8__pclm_diff_37=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 038, W = 0.42, L = 4.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__pclm_diff_38=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_38=-5.0764e-8
+  sky130_fd_pr__pfet_01v8__agidl_diff_38=1.6018e-10
+  sky130_fd_pr__pfet_01v8__b1_diff_38=1.5533e-10
+  sky130_fd_pr__pfet_01v8__ua_diff_38=-3.8513e-13
+  sky130_fd_pr__pfet_01v8__bgidl_diff_38=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_38=4.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_38=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_38=0.0
+  sky130_fd_pr__pfet_01v8__ub_diff_38=6.0269e-19
+  sky130_fd_pr__pfet_01v8__k2_diff_38=-0.012379
+  sky130_fd_pr__pfet_01v8__pdits_diff_38=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_38=-0.4
+  sky130_fd_pr__pfet_01v8__eta0_diff_38=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_38=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_38=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_38=0.0029622
+  sky130_fd_pr__pfet_01v8__vsat_diff_38=0.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_38=0.00040399
+  sky130_fd_pr__pfet_01v8__cgidl_diff_38=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_38=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_38=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_38=-0.37766
*
* sky130_fd_pr__pfet_01v8, Bin 039, W = 0.42, L = 8.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__kt1_diff_39=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_39=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_39=3.2804e-8
+  sky130_fd_pr__pfet_01v8__agidl_diff_39=1.0718e-8
+  sky130_fd_pr__pfet_01v8__b1_diff_39=9.5861e-11
+  sky130_fd_pr__pfet_01v8__bgidl_diff_39=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_39=4.0
+  sky130_fd_pr__pfet_01v8__ua_diff_39=-6.752e-11
+  sky130_fd_pr__pfet_01v8__tvoff_diff_39=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_39=0.0
+  sky130_fd_pr__pfet_01v8__ub_diff_39=7.8184e-19
+  sky130_fd_pr__pfet_01v8__k2_diff_39=-0.01397
+  sky130_fd_pr__pfet_01v8__pdits_diff_39=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_39=-0.4
+  sky130_fd_pr__pfet_01v8__eta0_diff_39=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_39=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_39=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_39=0.0035533
+  sky130_fd_pr__pfet_01v8__vsat_diff_39=20051.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_39=0.0027392
+  sky130_fd_pr__pfet_01v8__cgidl_diff_39=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_39=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_39=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 040, W = 0.42, L = 0.15
* -----------------------------------
+  sky130_fd_pr__pfet_01v8__rdsw_diff_40=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_40=-0.43866
+  sky130_fd_pr__pfet_01v8__pclm_diff_40=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_40=3.2204e-7
+  sky130_fd_pr__pfet_01v8__b1_diff_40=2.0586e-8
+  sky130_fd_pr__pfet_01v8__agidl_diff_40=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_40=-7.7662e-11
+  sky130_fd_pr__pfet_01v8__bgidl_diff_40=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_40=7.0
+  sky130_fd_pr__pfet_01v8__ub_diff_40=6.1327e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_40=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_40=0.0052792
+  sky130_fd_pr__pfet_01v8__ags_diff_40=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_40=-0.0067948
+  sky130_fd_pr__pfet_01v8__voff_diff_40=-0.21256
+  sky130_fd_pr__pfet_01v8__a0_diff_40=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_40=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_40=0.13689
+  sky130_fd_pr__pfet_01v8__vsat_diff_40=-50000.0
+  sky130_fd_pr__pfet_01v8__u0_diff_40=0.00074341
+  sky130_fd_pr__pfet_01v8__vth0_diff_40=-0.013683
+  sky130_fd_pr__pfet_01v8__cgidl_diff_40=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_40=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 041, W = 0.42, L = 0.18
* -----------------------------------
+  sky130_fd_pr__pfet_01v8__cgidl_diff_41=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_41=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_41=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_41=-0.39913
+  sky130_fd_pr__pfet_01v8__pclm_diff_41=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_41=2.4612e-7
+  sky130_fd_pr__pfet_01v8__b1_diff_41=3.3783e-9
+  sky130_fd_pr__pfet_01v8__agidl_diff_41=-4.3155e-9
+  sky130_fd_pr__pfet_01v8__ua_diff_41=-4.9909e-10
+  sky130_fd_pr__pfet_01v8__bgidl_diff_41=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_41=-0.2
+  sky130_fd_pr__pfet_01v8__ub_diff_41=9.3187e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_41=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_41=6.198e-7
+  sky130_fd_pr__pfet_01v8__ags_diff_41=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_41=0.011456
+  sky130_fd_pr__pfet_01v8__voff_diff_41=-0.5
+  sky130_fd_pr__pfet_01v8__a0_diff_41=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_41=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_41=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_41=5887.7
+  sky130_fd_pr__pfet_01v8__u0_diff_41=-0.00039577
+  sky130_fd_pr__pfet_01v8__vth0_diff_41=0.10661
*
* sky130_fd_pr__pfet_01v8, Bin 042, W = 0.42, L = 0.5
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__u0_diff_42=0.0018823
+  sky130_fd_pr__pfet_01v8__vth0_diff_42=0.037859
+  sky130_fd_pr__pfet_01v8__cgidl_diff_42=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_42=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_42=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_42=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_42=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_42=3.6809e-8
+  sky130_fd_pr__pfet_01v8__b1_diff_42=-2.2779e-9
+  sky130_fd_pr__pfet_01v8__agidl_diff_42=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_42=-1.0153e-11
+  sky130_fd_pr__pfet_01v8__bgidl_diff_42=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_42=0.3823
+  sky130_fd_pr__pfet_01v8__ub_diff_42=5.6326e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_42=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_42=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_42=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_42=-0.0070988
+  sky130_fd_pr__pfet_01v8__voff_diff_42=-1.0162
+  sky130_fd_pr__pfet_01v8__a0_diff_42=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_42=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_42=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_42=19837.0
*
* sky130_fd_pr__pfet_01v8, Bin 043, W = 0.55, L = 1.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__pditsd_diff_43=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_43=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_43=119930.0
+  sky130_fd_pr__pfet_01v8__u0_diff_43=7.5664e-5
+  sky130_fd_pr__pfet_01v8__vth0_diff_43=0.0014854
+  sky130_fd_pr__pfet_01v8__cgidl_diff_43=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_43=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_43=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_43=-2.7282e-6
+  sky130_fd_pr__pfet_01v8__pclm_diff_43=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_43=7.5463e-8
+  sky130_fd_pr__pfet_01v8__b1_diff_43=3.7039e-12
+  sky130_fd_pr__pfet_01v8__agidl_diff_43=-1.3767e-10
+  sky130_fd_pr__pfet_01v8__ua_diff_43=-4.9877e-10
+  sky130_fd_pr__pfet_01v8__bgidl_diff_43=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_43=2.7489
+  sky130_fd_pr__pfet_01v8__ub_diff_43=7.6183e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_43=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_43=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_43=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_43=-0.0061079
+  sky130_fd_pr__pfet_01v8__voff_diff_43=-0.39681
+  sky130_fd_pr__pfet_01v8__a0_diff_43=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 044, W = 0.55, L = 2.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__voff_diff_44=-0.39995
+  sky130_fd_pr__pfet_01v8__a0_diff_44=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_44=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_44=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_44=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_44=0.0030766
+  sky130_fd_pr__pfet_01v8__vth0_diff_44=0.027061
+  sky130_fd_pr__pfet_01v8__cgidl_diff_44=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_44=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_44=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_44=-8.5609e-7
+  sky130_fd_pr__pfet_01v8__pclm_diff_44=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_44=-1.9527e-8
+  sky130_fd_pr__pfet_01v8__b1_diff_44=-1.746e-9
+  sky130_fd_pr__pfet_01v8__agidl_diff_44=1.1392e-10
+  sky130_fd_pr__pfet_01v8__ua_diff_44=9.5215e-12
+  sky130_fd_pr__pfet_01v8__bgidl_diff_44=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_44=3.9606
+  sky130_fd_pr__pfet_01v8__ub_diff_44=6.6875e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_44=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_44=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_44=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_44=-0.0090663
*
* sky130_fd_pr__pfet_01v8, Bin 045, W = 0.55, L = 4.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__pdits_diff_45=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_45=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_45=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_45=-0.0099384
+  sky130_fd_pr__pfet_01v8__voff_diff_45=-0.4
+  sky130_fd_pr__pfet_01v8__a0_diff_45=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_45=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_45=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_45=20111.0
+  sky130_fd_pr__pfet_01v8__u0_diff_45=0.0028513
+  sky130_fd_pr__pfet_01v8__vth0_diff_45=-0.0079656
+  sky130_fd_pr__pfet_01v8__cgidl_diff_45=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_45=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_45=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_45=-0.31682
+  sky130_fd_pr__pfet_01v8__pclm_diff_45=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_45=-2.7446e-8
+  sky130_fd_pr__pfet_01v8__b1_diff_45=7.2475e-8
+  sky130_fd_pr__pfet_01v8__agidl_diff_45=6.5747e-9
+  sky130_fd_pr__pfet_01v8__ua_diff_45=-5.5618e-11
+  sky130_fd_pr__pfet_01v8__bgidl_diff_45=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_45=4.0
+  sky130_fd_pr__pfet_01v8__ub_diff_45=7.0725e-19
*
* sky130_fd_pr__pfet_01v8, Bin 046, W = 0.55, L = 8.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__bgidl_diff_46=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_46=4.0
+  sky130_fd_pr__pfet_01v8__ub_diff_46=6.9222e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_46=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_46=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_46=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_46=-0.013366
+  sky130_fd_pr__pfet_01v8__voff_diff_46=-0.4
+  sky130_fd_pr__pfet_01v8__a0_diff_46=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_46=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_46=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_46=0.00349
+  sky130_fd_pr__pfet_01v8__vsat_diff_46=0.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_46=0.0039395
+  sky130_fd_pr__pfet_01v8__cgidl_diff_46=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_46=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_46=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_46=-0.58418
+  sky130_fd_pr__pfet_01v8__pclm_diff_46=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_46=-2.1294e-8
+  sky130_fd_pr__pfet_01v8__b1_diff_46=-1.2248e-10
+  sky130_fd_pr__pfet_01v8__agidl_diff_46=-1.7596e-10
+  sky130_fd_pr__pfet_01v8__ua_diff_46=-2.4775e-12
*
* sky130_fd_pr__pfet_01v8, Bin 047, W = 0.55, L = 0.15
* -----------------------------------
+  sky130_fd_pr__pfet_01v8__agidl_diff_47=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_47=2.3324e-8
+  sky130_fd_pr__pfet_01v8__ua_diff_47=-4.2037e-11
+  sky130_fd_pr__pfet_01v8__bgidl_diff_47=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_47=1.0273
+  sky130_fd_pr__pfet_01v8__ub_diff_47=5.792e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_47=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_47=-6.8313e-7
+  sky130_fd_pr__pfet_01v8__ags_diff_47=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_47=0.0089906
+  sky130_fd_pr__pfet_01v8__voff_diff_47=-0.34706
+  sky130_fd_pr__pfet_01v8__eta0_diff_47=0.18556
+  sky130_fd_pr__pfet_01v8__a0_diff_47=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_47=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_47=0.00075996
+  sky130_fd_pr__pfet_01v8__vsat_diff_47=-34891.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_47=-0.015495
+  sky130_fd_pr__pfet_01v8__cgidl_diff_47=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_47=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_47=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_47=0.1866
+  sky130_fd_pr__pfet_01v8__pclm_diff_47=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_47=6.8027e-7
*
* sky130_fd_pr__pfet_01v8, Bin 048, W = 0.55, L = 0.5
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__b0_diff_48=2.4391e-8
+  sky130_fd_pr__pfet_01v8__agidl_diff_48=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_48=1.6514e-8
+  sky130_fd_pr__pfet_01v8__ua_diff_48=-4.9634e-12
+  sky130_fd_pr__pfet_01v8__bgidl_diff_48=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_48=0.37279
+  sky130_fd_pr__pfet_01v8__ub_diff_48=4.8904e-19
+  sky130_fd_pr__pfet_01v8__tvoff_diff_48=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_48=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_48=-0.016336
+  sky130_fd_pr__pfet_01v8__pdits_diff_48=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_48=-0.94461
+  sky130_fd_pr__pfet_01v8__eta0_diff_48=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_48=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_48=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_48=0.0015741
+  sky130_fd_pr__pfet_01v8__vsat_diff_48=19810.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_48=0.038899
+  sky130_fd_pr__pfet_01v8__cgidl_diff_48=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_48=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_48=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_48=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_48=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 049, W = 0.64, L = 0.15
* -----------------------------------
+  sky130_fd_pr__pfet_01v8__pclm_diff_49=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_49=8.6951e-7
+  sky130_fd_pr__pfet_01v8__agidl_diff_49=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_49=9.8831e-9
+  sky130_fd_pr__pfet_01v8__ua_diff_49=-2.0555e-10
+  sky130_fd_pr__pfet_01v8__bgidl_diff_49=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_49=4.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_49=-4.1951e-7
+  sky130_fd_pr__pfet_01v8__ags_diff_49=0.0
+  sky130_fd_pr__pfet_01v8__ub_diff_49=6.2299e-19
+  sky130_fd_pr__pfet_01v8__k2_diff_49=0.014274
+  sky130_fd_pr__pfet_01v8__pdits_diff_49=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_49=-0.4
+  sky130_fd_pr__pfet_01v8__eta0_diff_49=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_49=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_49=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_49=0.000184
+  sky130_fd_pr__pfet_01v8__vsat_diff_49=23896.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_49=-0.10123
+  sky130_fd_pr__pfet_01v8__cgidl_diff_49=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_49=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_49=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_49=0.21394
*
* sky130_fd_pr__pfet_01v8, Bin 050, W = 0.84, L = 0.15
* -----------------------------------
+  sky130_fd_pr__pfet_01v8__kt1_diff_50=0.14725
+  sky130_fd_pr__pfet_01v8__pclm_diff_50=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_50=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_50=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_50=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_50=-2.4122e-10
+  sky130_fd_pr__pfet_01v8__bgidl_diff_50=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_50=-0.22096
+  sky130_fd_pr__pfet_01v8__ub_diff_50=6.4451e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_50=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_50=-2.192e-5
+  sky130_fd_pr__pfet_01v8__ags_diff_50=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_50=-0.024696
+  sky130_fd_pr__pfet_01v8__voff_diff_50=0.0072572
+  sky130_fd_pr__pfet_01v8__a0_diff_50=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_50=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_50=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_50=-20000.0
+  sky130_fd_pr__pfet_01v8__u0_diff_50=0.00025044
+  sky130_fd_pr__pfet_01v8__vth0_diff_50=-0.11705
+  sky130_fd_pr__pfet_01v8__cgidl_diff_50=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_50=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_50=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 051, W = 1.65, L = 0.15
* -----------------------------------
+  sky130_fd_pr__pfet_01v8__rdsw_diff_51=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_51=0.2841
+  sky130_fd_pr__pfet_01v8__pclm_diff_51=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_51=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_51=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_51=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_51=-2.8822e-11
+  sky130_fd_pr__pfet_01v8__bgidl_diff_51=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_51=1.3308
+  sky130_fd_pr__pfet_01v8__ub_diff_51=3.1525e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_51=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_51=0.00036195
+  sky130_fd_pr__pfet_01v8__ags_diff_51=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_51=-0.0044952
+  sky130_fd_pr__pfet_01v8__voff_diff_51=-0.16115
+  sky130_fd_pr__pfet_01v8__a0_diff_51=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_51=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_51=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_51=-16955.0
+  sky130_fd_pr__pfet_01v8__u0_diff_51=0.00035368
+  sky130_fd_pr__pfet_01v8__vth0_diff_51=-0.10495
+  sky130_fd_pr__pfet_01v8__cgidl_diff_51=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_51=0.0
.include "sky130_fd_pr__pfet_01v8.pm3.spice"
