* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param sky130_fd_pr__special_nfet_pass_flash__tox_slope_spectre=0.0
.param sky130_fd_pr__special_nfet_pass_flash__vth0_slope_spectre=0.0
* statistics {
*   process {
*   }
*   mismatch {
*     vary sky130_fd_pr__special_nfet_pass_flash__tox_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__special_nfet_pass_flash__vth0_slope_spectre dist=gauss std = 1.0
*   }
* }
.subckt sky130_fd_pr__special_nfet_pass_flash d g s b
.param l=1 w=1 ad=0 as=0 pd=0 ps=0 nrd=0 nrs=0 mult=1.0
Msky130_fd_pr__special_nfet_pass_flash d g s b sky130_fd_pr__special_nfet_pass_flash__model l={l} w={w} ad={ad} as={as} pd={pd} ps={ps} nrd={nrd} nrs={nrs}
.model sky130_fd_pr__special_nfet_pass_flash__model.0 nmos
+  lmin=1.495e-007 lmax=1.505e-007 wmin=4.495e-007 wmax=4.505e-7
+  level=49.0
+  tnom=30.0
+  version=3.2
+  tox={1.1628e-008*sky130_fd_pr__special_nfet_pass_flash__tox_mult+sky130_fd_pr__special_nfet_pass_flash__tox_slope_spectre*(1.1628e-008*sky130_fd_pr__special_nfet_pass_flash__tox_mult*(sky130_fd_pr__special_nfet_pass_flash__tox_slope/sqrt(l*w*mult)))}
+  toxm=1.1628e-8
+  xj=1.2e-7
+  nch=1.1247e+18
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint={0+sky130_fd_pr__special_nfet_pass_flash__lint_diff}
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint={0+sky130_fd_pr__special_nfet_pass_flash__wint_diff}
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  mobmod=1.0
+  binunit=2.0
+  dwg={0+sky130_fd_pr__special_nfet_pass_flash__dwg_diff}
+  dwb=0.0
* Diode Parameters
+  ldif=0.0
+  hdif=0.0
+  rd=0.0
+  rs=0.0
+  rsc=0.0
+  rdc=0.0
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={1.1466+sky130_fd_pr__special_nfet_pass_flash__vth0_diff_0+sky130_fd_pr__special_nfet_pass_flash__vth0_slope_spectre*(sky130_fd_pr__special_nfet_pass_flash__vth0_slope/sqrt(w*l*mult))}
+  k1=0.60764
+  k2={-0.12236+sky130_fd_pr__special_nfet_pass_flash__k2_diff_0}
+  k3={0+sky130_fd_pr__special_nfet_pass_flash__k3_diff}
+  dvt0={0+sky130_fd_pr__special_nfet_pass_flash__dvt0_diff}
+  dvt1=0.53
+  dvt2=0.0
+  dvt0w={0+sky130_fd_pr__special_nfet_pass_flash__dvt0w_diff}
+  dvt1w=400000.0
+  dvt2w=0.0
+  nlx={0+sky130_fd_pr__special_nfet_pass_flash__nlx_diff}
+  w0=1.0e-9
+  k3b=0.0
+  ngate=1.0e+30
+  vfb=-0.9693
* Mobility Parameters
+  vsat={93196+sky130_fd_pr__special_nfet_pass_flash__vsat_diff_0}
+  ua=1.0846e-9
+  ub=1.2522e-18
+  uc=7.8332e-11
+  rdsw=251.69
+  prwb=0.0
+  prwg=0.0
+  wr=1.0
+  u0={0.038044+sky130_fd_pr__special_nfet_pass_flash__u0_diff_0}
+  a0=0.4436
+  keta=0.073859
+  a1=0.0
+  a2=0.99
+  ags=0.0
+  b0=0.0
+  b1=0.0
* Subthreshold Current Parameters
+  voff={-0.25275+sky130_fd_pr__special_nfet_pass_flash__voff_diff_0}
+  nfactor={0.94875+sky130_fd_pr__special_nfet_pass_flash__nfactor_diff_0}
+  cit={0+sky130_fd_pr__special_nfet_pass_flash__cit_diff}
+  cdsc={0+sky130_fd_pr__special_nfet_pass_flash__cdsc_diff}
+  cdscb={0+sky130_fd_pr__special_nfet_pass_flash__cdscb_diff}
+  cdscd={0+sky130_fd_pr__special_nfet_pass_flash__cdscd_diff}
+  eta0=0.09373
+  etab=-0.01485
+  dsub=0.176
* Rout Parameters
+  pclm=0.080615
+  pdiblc1=0.025
+  pdiblc2=0.085152
+  pdiblcb=0.055737
+  drout=0.16
+  pscbe1=7.8166e+8
+  pscbe2=1.0e-20
+  pvag=0.0
+  delta=0.02553
+  alpha0=0.00019736
+  alpha1=0.0
+  beta0=24.801
* Temperature Effects Parameters
+  kt1={-0.31006+sky130_fd_pr__special_nfet_pass_flash__kt1_diff_0}
+  kt2={-0.041175+sky130_fd_pr__special_nfet_pass_flash__kt2_diff}
+  at=13357.0
+  ute=-0.81863
+  ua1=2.3327e-9
+  ub1=-1.6577e-18
+  uc1=6.275e-11
+  kt1l={0+sky130_fd_pr__special_nfet_pass_flash__kt1l_diff}
+  prt=0.0
* Capacitance Parameters
+  cj={0.0012651*sky130_fd_pr__special_nfet_pass_flash__ajunction_mult}
+  mj=0.3608
+  pb=0.729
+  cjsw={7.3442e-011*sky130_fd_pr__special_nfet_pass_flash__pjunction_mult}
+  mjsw=0.13
+  pbsw=0.729
+  cjswg={7.3442e-011*sky130_fd_pr__special_nfet_pass_flash__pjunction_mult}
+  mjswg=0.13
+  pbswg=0.729
+  tpb=0.0012287
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.0
+  tcjsw=0.0
+  tcjswg=0.0
+  js=0.000375
+  jsw=6.0e-10
+  nj=1.3574
+  xti=0.13
+  cgdo={3.0674e-010*sky130_fd_pr__special_nfet_pass_flash__overlap_mult}
+  cgso={3.0674e-010*sky130_fd_pr__special_nfet_pass_flash__overlap_mult}
+  cgbo=0.0
+  capmod=3.0
+  nqsmod=0.0
+  elm=0.0
+  xpart=0.0
+  cgsl={5e-011*sky130_fd_pr__special_nfet_pass_flash__overlap_mult}
+  cgdl={5e-011*sky130_fd_pr__special_nfet_pass_flash__overlap_mult}
+  ckappa=0.6
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc={1.8739e-008+sky130_fd_pr__special_nfet_pass_flash__dlc_diff+sky130_fd_pr__special_nfet_pass_flash__dlc_rotweak}
+  dwc={0+sky130_fd_pr__special_nfet_pass_flash__dwc_diff}
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
+  noimod=2.0
+  noia={2.1700000e+41*1.6e-21}
+  noib={3.2000000e+24*1.6e-21}
+  noic={-1.7200000e+06*1.6e-21}
+  em=4.1000000e+7
+  ef=0.89
.model sky130_fd_pr__special_nfet_pass_flash__model.1 nmos
+  lmin=1.49e-007 lmax=1.51e-007 wmin=3.45e-007 wmax=3.55e-7
+  level=49.0
+  tnom=30.0
+  version=3.2
+  tox={1.1628e-008*sky130_fd_pr__special_nfet_pass_flash__tox_mult+sky130_fd_pr__special_nfet_pass_flash__tox_slope_spectre*(1.1628e-008*sky130_fd_pr__special_nfet_pass_flash__tox_mult*(sky130_fd_pr__special_nfet_pass_flash__tox_slope/sqrt(l*w*mult)))}
+  toxm=1.1628e-8
+  xj=1.2e-7
+  nch=1.1247e+18
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint={0+sky130_fd_pr__special_nfet_pass_flash__lint_diff}
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint={0+sky130_fd_pr__special_nfet_pass_flash__wint_diff}
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  mobmod=1.0
+  binunit=2.0
+  dwg={0+sky130_fd_pr__special_nfet_pass_flash__dwg_diff}
+  dwb=0.0
* Diode Parameters
+  ldif=0.0
+  hdif=0.0
+  rd=0.0
+  rs=0.0
+  rsc=0.0
+  rdc=0.0
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.97306+sky130_fd_pr__special_nfet_pass_flash__vth0_diff_1+sky130_fd_pr__special_nfet_pass_flash__vth0_slope_spectre*(sky130_fd_pr__special_nfet_pass_flash__vth0_slope/sqrt(w*l*mult))}
+  k1=0.60764
+  k2={-0.14289+sky130_fd_pr__special_nfet_pass_flash__k2_diff_1}
+  k3={0+sky130_fd_pr__special_nfet_pass_flash__k3_diff}
+  dvt0={0+sky130_fd_pr__special_nfet_pass_flash__dvt0_diff}
+  dvt1=0.53
+  dvt2=0.0
+  dvt0w={0+sky130_fd_pr__special_nfet_pass_flash__dvt0w_diff}
+  dvt1w=400000.0
+  dvt2w=0.0
+  nlx={0+sky130_fd_pr__special_nfet_pass_flash__nlx_diff}
+  w0=1.0e-9
+  k3b=0.0
+  ngate=1.0e+23
+  vfb=-0.9693
* Mobility Parameters
+  vsat={82954+sky130_fd_pr__special_nfet_pass_flash__vsat_diff_1}
+  ua=1.7786e-9
+  ub=-2.0e-19
+  uc=7.8332e-11
+  rdsw=251.69
+  prwb=0.0
+  prwg=0.0
+  wr=1.0
+  u0={0.038274+sky130_fd_pr__special_nfet_pass_flash__u0_diff_1}
+  a0=1.0
+  keta=0.073859
+  a1=0.0
+  a2=0.99
+  ags=0.1
+  b0=0.0
+  b1=0.0
* Subthreshold Current Parameters
+  voff={-0.1198+sky130_fd_pr__special_nfet_pass_flash__voff_diff_1}
+  nfactor={0.85834+sky130_fd_pr__special_nfet_pass_flash__nfactor_diff_1}
+  cit={0+sky130_fd_pr__special_nfet_pass_flash__cit_diff}
+  cdsc={0+sky130_fd_pr__special_nfet_pass_flash__cdsc_diff}
+  cdscb={0+sky130_fd_pr__special_nfet_pass_flash__cdscb_diff}
+  cdscd={0+sky130_fd_pr__special_nfet_pass_flash__cdscd_diff}
+  eta0=0.09373
+  etab=-0.01485
+  dsub=0.176
* Rout Parameters
+  pclm=0.080615
+  pdiblc1=0.025
+  pdiblc2=0.085152
+  pdiblcb=0.055737
+  drout=0.16
+  pscbe1=7.8166e+8
+  pscbe2=1.0e-20
+  pvag=0.0
+  delta=0.02553
+  alpha0=0.00019736
+  alpha1=0.0
+  beta0=24.801
* Temperature Effects Parameters
+  kt1={-0.30763+sky130_fd_pr__special_nfet_pass_flash__kt1_diff_1}
+  kt2={-0.041175+sky130_fd_pr__special_nfet_pass_flash__kt2_diff}
+  at=33000.0
+  ute=-0.6
+  ua1=2.3327e-9
+  ub1=-1.6577e-18
+  uc1=6.275e-11
+  kt1l={0+sky130_fd_pr__special_nfet_pass_flash__kt1l_diff}
+  prt=0.0
* Capacitance Parameters
+  cj={0.00106*sky130_fd_pr__special_nfet_pass_flash__ajunction_mult}
+  mj=0.4
+  pb=0.729
+  cjsw={2.3162e-011*sky130_fd_pr__special_nfet_pass_flash__pjunction_mult}
+  mjsw=0.4
+  pbsw=0.729
+  cjswg={2.3162e-011*sky130_fd_pr__special_nfet_pass_flash__pjunction_mult}
+  mjswg=0.4
+  pbswg=0.729
+  tpb=0.0012287
+  tpbsw=0.0
+  tpbswg=0.0
+  tcj=0.0007
+  tcjsw=0.0015
+  tcjswg=0.0015
+  js=0.000375
+  jsw=6.0e-10
+  nj=1.3574
+  xti=0.13
+  cgdo={1.97e-010*sky130_fd_pr__special_nfet_pass_flash__overlap_mult}
+  cgso={1.97e-010*sky130_fd_pr__special_nfet_pass_flash__overlap_mult}
+  cgbo=0.0
+  capmod=3.0
+  nqsmod=0.0
+  elm=0.0
+  xpart=0.0
+  cgsl={0*sky130_fd_pr__special_nfet_pass_flash__overlap_mult}
+  cgdl={0*sky130_fd_pr__special_nfet_pass_flash__overlap_mult}
+  ckappa=0.6
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc={2.3232e-008+sky130_fd_pr__special_nfet_pass_flash__dlc_diff+sky130_fd_pr__special_nfet_pass_flash__dlc_rotweak}
+  dwc={0+sky130_fd_pr__special_nfet_pass_flash__dwc_diff}
+  vfbcv=-1.0
+  acde=0.4
+  moin=15.0
+  noff=4.0
+  voffcv=-0.24172
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
+  noimod=2.0
+  noia=3.472e+20
+  noib=5120.0
+  noic=-2.752e-15
+  em=4.1000000e+7
+  ef=0.89
.ends sky130_fd_pr__special_nfet_pass_flash
