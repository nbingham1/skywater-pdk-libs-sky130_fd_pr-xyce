* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 63
.param
+  sky130_fd_pr__nfet_01v8__toxe_mult=1.0
+  sky130_fd_pr__nfet_01v8__rshn_mult=1.0
+  sky130_fd_pr__nfet_01v8__overlap_mult=1.0
+  sky130_fd_pr__nfet_01v8__lint_diff=0.0
+  sky130_fd_pr__nfet_01v8__wint_diff=0.0
+  sky130_fd_pr__nfet_01v8__dlc_diff=0.0
+  sky130_fd_pr__nfet_01v8__dwc_diff=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 000, W = 1.26, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__voff_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_0=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 001, W = 1.68, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__eta0_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_1=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 002, W = 1.0, L = 1.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__nfactor_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_2=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 003, W = 1.0, L = 2.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__keta_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_3=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 004, W = 1.0, L = 4.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__pdits_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_4=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 005, W = 1.0, L = 8.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__pdits_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_5=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 006, W = 1.0, L = 0.15
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__pclm_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_6=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 007, W = 1.0, L = 0.18
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__b0_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_7=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 008, W = 1.0, L = 0.25
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__a0_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_8=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 009, W = 1.0, L = 0.5
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__kt1_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_9=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 010, W = 2.0, L = 0.15
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__ags_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_10=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 011, W = 3.0, L = 1.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__pclm_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_11=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 012, W = 3.0, L = 2.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__pditsd_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_12=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 013, W = 3.0, L = 4.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__pdits_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_13=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 014, W = 3.0, L = 8.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__b0_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_14=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 015, W = 3.0, L = 0.15
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__kt1_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_15=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 016, W = 3.0, L = 0.18
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__a0_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_16=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 017, W = 3.0, L = 0.25
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__a0_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_17=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 018, W = 3.0, L = 0.5
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__ub_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_18=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 019, W = 5.0, L = 1.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__eta0_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_19=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 020, W = 5.0, L = 2.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__ua_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_20=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 021, W = 5.0, L = 4.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__ags_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_21=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 022, W = 5.0, L = 8.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__pclm_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_22=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 023, W = 5.0, L = 0.15
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__pditsd_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_23=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 024, W = 5.0, L = 0.18
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__pdits_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_24=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 025, W = 5.0, L = 0.25
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__b0_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_25=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 026, W = 5.0, L = 0.5
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__kt1_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_26=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 027, W = 7.0, L = 1.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__a0_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_27=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 028, W = 7.0, L = 2.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__a0_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_28=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 029, W = 7.0, L = 4.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__ub_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_29=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 030, W = 7.0, L = 8.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__eta0_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_30=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 031, W = 7.0, L = 0.15
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__ua_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_31=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 032, W = 7.0, L = 0.18
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__ags_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_32=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 033, W = 7.0, L = 0.25
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__pclm_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_33=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 034, W = 7.0, L = 0.5
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__pditsd_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_34=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 035, W = 0.42, L = 1.0
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__pdits_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_35=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 036, W = 0.42, L = 20.0
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__b0_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_36=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 037, W = 0.42, L = 2.0
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__kt1_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_37=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 038, W = 0.42, L = 4.0
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__a0_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_38=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 039, W = 0.42, L = 8.0
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__a0_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_39=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 040, W = 0.42, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__a0_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_40=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 041, W = 0.42, L = 0.18
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__eta0_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_41=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 042, W = 0.42, L = 0.5
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__ua_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_42=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 043, W = 0.55, L = 1.0
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__ags_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_43=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 044, W = 0.55, L = 2.0
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__pclm_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_44=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 045, W = 0.55, L = 4.0
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__pditsd_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_45=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 046, W = 0.55, L = 8.0
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__pdits_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_46=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 047, W = 0.55, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__b0_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_47=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 048, W = 0.55, L = 0.5
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__kt1_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_48=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 049, W = 0.64, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__a0_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_49=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 050, W = 0.84, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__a0_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_50=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 051, W = 0.74, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__nfactor_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_51=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 052, W = 0.36, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__nfactor_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_52=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 053, W = 0.39, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__nfactor_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_53=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 054, W = 0.52, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__nfactor_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_54=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 055, W = 0.54, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__nfactor_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_55=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 056, W = 0.58, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__nfactor_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_56=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 057, W = 0.6, L = 0.15
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__nfactor_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_57=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 058, W = 0.61, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__nfactor_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_58=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 059, W = 0.65, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__nfactor_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_59=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 060, W = 0.65, L = 0.18
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__nfactor_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_60=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 061, W = 0.65, L = 0.25
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__nfactor_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_61=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 062, W = 0.65, L = 0.5
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__nfactor_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_62=0.0
.include "sky130_fd_pr__nfet_01v8.pm3.spice"
