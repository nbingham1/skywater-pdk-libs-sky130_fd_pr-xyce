* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* statistics {
* 	mismatch {
*     	}
*         process {
* 		vary sky130_fd_pr__res_xhigh_po__var_mult dist=gauss std=0.025
* 		vary sky130_fd_pr__res_high_po__var       dist=gauss std=0.025
*         }
* }
.subckt sky130_fd_pr__res_xhigh_po_1p41 r0 r1 b
.param w=1.41 l=5 mult=1.0
Xsky130_fd_pr__res_xhigh_po_1p41 r0 r1 b sky130_fd_pr__res_xhigh_po__base w={w} l={l} mult={mult}
.ends sky130_fd_pr__res_xhigh_po_1p41
