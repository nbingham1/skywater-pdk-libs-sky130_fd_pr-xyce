* SKY130 Spice File.
* Number of bins: 1
* 9 parameters
.param
+  sky130_fd_bs_flash__special_sonosfet_original__tox_mult=1.0
+  sky130_fd_bs_flash__special_sonosfet_original__ajunction_mult=1.0
+  sky130_fd_bs_flash__special_sonosfet_original__pjunction_mult=1.0
+  sky130_fd_bs_flash__special_sonosfet_original__overlap_mult=1.0
+  sky130_fd_bs_flash__special_sonosfet_original__lint_diff=0.0
+  sky130_fd_bs_flash__special_sonosfet_original__wint_diff=0.0
+  sky130_fd_bs_flash__special_sonosfet_original__dlc_diff=0.0
+  sky130_fd_bs_flash__special_sonosfet_original__dwc_diff=0.0
*
* sky130_fd_bs_flash__special_sonosfet_original, Bin 000, W = 0.45, L = 0.22
* ------------------------------------
+  sky130_fd_bs_flash__special_sonosfet_original__rdsw_diff_0=0.0
+  sky130_fd_bs_flash__special_sonosfet_original__vth0_diff_0=-1.6077
+  sky130_fd_bs_flash__special_sonosfet_original__u0_diff_0=-4.4130e-3
+  sky130_fd_bs_flash__special_sonosfet_original__vsat_diff_0=0.0
+  sky130_fd_bs_flash__special_sonosfet_original__voff_diff_0=0.0
+  sky130_fd_bs_flash__special_sonosfet_original__k2_diff_0=0.0
+  sky130_fd_bs_flash__special_sonosfet_original__nfactor_diff_0=6.4427e-2
+  sky130_fd_bs_flash__special_sonosfet_original__kt1_diff_0=-3.5697e-1
*
* sky130_fd_bs_flash__special_sonosfet_original, Bin 001, W = 1.00, L = 0.50
* ------------------------------------
+  sky130_fd_bs_flash__special_sonosfet_original__k2_diff_1=0.0
+  sky130_fd_bs_flash__special_sonosfet_original__vth0_diff_1=-1.3466
+  sky130_fd_bs_flash__special_sonosfet_original__vsat_diff_1=0.0
+  sky130_fd_bs_flash__special_sonosfet_original__kt1_diff_1=-3.1940e-2
+  sky130_fd_bs_flash__special_sonosfet_original__u0_diff_1=-2.0e-3
+  sky130_fd_bs_flash__special_sonosfet_original__nfactor_diff_1=-5.1568e-1
+  sky130_fd_bs_flash__special_sonosfet_original__rdsw_diff_1=0.0
+  sky130_fd_bs_flash__special_sonosfet_original__voff_diff_1=0.0
*
* sky130_fd_bs_flash__special_sonosfet_original, Bin 002, W = 0.35, L = 0.15
* ------------------------------------
+  sky130_fd_bs_flash__special_sonosfet_original__rdsw_diff_2=0.0
+  sky130_fd_bs_flash__special_sonosfet_original__vth0_diff_2=-1.3168
+  sky130_fd_bs_flash__special_sonosfet_original__u0_diff_2=1.4377e-3
+  sky130_fd_bs_flash__special_sonosfet_original__vsat_diff_2=0.0
+  sky130_fd_bs_flash__special_sonosfet_original__voff_diff_2=-3.2704e-1
+  sky130_fd_bs_flash__special_sonosfet_original__k2_diff_2=0.0
+  sky130_fd_bs_flash__special_sonosfet_original__nfactor_diff_2=2.2633
+  sky130_fd_bs_flash__special_sonosfet_original__kt1_diff_2=-6.2632e-1
