* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 49
.param
+  sky130_fd_pr__nfet_g5v0d10v5__toxe_mult=0.94
+  sky130_fd_pr__nfet_g5v0d10v5__rshn_mult=1.0
+  sky130_fd_pr__nfet_g5v0d10v5__overlap_mult=0.76246
+  sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult=8.1753e-1
+  sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult=7.7786e-1
+  sky130_fd_pr__nfet_g5v0d10v5__lint_diff=1.7325e-8
+  sky130_fd_pr__nfet_g5v0d10v5__wint_diff=-3.2175e-8
+  sky130_fd_pr__nfet_g5v0d10v5__dlc_diff=1.7325e-8
+  sky130_fd_pr__nfet_g5v0d10v5__dwc_diff=-3.2175e-8
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 000, W = 10.0, L = 0.5
* -------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_0=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_0=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_0=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_0=-0.001744
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_0=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_0=0.00067346
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_0=-0.11533
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_0=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_0=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_0=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_0=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_0=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_0=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_0=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_0=-7.2729e-13
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_0=-10837.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_0=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_0=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_0=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_0=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_0=0.017751
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_0=-8.9194e-20
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_0=0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 001, W = 15.0, L = 1.0
* -------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_1=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_1=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_1=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_1=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_1=0.0065028
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_1=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_1=-0.00072595
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_1=-0.03773
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_1=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_1=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_1=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_1=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_1=-0.17178
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_1=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_1=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_1=-2.9245e-12
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_1=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_1=0.096329
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_1=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_1=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_1=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_1=0.22524
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_1=-5.5898e-19
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 002, W = 15.0, L = 0.5
* -------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_2=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_2=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_2=0.012894
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_2=-2.1053e-19
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_2=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_2=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_2=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_2=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_2=-0.0025359
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_2=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_2=0.0018816
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_2=-0.10296
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_2=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_2=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_2=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_2=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_2=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_2=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_2=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_2=-6.098e-12
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_2=-6890.7
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_2=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_2=0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 003, W = 1.5, L = 1.0
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_3=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_3=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_3=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_3=0.45157
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_3=-2.8366e-19
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_3=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_3=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_3=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_3=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_3=-0.0024725
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_3=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_3=-0.0031377
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_3=-0.067755
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_3=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_3=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_3=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_3=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_3=-0.11561
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_3=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_3=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_3=3.524e-12
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_3=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_3=0.041256
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 004, W = 1.5, L = 2.0
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_4=0.0010053
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_4=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_4=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_4=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_4=0.42135
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_4=-2.4973e-19
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_4=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_4=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_4=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_4=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_4=-0.012359
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_4=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_4=-0.0025723
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_4=-0.042901
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_4=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_4=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_4=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_4=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_4=-0.019831
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_4=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_4=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_4=2.6852e-12
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_4=0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 005, W = 1.5, L = 4.0
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_5=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_5=2.0835e-12
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_5=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_5=0.0022408
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_5=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_5=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_5=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_5=-1.6048e-19
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_5=0.49358
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_5=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_5=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_5=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_5=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_5=-0.015725
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_5=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_5=-0.0016407
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_5=-0.023862
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_5=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_5=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_5=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_5=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_5=-0.018345
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_5=0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 006, W = 1.5, L = 0.5
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_6=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_6=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_6=9.6095e-12
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_6=-17518.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_6=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_6=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_6=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_6=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_6=2.1831e-19
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_6=0.63002
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_6=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_6=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_6=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_6=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_6=0.0086273
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_6=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_6=-0.0017875
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_6=-0.14935
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_6=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_6=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_6=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_6=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_6=0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 007, W = 1.0, L = 1.0
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_7=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_7=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_7=-0.53824
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_7=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_7=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_7=9.0617e-11
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_7=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_7=-0.59992
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_7=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_7=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_7=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_7=-4.0753e-20
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_7=0.51381
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_7=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_7=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_7=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_7=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_7=0.005737
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_7=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_7=-0.00061823
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_7=-0.050984
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_7=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_7=0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 008, W = 1.0, L = 2.0
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_8=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_8=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_8=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_8=-0.045086
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_8=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_8=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_8=2.8087e-12
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_8=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_8=0.0065931
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_8=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_8=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_8=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_8=3.9997e-20
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_8=0.51123
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_8=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_8=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_8=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_8=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_8=-0.01817
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_8=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_8=-0.00080585
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_8=-0.040224
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_8=0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 009, W = 1.0, L = 4.0
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_9=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_9=-0.0012822
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_9=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_9=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_9=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_9=-0.05098
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_9=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_9=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_9=1.4474e-12
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_9=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_9=0.0068253
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_9=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_9=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_9=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_9=-1.5723e-19
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_9=0.50278
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_9=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_9=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_9=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_9=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_9=-0.011513
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_9=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_9=-0.029678
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 010, W = 1.0, L = 8.0
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_10=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_10=0.0033427
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_10=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_10=-0.00063338
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_10=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_10=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_10=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_10=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_10=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_10=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_10=-0.020704
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_10=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_10=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_10=-0.02653
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_10=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_10=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_10=-0.013333
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_10=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_10=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_10=0.62425
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_10=1.0675e-12
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_10=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_10=3.155e-20
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 011, W = 1.0, L = 0.5
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_11=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_11=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_11=6.1171e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_11=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_11=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_11=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_11=-0.0015314
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_11=-16625.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_11=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_11=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_11=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_11=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_11=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_11=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_11=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_11=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_11=-0.12897
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_11=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_11=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_11=0.012032
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_11=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_11=0.72734
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_11=1.6344e-11
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 012, W = 1.0, L = 0.6
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_12=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_12=0.6374
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_12=5.7445e-12
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_12=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_12=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_12=2.1575e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_12=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_12=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_12=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_12=-0.00080036
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_12=-16866.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_12=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_12=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_12=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_12=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_12=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_12=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_12=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_12=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_12=-0.096744
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_12=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_12=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_12=0.00028865
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 013, W = 1.0, L = 0.8
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_13=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_13=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_13=-0.0036231
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_13=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_13=0.52162
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_13=5.462e-12
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_13=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_13=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_13=1.5753e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_13=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_13=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_13=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_13=-0.0011108
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_13=-15059.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_13=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_13=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_13=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_13=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_13=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_13=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_13=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_13=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_13=-0.050378
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 014, W = 20.0, L = 1.0
* -------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_14=-0.033499
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_14=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_14=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_14=0.0059175
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_14=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_14=0.22163
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_14=-1.7474e-13
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_14=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_14=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_14=-5.8145e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_14=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_14=0.043819
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_14=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_14=-0.0003715
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_14=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_14=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_14=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_14=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_14=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_14=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_14=-0.084668
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_14=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_14=0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 015, W = 20.0, L = 0.5
* -------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_15=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_15=-0.10402
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_15=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_15=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_15=-0.0066134
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_15=-0.07294
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_15=-3.1989e-12
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_15=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_15=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_15=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_15=-1.1952e-18
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_15=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_15=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_15=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_15=-0.0011793
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_15=-12316.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_15=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_15=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_15=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_15=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_15=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_15=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_15=0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 016, W = 3.0, L = 1.0
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_16=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_16=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_16=-0.046379
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_16=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_16=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_16=-0.0029649
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_16=0.31805
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_16=5.1967e-12
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_16=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_16=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_16=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_16=-2.5784e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_16=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_16=0.037966
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_16=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_16=-0.0027377
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_16=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_16=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_16=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_16=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_16=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_16=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_16=-0.10779
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 017, W = 3.0, L = 2.0
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_17=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_17=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_17=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_17=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_17=-0.04734
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_17=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_17=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_17=-0.036778
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_17=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_17=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_17=-0.012322
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_17=0.30533
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_17=3.4276e-12
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_17=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_17=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_17=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_17=-2.2984e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_17=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_17=0.0074847
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_17=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_17=-0.0021369
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_17=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_17=0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 018, W = 3.0, L = 4.0
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_18=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_18=-0.0019436
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_18=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_18=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_18=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_18=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_18=-0.015327
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_18=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_18=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_18=-0.025357
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_18=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_18=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_18=-0.016989
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_18=0.39135
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_18=2.6195e-12
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_18=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_18=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_18=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_18=-2.1799e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_18=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_18=0.0014114
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_18=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_18=0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 019, W = 3.0, L = 8.0
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_19=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_19=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_19=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_19=-0.001547
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_19=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_19=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_19=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_19=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_19=-0.0093411
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_19=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_19=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_19=-0.026953
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_19=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_19=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_19=-0.01926
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_19=0.4283
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_19=2.6177e-12
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_19=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_19=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_19=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_19=-1.1567e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_19=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_19=0.00015762
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 020, W = 3.0, L = 0.5
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_20=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_20=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_20=-0.0008493
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_20=-11352.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_20=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_20=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_20=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_20=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_20=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_20=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_20=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_20=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_20=-0.10938
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_20=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_20=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_20=0.0013192
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_20=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_20=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_20=0.41548
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_20=6.6964e-12
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_20=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_20=2.9253e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_20=0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 021, W = 3.0, L = 0.6
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_21=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_21=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_21=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_21=-0.00014915
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_21=-11412.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_21=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_21=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_21=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_21=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_21=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_21=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_21=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_21=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_21=-0.058628
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_21=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_21=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_21=-0.0042354
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_21=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_21=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_21=0.30725
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_21=4.9625e-12
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_21=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_21=3.3096e-19
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 022, W = 5.0, L = 1.0
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_22=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_22=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_22=-2.3943e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_22=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_22=0.032162
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_22=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_22=-0.0018579
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_22=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_22=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_22=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_22=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_22=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_22=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_22=-0.093515
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_22=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_22=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_22=-0.047103
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_22=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_22=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_22=0.0079029
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_22=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_22=0.2517
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_22=1.9974e-12
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 023, W = 5.0, L = 2.0
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_23=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_23=0.31695
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_23=4.9398e-12
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_23=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_23=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_23=-3.2795e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_23=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_23=0.00028143
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_23=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_23=-0.0030795
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_23=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_23=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_23=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_23=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_23=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_23=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_23=-0.014367
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_23=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_23=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_23=-0.032842
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_23=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_23=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_23=-0.0030642
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 024, W = 5.0, L = 4.0
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_24=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_24=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_24=-0.0067096
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_24=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_24=0.37141
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_24=4.2158e-12
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_24=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_24=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_24=-4.0315e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_24=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_24=0.001735
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_24=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_24=-0.0031364
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_24=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_24=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_24=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_24=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_24=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_24=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_24=-0.013816
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_24=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_24=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_24=-0.026088
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 025, W = 5.0, L = 8.0
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_25=-0.020915
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_25=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_25=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_25=-0.0098344
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_25=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_25=0.41226
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_25=4.1901e-12
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_25=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_25=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_25=-3.0855e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_25=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_25=0.00053738
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_25=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_25=-0.0028418
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_25=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_25=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_25=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_25=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_25=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_25=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_25=-0.0054488
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_25=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_25=0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 026, W = 5.0, L = 0.5
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_26=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_26=-0.10884
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_26=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_26=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_26=-0.0055458
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_26=0.26606
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_26=4.2929e-12
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_26=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_26=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_26=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_26=2.7713e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_26=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_26=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_26=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_26=-3.6655e-5
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_26=-10490.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_26=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_26=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_26=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_26=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_26=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_26=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_26=0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 027, W = 5.0, L = 0.6
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_27=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_27=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_27=-0.048477
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_27=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_27=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_27=0.0035792
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_27=0.2633
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_27=2.7136e-12
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_27=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_27=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_27=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_27=2.5526e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_27=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_27=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_27=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_27=0.00031269
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_27=-9644.7
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_27=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_27=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_27=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_27=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_27=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_27=0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 028, W = 5.0, L = 0.8
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_28=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_28=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_28=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_28=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_28=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_28=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_28=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_28=-0.050601
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_28=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_28=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_28=0.010605
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_28=0.2468
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_28=3.1807e-12
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_28=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_28=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_28=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_28=-1.0796e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_28=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_28=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_28=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_28=-0.0013987
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_28=-9154.7
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_28=0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 029, W = 7.0, L = 1.0
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_29=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_29=-0.0030942
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_29=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_29=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_29=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_29=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_29=-0.092123
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_29=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_29=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_29=-0.046919
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_29=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_29=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_29=0.0068682
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_29=0.24381
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_29=4.5534e-12
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_29=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_29=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_29=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_29=-4.414e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_29=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_29=0.027943
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_29=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_29=0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 030, W = 7.0, L = 2.0
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_30=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_30=-0.0038175
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_30=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_30=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_30=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_30=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_30=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_30=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_30=-0.023244
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_30=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_30=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_30=-0.033621
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_30=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_30=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_30=-0.0031254
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_30=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_30=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_30=0.30066
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_30=5.2436e-12
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_30=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_30=-5.357e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_30=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_30=0.0020451
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 031, W = 7.0, L = 4.0
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_31=0.0022363
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_31=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_31=-0.0032561
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_31=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_31=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_31=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_31=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_31=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_31=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_31=-0.016796
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_31=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_31=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_31=-0.027828
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_31=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_31=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_31=-0.0080288
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_31=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_31=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_31=0.34407
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_31=4.1919e-12
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_31=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_31=-4.5483e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_31=0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 032, W = 7.0, L = 8.0
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_32=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_32=-0.00033374
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_32=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_32=-0.0031495
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_32=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_32=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_32=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_32=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_32=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_32=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_32=-0.0063838
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_32=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_32=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_32=-0.023919
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_32=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_32=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_32=-0.0092581
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_32=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_32=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_32=0.38353
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_32=4.4861e-12
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_32=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_32=-3.862e-19
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 033, W = 7.0, L = 0.5
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_33=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_33=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_33=3.1635e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_33=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_33=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_33=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_33=0.00076765
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_33=-8082.5
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_33=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_33=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_33=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_33=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_33=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_33=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_33=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_33=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_33=-0.11157
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_33=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_33=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_33=-0.0049124
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_33=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_33=0.10731
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_33=2.5342e-12
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 034, W = 7.0, L = 0.8
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_34=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_34=0.23476
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_34=3.4845e-12
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_34=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_34=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_34=-4.3629e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_34=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_34=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_34=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_34=-0.0028047
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_34=-11258.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_34=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_34=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_34=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_34=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_34=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_34=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_34=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_34=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_34=-0.046501
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_34=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_34=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_34=0.0096808
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 035, W = 0.42, L = 1.0
* -------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_35=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_35=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_35=-0.013148
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_35=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_35=0.32428
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_35=1.2125e-11
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_35=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_35=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_35=4.7539e-20
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_35=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_35=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_35=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_35=-0.003457
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_35=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_35=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_35=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_35=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_35=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_35=2.6925e-7
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_35=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_35=-2.4215e-9
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_35=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_35=-0.12179
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 036, W = 0.42, L = 20.0
* --------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_36=-0.058622
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_36=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_36=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_36=-0.01786
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_36=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_36=0.95348
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_36=6.4917e-12
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_36=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_36=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_36=-1.8362e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_36=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_36=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_36=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_36=-0.003775
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_36=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_36=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_36=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_36=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_36=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_36=5.9604e-8
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_36=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_36=4.2551e-10
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_36=0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 037, W = 0.42, L = 2.0
* -------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_37=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_37=-0.065972
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_37=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_37=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_37=-0.019646
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_37=0.48194
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_37=7.1708e-12
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_37=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_37=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_37=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_37=-1.1404e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_37=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_37=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_37=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_37=-0.0026716
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_37=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_37=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_37=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_37=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_37=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_37=9.5177e-8
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_37=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_37=-1.5823e-9
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 038, W = 0.42, L = 4.0
* -------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_38=-3.398e-9
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_38=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_38=-0.068355
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_38=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_38=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_38=-0.016156
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_38=0.54072
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_38=1.0732e-11
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_38=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_38=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_38=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_38=-1.6411e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_38=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_38=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_38=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_38=-0.0042034
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_38=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_38=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_38=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_38=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_38=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_38=4.885e-8
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_38=0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 039, W = 0.42, L = 8.0
* -------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_39=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_39=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_39=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_39=5.7403e-8
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_39=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_39=3.3719e-8
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_39=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_39=-0.064182
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_39=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_39=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_39=-0.02017
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_39=0.72934
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_39=8.1318e-12
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_39=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_39=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_39=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_39=-3.653e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_39=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_39=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_39=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_39=-0.0041811
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_39=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_39=0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 040, W = 0.42, L = 0.5
* -------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_40=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_40=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_40=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_40=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_40=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_40=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_40=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_40=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_40=-0.14814
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_40=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_40=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_40=0.0011713
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_40=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_40=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_40=0.62698
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_40=3.7351e-12
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_40=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_40=2.2029e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_40=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_40=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_40=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_40=-0.0027234
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_40=-23997.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 041, W = 0.42, L = 0.6
* -------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_41=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_41=-0.0025844
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_41=-21982.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_41=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_41=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_41=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_41=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_41=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_41=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_41=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_41=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_41=-0.12926
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_41=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_41=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_41=-0.015942
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_41=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_41=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_41=0.47265
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_41=3.912e-12
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_41=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_41=3.6155e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_41=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_41=0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 042, W = 0.42, L = 0.8
* -------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_42=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_42=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_42=-0.0021575
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_42=-17815.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_42=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_42=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_42=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_42=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_42=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_42=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_42=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_42=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_42=-0.1332
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_42=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_42=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_42=-0.022906
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_42=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_42=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_42=0.43487
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_42=1.2974e-12
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_42=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_42=1.7324e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_42=0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 043, W = 0.75, L = 1.0
* -------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_43=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_43=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_43=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_43=-0.0015022
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_43=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_43=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_43=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_43=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_43=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_43=2.5083e-7
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_43=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_43=1.8595e-9
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_43=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_43=-0.057005
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_43=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_43=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_43=-0.00361
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_43=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_43=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_43=0.5045
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_43=5.6688e-12
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_43=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_43=9.2328e-20
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 044, W = 0.75, L = 2.0
* -------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_44=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_44=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_44=1.4394e-20
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_44=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_44=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_44=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_44=-0.001027
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_44=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_44=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_44=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_44=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_44=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_44=1.2039e-7
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_44=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_44=-2.0663e-10
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_44=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_44=-0.062588
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_44=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_44=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_44=-0.013153
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_44=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_44=0.51157
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_44=3.7152e-12
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 045, W = 0.75, L = 4.0
* -------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_45=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_45=0.60809
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_45=2.6165e-12
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_45=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_45=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_45=-2.3003e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_45=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_45=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_45=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_45=-0.0020521
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_45=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_45=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_45=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_45=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_45=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_45=1.597e-7
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_45=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_45=-1.606e-10
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_45=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_45=-0.037911
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_45=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_45=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_45=-0.018074
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 046, W = 0.75, L = 0.5
* -------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_46=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_46=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_46=0.0035731
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_46=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_46=0.68272
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_46=1.293e-11
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_46=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_46=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_46=6.3502e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_46=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_46=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_46=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_46=-0.001157
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_46=-17789.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_46=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_46=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_46=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_46=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_46=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_46=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_46=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_46=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_46=-0.12821
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 047, W = 0.75, L = 0.8
* -------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_47=-0.064169
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_47=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_47=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_47=-0.00085911
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_47=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_47=0.60536
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_47=4.9518e-12
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_47=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_47=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_47=8.6671e-20
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_47=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_47=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_47=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_47=-0.0011573
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_47=-17521.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_47=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_47=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_47=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_47=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_47=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_47=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_47=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_47=0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 048, W = 0.7, L = 0.6
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_48=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_48=-0.096097
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_48=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_48=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_48=5.4148e-5
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_48=0.7055
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_48=8.8919e-12
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_48=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_48=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_48=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_48=2.3132e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_48=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_48=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_48=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_48=-0.0018033
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_48=-20000.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_48=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_48=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_48=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_48=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_48=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_48=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_48=0.0
.include "sky130_fd_pr__nfet_g5v0d10v5.pm3.spice"
