* Pwell-isolated Transistor Vth and I-V characteristic

* Include SkyWater sky130 device models
.lib "../../../models/sky130.lib.spice" tt
.include "../../nfet_20v0/sky130_fd_pr__nfet_20v0__tt_discrete.corner.spice"
.include "../sky130_fd_pr__nfet_20v0_nvt_iso__tt_discrete.corner.spice"

* Gate bias
Rg 1 2 680
X1 3 2 0 4 0 sky130_fd_pr__nfet_20v0_nvt_iso W=20 L=1 M=1
Rd 3 4 100

* DC source for current measure
Vid 5 4 DC 0V
Vgb 1 0 DC 0V
Vdd 5 0 DC 3.3V

.control
* Sweep Vds from 0 to 1.8V
dc Vdd 0 1.8 0.01 Vgb 0 1.2 0.01
wrdata sky130_fd_pr__nfet_20v0_nvt_iso__iv.data Vid#branch V ( 1 ) V ( 3 )

* Sweep Vgs from 0 to 1.2V
dc Vgb 0 1.2 0.01
+ # Find threshold
let ih=Vid#branch[98]
let il=Vid#branch[85]
let vh=V(2)[98]
let vl=V(2)[85]
let vth=((vl - vh ) / ( ih - il ) ) * ih vh
echo threshold voltage
print vth
quit
.endc
.end
