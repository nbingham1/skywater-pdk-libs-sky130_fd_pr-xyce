* SKY130 Spice File.
.param globalk=1
.param localkswitch=1
.param capunits='1.0*1e-6'
.param
+  mcp1f_ca_w_0_150_s_0_210=1.55e-04 mcp1f_cc_w_0_150_s_0_210=8.91e-11 mcp1f_cf_w_0_150_s_0_210=1.33e-11
+  mcp1f_ca_w_0_150_s_0_263=1.55e-04 mcp1f_cc_w_0_150_s_0_263=6.96e-11 mcp1f_cf_w_0_150_s_0_263=1.63e-11
+  mcp1f_ca_w_0_150_s_0_315=1.55e-04 mcp1f_cc_w_0_150_s_0_315=5.79e-11 mcp1f_cf_w_0_150_s_0_315=1.91e-11
+  mcp1f_ca_w_0_150_s_0_420=1.55e-04 mcp1f_cc_w_0_150_s_0_420=4.29e-11 mcp1f_cf_w_0_150_s_0_420=2.41e-11
+  mcp1f_ca_w_0_150_s_0_525=1.55e-04 mcp1f_cc_w_0_150_s_0_525=3.42e-11 mcp1f_cf_w_0_150_s_0_525=2.82e-11
+  mcp1f_ca_w_0_150_s_0_630=1.55e-04 mcp1f_cc_w_0_150_s_0_630=2.83e-11 mcp1f_cf_w_0_150_s_0_630=3.16e-11
+  mcp1f_ca_w_0_150_s_0_840=1.55e-04 mcp1f_cc_w_0_150_s_0_840=2.04e-11 mcp1f_cf_w_0_150_s_0_840=3.71e-11
+  mcp1f_ca_w_0_150_s_1_260=1.55e-04 mcp1f_cc_w_0_150_s_1_260=1.15e-11 mcp1f_cf_w_0_150_s_1_260=4.44e-11
+  mcp1f_ca_w_0_150_s_2_310=1.55e-04 mcp1f_cc_w_0_150_s_2_310=4.85e-12 mcp1f_cf_w_0_150_s_2_310=5.06e-11
+  mcp1f_ca_w_0_150_s_5_250=1.55e-04 mcp1f_cc_w_0_150_s_5_250=1.10e-12 mcp1f_cf_w_0_150_s_5_250=5.43e-11
+  mcp1f_ca_w_1_200_s_0_210=1.55e-04 mcp1f_cc_w_1_200_s_0_210=1.08e-10 mcp1f_cf_w_1_200_s_0_210=1.32e-11
+  mcp1f_ca_w_1_200_s_0_263=1.55e-04 mcp1f_cc_w_1_200_s_0_263=8.71e-11 mcp1f_cf_w_1_200_s_0_263=1.63e-11
+  mcp1f_ca_w_1_200_s_0_315=1.55e-04 mcp1f_cc_w_1_200_s_0_315=7.40e-11 mcp1f_cf_w_1_200_s_0_315=1.91e-11
+  mcp1f_ca_w_1_200_s_0_420=1.55e-04 mcp1f_cc_w_1_200_s_0_420=5.78e-11 mcp1f_cf_w_1_200_s_0_420=2.40e-11
+  mcp1f_ca_w_1_200_s_0_525=1.55e-04 mcp1f_cc_w_1_200_s_0_525=4.76e-11 mcp1f_cf_w_1_200_s_0_525=2.82e-11
+  mcp1f_ca_w_1_200_s_0_630=1.55e-04 mcp1f_cc_w_1_200_s_0_630=4.07e-11 mcp1f_cf_w_1_200_s_0_630=3.18e-11
+  mcp1f_ca_w_1_200_s_0_840=1.55e-04 mcp1f_cc_w_1_200_s_0_840=3.14e-11 mcp1f_cf_w_1_200_s_0_840=3.76e-11
+  mcp1f_ca_w_1_200_s_1_260=1.55e-04 mcp1f_cc_w_1_200_s_1_260=2.11e-11 mcp1f_cf_w_1_200_s_1_260=4.54e-11
+  mcp1f_ca_w_1_200_s_2_310=1.55e-04 mcp1f_cc_w_1_200_s_2_310=1.03e-11 mcp1f_cf_w_1_200_s_2_310=5.50e-11
+  mcp1f_ca_w_1_200_s_5_250=1.55e-04 mcp1f_cc_w_1_200_s_5_250=3.25e-12 mcp1f_cf_w_1_200_s_5_250=6.19e-11
+  mcl1f_ca_w_0_170_s_0_180=4.97e-05 mcl1f_cc_w_0_170_s_0_180=1.01e-10 mcl1f_cf_w_0_170_s_0_180=3.56e-12
+  mcl1f_ca_w_0_170_s_0_225=4.97e-05 mcl1f_cc_w_0_170_s_0_225=8.20e-11 mcl1f_cf_w_0_170_s_0_225=4.63e-12
+  mcl1f_ca_w_0_170_s_0_270=4.97e-05 mcl1f_cc_w_0_170_s_0_270=7.04e-11 mcl1f_cf_w_0_170_s_0_270=5.66e-12
+  mcl1f_ca_w_0_170_s_0_360=4.97e-05 mcl1f_cc_w_0_170_s_0_360=5.55e-11 mcl1f_cf_w_0_170_s_0_360=7.72e-12
+  mcl1f_ca_w_0_170_s_0_450=4.97e-05 mcl1f_cc_w_0_170_s_0_450=4.65e-11 mcl1f_cf_w_0_170_s_0_450=9.60e-12
+  mcl1f_ca_w_0_170_s_0_540=4.97e-05 mcl1f_cc_w_0_170_s_0_540=3.97e-11 mcl1f_cf_w_0_170_s_0_540=1.17e-11
+  mcl1f_ca_w_0_170_s_0_720=4.97e-05 mcl1f_cc_w_0_170_s_0_720=3.10e-11 mcl1f_cf_w_0_170_s_0_720=1.51e-11
+  mcl1f_ca_w_0_170_s_1_080=4.97e-05 mcl1f_cc_w_0_170_s_1_080=2.08e-11 mcl1f_cf_w_0_170_s_1_080=2.07e-11
+  mcl1f_ca_w_0_170_s_1_980=4.97e-05 mcl1f_cc_w_0_170_s_1_980=1.03e-11 mcl1f_cf_w_0_170_s_1_980=2.88e-11
+  mcl1f_ca_w_0_170_s_4_500=4.97e-05 mcl1f_cc_w_0_170_s_4_500=2.87e-12 mcl1f_cf_w_0_170_s_4_500=3.57e-11
+  mcl1f_ca_w_1_360_s_0_180=4.97e-05 mcl1f_cc_w_1_360_s_0_180=1.21e-10 mcl1f_cf_w_1_360_s_0_180=3.56e-12
+  mcl1f_ca_w_1_360_s_0_225=4.97e-05 mcl1f_cc_w_1_360_s_0_225=1.01e-10 mcl1f_cf_w_1_360_s_0_225=4.62e-12
+  mcl1f_ca_w_1_360_s_0_270=4.97e-05 mcl1f_cc_w_1_360_s_0_270=8.77e-11 mcl1f_cf_w_1_360_s_0_270=5.66e-12
+  mcl1f_ca_w_1_360_s_0_360=4.97e-05 mcl1f_cc_w_1_360_s_0_360=7.11e-11 mcl1f_cf_w_1_360_s_0_360=7.69e-12
+  mcl1f_ca_w_1_360_s_0_450=4.97e-05 mcl1f_cc_w_1_360_s_0_450=6.07e-11 mcl1f_cf_w_1_360_s_0_450=9.64e-12
+  mcl1f_ca_w_1_360_s_0_540=4.97e-05 mcl1f_cc_w_1_360_s_0_540=5.32e-11 mcl1f_cf_w_1_360_s_0_540=1.15e-11
+  mcl1f_ca_w_1_360_s_0_720=4.97e-05 mcl1f_cc_w_1_360_s_0_720=4.30e-11 mcl1f_cf_w_1_360_s_0_720=1.50e-11
+  mcl1f_ca_w_1_360_s_1_080=4.97e-05 mcl1f_cc_w_1_360_s_1_080=3.12e-11 mcl1f_cf_w_1_360_s_1_080=2.08e-11
+  mcl1f_ca_w_1_360_s_1_980=4.97e-05 mcl1f_cc_w_1_360_s_1_980=1.74e-11 mcl1f_cf_w_1_360_s_1_980=3.06e-11
+  mcl1f_ca_w_1_360_s_4_500=4.97e-05 mcl1f_cc_w_1_360_s_4_500=6.15e-12 mcl1f_cf_w_1_360_s_4_500=4.08e-11
+  mcl1d_ca_w_0_170_s_0_180=7.09e-05 mcl1d_cc_w_0_170_s_0_180=9.83e-11 mcl1d_cf_w_0_170_s_0_180=5.04e-12
+  mcl1d_ca_w_0_170_s_0_225=7.09e-05 mcl1d_cc_w_0_170_s_0_225=7.93e-11 mcl1d_cf_w_0_170_s_0_225=6.52e-12
+  mcl1d_ca_w_0_170_s_0_270=7.09e-05 mcl1d_cc_w_0_170_s_0_270=6.75e-11 mcl1d_cf_w_0_170_s_0_270=7.95e-12
+  mcl1d_ca_w_0_170_s_0_360=7.09e-05 mcl1d_cc_w_0_170_s_0_360=5.24e-11 mcl1d_cf_w_0_170_s_0_360=1.08e-11
+  mcl1d_ca_w_0_170_s_0_450=7.09e-05 mcl1d_cc_w_0_170_s_0_450=4.33e-11 mcl1d_cf_w_0_170_s_0_450=1.33e-11
+  mcl1d_ca_w_0_170_s_0_540=7.09e-05 mcl1d_cc_w_0_170_s_0_540=3.63e-11 mcl1d_cf_w_0_170_s_0_540=1.60e-11
+  mcl1d_ca_w_0_170_s_0_720=7.09e-05 mcl1d_cc_w_0_170_s_0_720=2.74e-11 mcl1d_cf_w_0_170_s_0_720=2.03e-11
+  mcl1d_ca_w_0_170_s_1_080=7.09e-05 mcl1d_cc_w_0_170_s_1_080=1.74e-11 mcl1d_cf_w_0_170_s_1_080=2.68e-11
+  mcl1d_ca_w_0_170_s_1_980=7.09e-05 mcl1d_cc_w_0_170_s_1_980=7.88e-12 mcl1d_cf_w_0_170_s_1_980=3.49e-11
+  mcl1d_ca_w_0_170_s_4_500=7.09e-05 mcl1d_cc_w_0_170_s_4_500=2.05e-12 mcl1d_cf_w_0_170_s_4_500=4.05e-11
+  mcl1d_ca_w_1_360_s_0_180=7.09e-05 mcl1d_cc_w_1_360_s_0_180=1.17e-10 mcl1d_cf_w_1_360_s_0_180=5.04e-12
+  mcl1d_ca_w_1_360_s_0_225=7.09e-05 mcl1d_cc_w_1_360_s_0_225=9.68e-11 mcl1d_cf_w_1_360_s_0_225=6.51e-12
+  mcl1d_ca_w_1_360_s_0_270=7.09e-05 mcl1d_cc_w_1_360_s_0_270=8.38e-11 mcl1d_cf_w_1_360_s_0_270=7.96e-12
+  mcl1d_ca_w_1_360_s_0_360=7.09e-05 mcl1d_cc_w_1_360_s_0_360=6.72e-11 mcl1d_cf_w_1_360_s_0_360=1.07e-11
+  mcl1d_ca_w_1_360_s_0_450=7.09e-05 mcl1d_cc_w_1_360_s_0_450=5.68e-11 mcl1d_cf_w_1_360_s_0_450=1.33e-11
+  mcl1d_ca_w_1_360_s_0_540=7.09e-05 mcl1d_cc_w_1_360_s_0_540=4.93e-11 mcl1d_cf_w_1_360_s_0_540=1.58e-11
+  mcl1d_ca_w_1_360_s_0_720=7.09e-05 mcl1d_cc_w_1_360_s_0_720=3.92e-11 mcl1d_cf_w_1_360_s_0_720=2.02e-11
+  mcl1d_ca_w_1_360_s_1_080=7.09e-05 mcl1d_cc_w_1_360_s_1_080=2.76e-11 mcl1d_cf_w_1_360_s_1_080=2.71e-11
+  mcl1d_ca_w_1_360_s_1_980=7.09e-05 mcl1d_cc_w_1_360_s_1_980=1.46e-11 mcl1d_cf_w_1_360_s_1_980=3.75e-11
+  mcl1d_ca_w_1_360_s_4_500=7.09e-05 mcl1d_cc_w_1_360_s_4_500=4.95e-12 mcl1d_cf_w_1_360_s_4_500=4.66e-11
+  mcl1p1_ca_w_0_170_s_0_180=1.74e-04 mcl1p1_cc_w_0_170_s_0_180=9.03e-11 mcl1p1_cf_w_0_170_s_0_180=1.18e-11
+  mcl1p1_ca_w_0_170_s_0_225=1.74e-04 mcl1p1_cc_w_0_170_s_0_225=7.11e-11 mcl1p1_cf_w_0_170_s_0_225=1.51e-11
+  mcl1p1_ca_w_0_170_s_0_270=1.74e-04 mcl1p1_cc_w_0_170_s_0_270=5.91e-11 mcl1p1_cf_w_0_170_s_0_270=1.81e-11
+  mcl1p1_ca_w_0_170_s_0_360=1.74e-04 mcl1p1_cc_w_0_170_s_0_360=4.36e-11 mcl1p1_cf_w_0_170_s_0_360=2.37e-11
+  mcl1p1_ca_w_0_170_s_0_450=1.74e-04 mcl1p1_cc_w_0_170_s_0_450=3.44e-11 mcl1p1_cf_w_0_170_s_0_450=2.82e-11
+  mcl1p1_ca_w_0_170_s_0_540=1.74e-04 mcl1p1_cc_w_0_170_s_0_540=2.72e-11 mcl1p1_cf_w_0_170_s_0_540=3.27e-11
+  mcl1p1_ca_w_0_170_s_0_720=1.74e-04 mcl1p1_cc_w_0_170_s_0_720=1.87e-11 mcl1p1_cf_w_0_170_s_0_720=3.88e-11
+  mcl1p1_ca_w_0_170_s_1_080=1.74e-04 mcl1p1_cc_w_0_170_s_1_080=1.03e-11 mcl1p1_cf_w_0_170_s_1_080=4.61e-11
+  mcl1p1_ca_w_0_170_s_1_980=1.74e-04 mcl1p1_cc_w_0_170_s_1_980=4.00e-12 mcl1p1_cf_w_0_170_s_1_980=5.21e-11
+  mcl1p1_ca_w_0_170_s_4_500=1.74e-04 mcl1p1_cc_w_0_170_s_4_500=1.00e-12 mcl1p1_cf_w_0_170_s_4_500=5.51e-11
+  mcl1p1_ca_w_1_360_s_0_180=1.74e-04 mcl1p1_cc_w_1_360_s_0_180=1.08e-10 mcl1p1_cf_w_1_360_s_0_180=1.20e-11
+  mcl1p1_ca_w_1_360_s_0_225=1.74e-04 mcl1p1_cc_w_1_360_s_0_225=8.78e-11 mcl1p1_cf_w_1_360_s_0_225=1.52e-11
+  mcl1p1_ca_w_1_360_s_0_270=1.74e-04 mcl1p1_cc_w_1_360_s_0_270=7.46e-11 mcl1p1_cf_w_1_360_s_0_270=1.82e-11
+  mcl1p1_ca_w_1_360_s_0_360=1.74e-04 mcl1p1_cc_w_1_360_s_0_360=5.80e-11 mcl1p1_cf_w_1_360_s_0_360=2.37e-11
+  mcl1p1_ca_w_1_360_s_0_450=1.74e-04 mcl1p1_cc_w_1_360_s_0_450=4.77e-11 mcl1p1_cf_w_1_360_s_0_450=2.85e-11
+  mcl1p1_ca_w_1_360_s_0_540=1.74e-04 mcl1p1_cc_w_1_360_s_0_540=4.04e-11 mcl1p1_cf_w_1_360_s_0_540=3.26e-11
+  mcl1p1_ca_w_1_360_s_0_720=1.74e-04 mcl1p1_cc_w_1_360_s_0_720=3.07e-11 mcl1p1_cf_w_1_360_s_0_720=3.91e-11
+  mcl1p1_ca_w_1_360_s_1_080=1.74e-04 mcl1p1_cc_w_1_360_s_1_080=2.03e-11 mcl1p1_cf_w_1_360_s_1_080=4.75e-11
+  mcl1p1_ca_w_1_360_s_1_980=1.74e-04 mcl1p1_cc_w_1_360_s_1_980=9.95e-12 mcl1p1_cf_w_1_360_s_1_980=5.71e-11
+  mcl1p1_ca_w_1_360_s_4_500=1.74e-04 mcl1p1_cc_w_1_360_s_4_500=3.20e-12 mcl1p1_cf_w_1_360_s_4_500=6.37e-11
+  mcm1f_ca_w_0_140_s_0_140=3.57e-05 mcm1f_cc_w_0_140_s_0_140=1.30e-10 mcm1f_cf_w_0_140_s_0_140=1.93e-12
+  mcm1f_ca_w_0_140_s_0_175=3.57e-05 mcm1f_cc_w_0_140_s_0_175=1.24e-10 mcm1f_cf_w_0_140_s_0_175=2.55e-12
+  mcm1f_ca_w_0_140_s_0_210=3.57e-05 mcm1f_cc_w_0_140_s_0_210=1.17e-10 mcm1f_cf_w_0_140_s_0_210=3.16e-12
+  mcm1f_ca_w_0_140_s_0_280=3.57e-05 mcm1f_cc_w_0_140_s_0_280=1.00e-10 mcm1f_cf_w_0_140_s_0_280=4.38e-12
+  mcm1f_ca_w_0_140_s_0_350=3.57e-05 mcm1f_cc_w_0_140_s_0_350=8.56e-11 mcm1f_cf_w_0_140_s_0_350=5.56e-12
+  mcm1f_ca_w_0_140_s_0_420=3.57e-05 mcm1f_cc_w_0_140_s_0_420=7.44e-11 mcm1f_cf_w_0_140_s_0_420=6.77e-12
+  mcm1f_ca_w_0_140_s_0_560=3.57e-05 mcm1f_cc_w_0_140_s_0_560=5.85e-11 mcm1f_cf_w_0_140_s_0_560=8.95e-12
+  mcm1f_ca_w_0_140_s_0_840=3.57e-05 mcm1f_cc_w_0_140_s_0_840=4.17e-11 mcm1f_cf_w_0_140_s_0_840=1.30e-11
+  mcm1f_ca_w_0_140_s_1_540=3.57e-05 mcm1f_cc_w_0_140_s_1_540=2.38e-11 mcm1f_cf_w_0_140_s_1_540=2.13e-11
+  mcm1f_ca_w_0_140_s_3_500=3.57e-05 mcm1f_cc_w_0_140_s_3_500=8.73e-12 mcm1f_cf_w_0_140_s_3_500=3.30e-11
+  mcm1f_ca_w_1_120_s_0_140=3.57e-05 mcm1f_cc_w_1_120_s_0_140=1.54e-10 mcm1f_cf_w_1_120_s_0_140=1.99e-12
+  mcm1f_ca_w_1_120_s_0_175=3.57e-05 mcm1f_cc_w_1_120_s_0_175=1.46e-10 mcm1f_cf_w_1_120_s_0_175=2.62e-12
+  mcm1f_ca_w_1_120_s_0_210=3.57e-05 mcm1f_cc_w_1_120_s_0_210=1.38e-10 mcm1f_cf_w_1_120_s_0_210=3.23e-12
+  mcm1f_ca_w_1_120_s_0_280=3.57e-05 mcm1f_cc_w_1_120_s_0_280=1.18e-10 mcm1f_cf_w_1_120_s_0_280=4.44e-12
+  mcm1f_ca_w_1_120_s_0_350=3.57e-05 mcm1f_cc_w_1_120_s_0_350=1.02e-10 mcm1f_cf_w_1_120_s_0_350=5.64e-12
+  mcm1f_ca_w_1_120_s_0_420=3.57e-05 mcm1f_cc_w_1_120_s_0_420=8.95e-11 mcm1f_cf_w_1_120_s_0_420=6.81e-12
+  mcm1f_ca_w_1_120_s_0_560=3.57e-05 mcm1f_cc_w_1_120_s_0_560=7.17e-11 mcm1f_cf_w_1_120_s_0_560=9.04e-12
+  mcm1f_ca_w_1_120_s_0_840=3.57e-05 mcm1f_cc_w_1_120_s_0_840=5.23e-11 mcm1f_cf_w_1_120_s_0_840=1.32e-11
+  mcm1f_ca_w_1_120_s_1_540=3.57e-05 mcm1f_cc_w_1_120_s_1_540=3.15e-11 mcm1f_cf_w_1_120_s_1_540=2.18e-11
+  mcm1f_ca_w_1_120_s_3_500=3.57e-05 mcm1f_cc_w_1_120_s_3_500=1.31e-11 mcm1f_cf_w_1_120_s_3_500=3.50e-11
+  mcm1d_ca_w_0_140_s_0_140=4.54e-05 mcm1d_cc_w_0_140_s_0_140=1.29e-10 mcm1d_cf_w_0_140_s_0_140=2.45e-12
+  mcm1d_ca_w_0_140_s_0_175=4.54e-05 mcm1d_cc_w_0_140_s_0_175=1.23e-10 mcm1d_cf_w_0_140_s_0_175=3.23e-12
+  mcm1d_ca_w_0_140_s_0_210=4.54e-05 mcm1d_cc_w_0_140_s_0_210=1.16e-10 mcm1d_cf_w_0_140_s_0_210=4.02e-12
+  mcm1d_ca_w_0_140_s_0_280=4.54e-05 mcm1d_cc_w_0_140_s_0_280=9.85e-11 mcm1d_cf_w_0_140_s_0_280=5.56e-12
+  mcm1d_ca_w_0_140_s_0_350=4.54e-05 mcm1d_cc_w_0_140_s_0_350=8.39e-11 mcm1d_cf_w_0_140_s_0_350=7.05e-12
+  mcm1d_ca_w_0_140_s_0_420=4.54e-05 mcm1d_cc_w_0_140_s_0_420=7.24e-11 mcm1d_cf_w_0_140_s_0_420=8.53e-12
+  mcm1d_ca_w_0_140_s_0_560=4.54e-05 mcm1d_cc_w_0_140_s_0_560=5.65e-11 mcm1d_cf_w_0_140_s_0_560=1.12e-11
+  mcm1d_ca_w_0_140_s_0_840=4.54e-05 mcm1d_cc_w_0_140_s_0_840=3.95e-11 mcm1d_cf_w_0_140_s_0_840=1.62e-11
+  mcm1d_ca_w_0_140_s_1_540=4.54e-05 mcm1d_cc_w_0_140_s_1_540=2.16e-11 mcm1d_cf_w_0_140_s_1_540=2.57e-11
+  mcm1d_ca_w_0_140_s_3_500=4.54e-05 mcm1d_cc_w_0_140_s_3_500=7.30e-12 mcm1d_cf_w_0_140_s_3_500=3.74e-11
+  mcm1d_ca_w_1_120_s_0_140=4.54e-05 mcm1d_cc_w_1_120_s_0_140=1.52e-10 mcm1d_cf_w_1_120_s_0_140=2.55e-12
+  mcm1d_ca_w_1_120_s_0_175=4.54e-05 mcm1d_cc_w_1_120_s_0_175=1.44e-10 mcm1d_cf_w_1_120_s_0_175=3.34e-12
+  mcm1d_ca_w_1_120_s_0_210=4.54e-05 mcm1d_cc_w_1_120_s_0_210=1.35e-10 mcm1d_cf_w_1_120_s_0_210=4.11e-12
+  mcm1d_ca_w_1_120_s_0_280=4.54e-05 mcm1d_cc_w_1_120_s_0_280=1.15e-10 mcm1d_cf_w_1_120_s_0_280=5.64e-12
+  mcm1d_ca_w_1_120_s_0_350=4.54e-05 mcm1d_cc_w_1_120_s_0_350=9.96e-11 mcm1d_cf_w_1_120_s_0_350=7.14e-12
+  mcm1d_ca_w_1_120_s_0_420=4.54e-05 mcm1d_cc_w_1_120_s_0_420=8.72e-11 mcm1d_cf_w_1_120_s_0_420=8.60e-12
+  mcm1d_ca_w_1_120_s_0_560=4.54e-05 mcm1d_cc_w_1_120_s_0_560=6.89e-11 mcm1d_cf_w_1_120_s_0_560=1.14e-11
+  mcm1d_ca_w_1_120_s_0_840=4.54e-05 mcm1d_cc_w_1_120_s_0_840=4.95e-11 mcm1d_cf_w_1_120_s_0_840=1.64e-11
+  mcm1d_ca_w_1_120_s_1_540=4.54e-05 mcm1d_cc_w_1_120_s_1_540=2.90e-11 mcm1d_cf_w_1_120_s_1_540=2.62e-11
+  mcm1d_ca_w_1_120_s_3_500=4.54e-05 mcm1d_cc_w_1_120_s_3_500=1.14e-11 mcm1d_cf_w_1_120_s_3_500=3.97e-11
+  mcm1p1_ca_w_0_140_s_0_140=7.32e-05 mcm1p1_cc_w_0_140_s_0_140=1.26e-10 mcm1p1_cf_w_0_140_s_0_140=3.92e-12
+  mcm1p1_ca_w_0_140_s_0_175=7.32e-05 mcm1p1_cc_w_0_140_s_0_175=1.19e-10 mcm1p1_cf_w_0_140_s_0_175=5.19e-12
+  mcm1p1_ca_w_0_140_s_0_210=7.32e-05 mcm1p1_cc_w_0_140_s_0_210=1.12e-10 mcm1p1_cf_w_0_140_s_0_210=6.44e-12
+  mcm1p1_ca_w_0_140_s_0_280=7.32e-05 mcm1p1_cc_w_0_140_s_0_280=9.46e-11 mcm1p1_cf_w_0_140_s_0_280=8.86e-12
+  mcm1p1_ca_w_0_140_s_0_350=7.32e-05 mcm1p1_cc_w_0_140_s_0_350=8.01e-11 mcm1p1_cf_w_0_140_s_0_350=1.12e-11
+  mcm1p1_ca_w_0_140_s_0_420=7.32e-05 mcm1p1_cc_w_0_140_s_0_420=6.79e-11 mcm1p1_cf_w_0_140_s_0_420=1.34e-11
+  mcm1p1_ca_w_0_140_s_0_560=7.32e-05 mcm1p1_cc_w_0_140_s_0_560=5.17e-11 mcm1p1_cf_w_0_140_s_0_560=1.74e-11
+  mcm1p1_ca_w_0_140_s_0_840=7.32e-05 mcm1p1_cc_w_0_140_s_0_840=3.46e-11 mcm1p1_cf_w_0_140_s_0_840=2.43e-11
+  mcm1p1_ca_w_0_140_s_1_540=7.32e-05 mcm1p1_cc_w_0_140_s_1_540=1.73e-11 mcm1p1_cf_w_0_140_s_1_540=3.57e-11
+  mcm1p1_ca_w_0_140_s_3_500=7.32e-05 mcm1p1_cc_w_0_140_s_3_500=5.25e-12 mcm1p1_cf_w_0_140_s_3_500=4.67e-11
+  mcm1p1_ca_w_1_120_s_0_140=7.32e-05 mcm1p1_cc_w_1_120_s_0_140=1.46e-10 mcm1p1_cf_w_1_120_s_0_140=4.17e-12
+  mcm1p1_ca_w_1_120_s_0_175=7.32e-05 mcm1p1_cc_w_1_120_s_0_175=1.38e-10 mcm1p1_cf_w_1_120_s_0_175=5.42e-12
+  mcm1p1_ca_w_1_120_s_0_210=7.32e-05 mcm1p1_cc_w_1_120_s_0_210=1.30e-10 mcm1p1_cf_w_1_120_s_0_210=6.66e-12
+  mcm1p1_ca_w_1_120_s_0_280=7.32e-05 mcm1p1_cc_w_1_120_s_0_280=1.10e-10 mcm1p1_cf_w_1_120_s_0_280=9.06e-12
+  mcm1p1_ca_w_1_120_s_0_350=7.32e-05 mcm1p1_cc_w_1_120_s_0_350=9.38e-11 mcm1p1_cf_w_1_120_s_0_350=1.14e-11
+  mcm1p1_ca_w_1_120_s_0_420=7.32e-05 mcm1p1_cc_w_1_120_s_0_420=8.11e-11 mcm1p1_cf_w_1_120_s_0_420=1.36e-11
+  mcm1p1_ca_w_1_120_s_0_560=7.32e-05 mcm1p1_cc_w_1_120_s_0_560=6.31e-11 mcm1p1_cf_w_1_120_s_0_560=1.77e-11
+  mcm1p1_ca_w_1_120_s_0_840=7.32e-05 mcm1p1_cc_w_1_120_s_0_840=4.41e-11 mcm1p1_cf_w_1_120_s_0_840=2.47e-11
+  mcm1p1_ca_w_1_120_s_1_540=7.32e-05 mcm1p1_cc_w_1_120_s_1_540=2.44e-11 mcm1p1_cf_w_1_120_s_1_540=3.65e-11
+  mcm1p1_ca_w_1_120_s_3_500=7.32e-05 mcm1p1_cc_w_1_120_s_3_500=9.10e-12 mcm1p1_cf_w_1_120_s_3_500=4.98e-11
+  mcm1l1_ca_w_0_140_s_0_140=2.15e-04 mcm1l1_cc_w_0_140_s_0_140=1.16e-10 mcm1l1_cf_w_0_140_s_0_140=1.06e-11
+  mcm1l1_ca_w_0_140_s_0_175=2.15e-04 mcm1l1_cc_w_0_140_s_0_175=1.09e-10 mcm1l1_cf_w_0_140_s_0_175=1.43e-11
+  mcm1l1_ca_w_0_140_s_0_210=2.15e-04 mcm1l1_cc_w_0_140_s_0_210=1.01e-10 mcm1l1_cf_w_0_140_s_0_210=1.78e-11
+  mcm1l1_ca_w_0_140_s_0_280=2.15e-04 mcm1l1_cc_w_0_140_s_0_280=8.36e-11 mcm1l1_cf_w_0_140_s_0_280=2.41e-11
+  mcm1l1_ca_w_0_140_s_0_350=2.15e-04 mcm1l1_cc_w_0_140_s_0_350=6.87e-11 mcm1l1_cf_w_0_140_s_0_350=2.96e-11
+  mcm1l1_ca_w_0_140_s_0_420=2.15e-04 mcm1l1_cc_w_0_140_s_0_420=5.68e-11 mcm1l1_cf_w_0_140_s_0_420=3.45e-11
+  mcm1l1_ca_w_0_140_s_0_560=2.15e-04 mcm1l1_cc_w_0_140_s_0_560=4.14e-11 mcm1l1_cf_w_0_140_s_0_560=4.23e-11
+  mcm1l1_ca_w_0_140_s_0_840=2.15e-04 mcm1l1_cc_w_0_140_s_0_840=2.55e-11 mcm1l1_cf_w_0_140_s_0_840=5.30e-11
+  mcm1l1_ca_w_0_140_s_1_540=2.15e-04 mcm1l1_cc_w_0_140_s_1_540=1.11e-11 mcm1l1_cf_w_0_140_s_1_540=6.59e-11
+  mcm1l1_ca_w_0_140_s_3_500=2.15e-04 mcm1l1_cc_w_0_140_s_3_500=3.05e-12 mcm1l1_cf_w_0_140_s_3_500=7.42e-11
+  mcm1l1_ca_w_1_120_s_0_140=2.15e-04 mcm1l1_cc_w_1_120_s_0_140=1.33e-10 mcm1l1_cf_w_1_120_s_0_140=1.08e-11
+  mcm1l1_ca_w_1_120_s_0_175=2.15e-04 mcm1l1_cc_w_1_120_s_0_175=1.25e-10 mcm1l1_cf_w_1_120_s_0_175=1.45e-11
+  mcm1l1_ca_w_1_120_s_0_210=2.15e-04 mcm1l1_cc_w_1_120_s_0_210=1.17e-10 mcm1l1_cf_w_1_120_s_0_210=1.80e-11
+  mcm1l1_ca_w_1_120_s_0_280=2.15e-04 mcm1l1_cc_w_1_120_s_0_280=9.73e-11 mcm1l1_cf_w_1_120_s_0_280=2.43e-11
+  mcm1l1_ca_w_1_120_s_0_350=2.15e-04 mcm1l1_cc_w_1_120_s_0_350=8.19e-11 mcm1l1_cf_w_1_120_s_0_350=2.98e-11
+  mcm1l1_ca_w_1_120_s_0_420=2.15e-04 mcm1l1_cc_w_1_120_s_0_420=6.93e-11 mcm1l1_cf_w_1_120_s_0_420=3.47e-11
+  mcm1l1_ca_w_1_120_s_0_560=2.15e-04 mcm1l1_cc_w_1_120_s_0_560=5.23e-11 mcm1l1_cf_w_1_120_s_0_560=4.25e-11
+  mcm1l1_ca_w_1_120_s_0_840=2.15e-04 mcm1l1_cc_w_1_120_s_0_840=3.48e-11 mcm1l1_cf_w_1_120_s_0_840=5.33e-11
+  mcm1l1_ca_w_1_120_s_1_540=2.15e-04 mcm1l1_cc_w_1_120_s_1_540=1.81e-11 mcm1l1_cf_w_1_120_s_1_540=6.72e-11
+  mcm1l1_ca_w_1_120_s_3_500=2.15e-04 mcm1l1_cc_w_1_120_s_3_500=6.30e-12 mcm1l1_cf_w_1_120_s_3_500=7.91e-11
+  mcm2f_ca_w_0_140_s_0_140=2.35e-05 mcm2f_cc_w_0_140_s_0_140=1.32e-10 mcm2f_cf_w_0_140_s_0_140=1.28e-12
+  mcm2f_ca_w_0_140_s_0_175=2.35e-05 mcm2f_cc_w_0_140_s_0_175=1.25e-10 mcm2f_cf_w_0_140_s_0_175=1.69e-12
+  mcm2f_ca_w_0_140_s_0_210=2.35e-05 mcm2f_cc_w_0_140_s_0_210=1.18e-10 mcm2f_cf_w_0_140_s_0_210=2.10e-12
+  mcm2f_ca_w_0_140_s_0_280=2.35e-05 mcm2f_cc_w_0_140_s_0_280=1.01e-10 mcm2f_cf_w_0_140_s_0_280=2.91e-12
+  mcm2f_ca_w_0_140_s_0_350=2.35e-05 mcm2f_cc_w_0_140_s_0_350=8.71e-11 mcm2f_cf_w_0_140_s_0_350=3.70e-12
+  mcm2f_ca_w_0_140_s_0_420=2.35e-05 mcm2f_cc_w_0_140_s_0_420=7.61e-11 mcm2f_cf_w_0_140_s_0_420=4.52e-12
+  mcm2f_ca_w_0_140_s_0_560=2.35e-05 mcm2f_cc_w_0_140_s_0_560=6.02e-11 mcm2f_cf_w_0_140_s_0_560=6.00e-12
+  mcm2f_ca_w_0_140_s_0_840=2.35e-05 mcm2f_cc_w_0_140_s_0_840=4.41e-11 mcm2f_cf_w_0_140_s_0_840=8.90e-12
+  mcm2f_ca_w_0_140_s_1_540=2.35e-05 mcm2f_cc_w_0_140_s_1_540=2.69e-11 mcm2f_cf_w_0_140_s_1_540=1.51e-11
+  mcm2f_ca_w_0_140_s_3_500=2.35e-05 mcm2f_cc_w_0_140_s_3_500=1.14e-11 mcm2f_cf_w_0_140_s_3_500=2.56e-11
+  mcm2f_ca_w_1_120_s_0_140=2.35e-05 mcm2f_cc_w_1_120_s_0_140=1.57e-10 mcm2f_cf_w_1_120_s_0_140=1.32e-12
+  mcm2f_ca_w_1_120_s_0_175=2.35e-05 mcm2f_cc_w_1_120_s_0_175=1.49e-10 mcm2f_cf_w_1_120_s_0_175=1.73e-12
+  mcm2f_ca_w_1_120_s_0_210=2.35e-05 mcm2f_cc_w_1_120_s_0_210=1.41e-10 mcm2f_cf_w_1_120_s_0_210=2.14e-12
+  mcm2f_ca_w_1_120_s_0_280=2.35e-05 mcm2f_cc_w_1_120_s_0_280=1.21e-10 mcm2f_cf_w_1_120_s_0_280=2.95e-12
+  mcm2f_ca_w_1_120_s_0_350=2.35e-05 mcm2f_cc_w_1_120_s_0_350=1.05e-10 mcm2f_cf_w_1_120_s_0_350=3.74e-12
+  mcm2f_ca_w_1_120_s_0_420=2.35e-05 mcm2f_cc_w_1_120_s_0_420=9.25e-11 mcm2f_cf_w_1_120_s_0_420=4.54e-12
+  mcm2f_ca_w_1_120_s_0_560=2.35e-05 mcm2f_cc_w_1_120_s_0_560=7.44e-11 mcm2f_cf_w_1_120_s_0_560=6.06e-12
+  mcm2f_ca_w_1_120_s_0_840=2.35e-05 mcm2f_cc_w_1_120_s_0_840=5.54e-11 mcm2f_cf_w_1_120_s_0_840=9.00e-12
+  mcm2f_ca_w_1_120_s_1_540=2.35e-05 mcm2f_cc_w_1_120_s_1_540=3.50e-11 mcm2f_cf_w_1_120_s_1_540=1.54e-11
+  mcm2f_ca_w_1_120_s_3_500=2.35e-05 mcm2f_cc_w_1_120_s_3_500=1.61e-11 mcm2f_cf_w_1_120_s_3_500=2.71e-11
+  mcm2d_ca_w_0_140_s_0_140=2.74e-05 mcm2d_cc_w_0_140_s_0_140=1.31e-10 mcm2d_cf_w_0_140_s_0_140=1.49e-12
+  mcm2d_ca_w_0_140_s_0_175=2.74e-05 mcm2d_cc_w_0_140_s_0_175=1.24e-10 mcm2d_cf_w_0_140_s_0_175=1.97e-12
+  mcm2d_ca_w_0_140_s_0_210=2.74e-05 mcm2d_cc_w_0_140_s_0_210=1.18e-10 mcm2d_cf_w_0_140_s_0_210=2.45e-12
+  mcm2d_ca_w_0_140_s_0_280=2.74e-05 mcm2d_cc_w_0_140_s_0_280=1.01e-10 mcm2d_cf_w_0_140_s_0_280=3.39e-12
+  mcm2d_ca_w_0_140_s_0_350=2.74e-05 mcm2d_cc_w_0_140_s_0_350=8.64e-11 mcm2d_cf_w_0_140_s_0_350=4.31e-12
+  mcm2d_ca_w_0_140_s_0_420=2.74e-05 mcm2d_cc_w_0_140_s_0_420=7.51e-11 mcm2d_cf_w_0_140_s_0_420=5.25e-12
+  mcm2d_ca_w_0_140_s_0_560=2.74e-05 mcm2d_cc_w_0_140_s_0_560=5.93e-11 mcm2d_cf_w_0_140_s_0_560=6.96e-12
+  mcm2d_ca_w_0_140_s_0_840=2.74e-05 mcm2d_cc_w_0_140_s_0_840=4.28e-11 mcm2d_cf_w_0_140_s_0_840=1.03e-11
+  mcm2d_ca_w_0_140_s_1_540=2.74e-05 mcm2d_cc_w_0_140_s_1_540=2.55e-11 mcm2d_cf_w_0_140_s_1_540=1.72e-11
+  mcm2d_ca_w_0_140_s_3_500=2.74e-05 mcm2d_cc_w_0_140_s_3_500=1.02e-11 mcm2d_cf_w_0_140_s_3_500=2.82e-11
+  mcm2d_ca_w_1_120_s_0_140=2.74e-05 mcm2d_cc_w_1_120_s_0_140=1.55e-10 mcm2d_cf_w_1_120_s_0_140=1.54e-12
+  mcm2d_ca_w_1_120_s_0_175=2.74e-05 mcm2d_cc_w_1_120_s_0_175=1.47e-10 mcm2d_cf_w_1_120_s_0_175=2.02e-12
+  mcm2d_ca_w_1_120_s_0_210=2.74e-05 mcm2d_cc_w_1_120_s_0_210=1.39e-10 mcm2d_cf_w_1_120_s_0_210=2.49e-12
+  mcm2d_ca_w_1_120_s_0_280=2.74e-05 mcm2d_cc_w_1_120_s_0_280=1.19e-10 mcm2d_cf_w_1_120_s_0_280=3.43e-12
+  mcm2d_ca_w_1_120_s_0_350=2.74e-05 mcm2d_cc_w_1_120_s_0_350=1.04e-10 mcm2d_cf_w_1_120_s_0_350=4.36e-12
+  mcm2d_ca_w_1_120_s_0_420=2.74e-05 mcm2d_cc_w_1_120_s_0_420=9.08e-11 mcm2d_cf_w_1_120_s_0_420=5.27e-12
+  mcm2d_ca_w_1_120_s_0_560=2.74e-05 mcm2d_cc_w_1_120_s_0_560=7.29e-11 mcm2d_cf_w_1_120_s_0_560=7.04e-12
+  mcm2d_ca_w_1_120_s_0_840=2.74e-05 mcm2d_cc_w_1_120_s_0_840=5.38e-11 mcm2d_cf_w_1_120_s_0_840=1.04e-11
+  mcm2d_ca_w_1_120_s_1_540=2.74e-05 mcm2d_cc_w_1_120_s_1_540=3.33e-11 mcm2d_cf_w_1_120_s_1_540=1.75e-11
+  mcm2d_ca_w_1_120_s_3_500=2.74e-05 mcm2d_cc_w_1_120_s_3_500=1.48e-11 mcm2d_cf_w_1_120_s_3_500=2.98e-11
+  mcm2p1_ca_w_0_140_s_0_140=3.55e-05 mcm2p1_cc_w_0_140_s_0_140=1.30e-10 mcm2p1_cf_w_0_140_s_0_140=1.94e-12
+  mcm2p1_ca_w_0_140_s_0_175=3.55e-05 mcm2p1_cc_w_0_140_s_0_175=1.23e-10 mcm2p1_cf_w_0_140_s_0_175=2.55e-12
+  mcm2p1_ca_w_0_140_s_0_210=3.55e-05 mcm2p1_cc_w_0_140_s_0_210=1.17e-10 mcm2p1_cf_w_0_140_s_0_210=3.17e-12
+  mcm2p1_ca_w_0_140_s_0_280=3.55e-05 mcm2p1_cc_w_0_140_s_0_280=9.92e-11 mcm2p1_cf_w_0_140_s_0_280=4.39e-12
+  mcm2p1_ca_w_0_140_s_0_350=3.55e-05 mcm2p1_cc_w_0_140_s_0_350=8.48e-11 mcm2p1_cf_w_0_140_s_0_350=5.57e-12
+  mcm2p1_ca_w_0_140_s_0_420=3.55e-05 mcm2p1_cc_w_0_140_s_0_420=7.32e-11 mcm2p1_cf_w_0_140_s_0_420=6.76e-12
+  mcm2p1_ca_w_0_140_s_0_560=3.55e-05 mcm2p1_cc_w_0_140_s_0_560=5.76e-11 mcm2p1_cf_w_0_140_s_0_560=8.95e-12
+  mcm2p1_ca_w_0_140_s_0_840=3.55e-05 mcm2p1_cc_w_0_140_s_0_840=4.08e-11 mcm2p1_cf_w_0_140_s_0_840=1.30e-11
+  mcm2p1_ca_w_0_140_s_1_540=3.55e-05 mcm2p1_cc_w_0_140_s_1_540=2.31e-11 mcm2p1_cf_w_0_140_s_1_540=2.12e-11
+  mcm2p1_ca_w_0_140_s_3_500=3.55e-05 mcm2p1_cc_w_0_140_s_3_500=8.47e-12 mcm2p1_cf_w_0_140_s_3_500=3.27e-11
+  mcm2p1_ca_w_1_120_s_0_140=3.55e-05 mcm2p1_cc_w_1_120_s_0_140=1.53e-10 mcm2p1_cf_w_1_120_s_0_140=2.02e-12
+  mcm2p1_ca_w_1_120_s_0_175=3.55e-05 mcm2p1_cc_w_1_120_s_0_175=1.44e-10 mcm2p1_cf_w_1_120_s_0_175=2.64e-12
+  mcm2p1_ca_w_1_120_s_0_210=3.55e-05 mcm2p1_cc_w_1_120_s_0_210=1.36e-10 mcm2p1_cf_w_1_120_s_0_210=3.26e-12
+  mcm2p1_ca_w_1_120_s_0_280=3.55e-05 mcm2p1_cc_w_1_120_s_0_280=1.17e-10 mcm2p1_cf_w_1_120_s_0_280=4.47e-12
+  mcm2p1_ca_w_1_120_s_0_350=3.55e-05 mcm2p1_cc_w_1_120_s_0_350=1.01e-10 mcm2p1_cf_w_1_120_s_0_350=5.66e-12
+  mcm2p1_ca_w_1_120_s_0_420=3.55e-05 mcm2p1_cc_w_1_120_s_0_420=8.78e-11 mcm2p1_cf_w_1_120_s_0_420=6.83e-12
+  mcm2p1_ca_w_1_120_s_0_560=3.55e-05 mcm2p1_cc_w_1_120_s_0_560=7.01e-11 mcm2p1_cf_w_1_120_s_0_560=9.04e-12
+  mcm2p1_ca_w_1_120_s_0_840=3.55e-05 mcm2p1_cc_w_1_120_s_0_840=5.08e-11 mcm2p1_cf_w_1_120_s_0_840=1.32e-11
+  mcm2p1_ca_w_1_120_s_1_540=3.55e-05 mcm2p1_cc_w_1_120_s_1_540=3.06e-11 mcm2p1_cf_w_1_120_s_1_540=2.16e-11
+  mcm2p1_ca_w_1_120_s_3_500=3.55e-05 mcm2p1_cc_w_1_120_s_3_500=1.28e-11 mcm2p1_cf_w_1_120_s_3_500=3.46e-11
+  mcm2l1_ca_w_0_140_s_0_140=5.23e-05 mcm2l1_cc_w_0_140_s_0_140=1.28e-10 mcm2l1_cf_w_0_140_s_0_140=2.79e-12
+  mcm2l1_ca_w_0_140_s_0_175=5.23e-05 mcm2l1_cc_w_0_140_s_0_175=1.21e-10 mcm2l1_cf_w_0_140_s_0_175=3.70e-12
+  mcm2l1_ca_w_0_140_s_0_210=5.23e-05 mcm2l1_cc_w_0_140_s_0_210=1.14e-10 mcm2l1_cf_w_0_140_s_0_210=4.60e-12
+  mcm2l1_ca_w_0_140_s_0_280=5.23e-05 mcm2l1_cc_w_0_140_s_0_280=9.69e-11 mcm2l1_cf_w_0_140_s_0_280=6.36e-12
+  mcm2l1_ca_w_0_140_s_0_350=5.23e-05 mcm2l1_cc_w_0_140_s_0_350=8.22e-11 mcm2l1_cf_w_0_140_s_0_350=8.06e-12
+  mcm2l1_ca_w_0_140_s_0_420=5.23e-05 mcm2l1_cc_w_0_140_s_0_420=7.06e-11 mcm2l1_cf_w_0_140_s_0_420=9.73e-12
+  mcm2l1_ca_w_0_140_s_0_560=5.23e-05 mcm2l1_cc_w_0_140_s_0_560=5.42e-11 mcm2l1_cf_w_0_140_s_0_560=1.28e-11
+  mcm2l1_ca_w_0_140_s_0_840=5.23e-05 mcm2l1_cc_w_0_140_s_0_840=3.72e-11 mcm2l1_cf_w_0_140_s_0_840=1.83e-11
+  mcm2l1_ca_w_0_140_s_1_540=5.23e-05 mcm2l1_cc_w_0_140_s_1_540=1.97e-11 mcm2l1_cf_w_0_140_s_1_540=2.82e-11
+  mcm2l1_ca_w_0_140_s_3_500=5.23e-05 mcm2l1_cc_w_0_140_s_3_500=6.44e-12 mcm2l1_cf_w_0_140_s_3_500=3.95e-11
+  mcm2l1_ca_w_1_120_s_0_140=5.23e-05 mcm2l1_cc_w_1_120_s_0_140=1.48e-10 mcm2l1_cf_w_1_120_s_0_140=2.83e-12
+  mcm2l1_ca_w_1_120_s_0_175=5.23e-05 mcm2l1_cc_w_1_120_s_0_175=1.40e-10 mcm2l1_cf_w_1_120_s_0_175=3.75e-12
+  mcm2l1_ca_w_1_120_s_0_210=5.23e-05 mcm2l1_cc_w_1_120_s_0_210=1.32e-10 mcm2l1_cf_w_1_120_s_0_210=4.65e-12
+  mcm2l1_ca_w_1_120_s_0_280=5.23e-05 mcm2l1_cc_w_1_120_s_0_280=1.13e-10 mcm2l1_cf_w_1_120_s_0_280=6.40e-12
+  mcm2l1_ca_w_1_120_s_0_350=5.23e-05 mcm2l1_cc_w_1_120_s_0_350=9.66e-11 mcm2l1_cf_w_1_120_s_0_350=8.10e-12
+  mcm2l1_ca_w_1_120_s_0_420=5.23e-05 mcm2l1_cc_w_1_120_s_0_420=8.37e-11 mcm2l1_cf_w_1_120_s_0_420=9.75e-12
+  mcm2l1_ca_w_1_120_s_0_560=5.23e-05 mcm2l1_cc_w_1_120_s_0_560=6.59e-11 mcm2l1_cf_w_1_120_s_0_560=1.29e-11
+  mcm2l1_ca_w_1_120_s_0_840=5.23e-05 mcm2l1_cc_w_1_120_s_0_840=4.68e-11 mcm2l1_cf_w_1_120_s_0_840=1.84e-11
+  mcm2l1_ca_w_1_120_s_1_540=5.23e-05 mcm2l1_cc_w_1_120_s_1_540=2.69e-11 mcm2l1_cf_w_1_120_s_1_540=2.87e-11
+  mcm2l1_ca_w_1_120_s_3_500=5.23e-05 mcm2l1_cc_w_1_120_s_3_500=1.05e-11 mcm2l1_cf_w_1_120_s_3_500=4.20e-11
+  mcm2m1_ca_w_0_140_s_0_140=3.13e-04 mcm2m1_cc_w_0_140_s_0_140=1.12e-10 mcm2m1_cf_w_0_140_s_0_140=1.45e-11
+  mcm2m1_ca_w_0_140_s_0_175=3.13e-04 mcm2m1_cc_w_0_140_s_0_175=1.05e-10 mcm2m1_cf_w_0_140_s_0_175=1.99e-11
+  mcm2m1_ca_w_0_140_s_0_210=3.13e-04 mcm2m1_cc_w_0_140_s_0_210=9.67e-11 mcm2m1_cf_w_0_140_s_0_210=2.47e-11
+  mcm2m1_ca_w_0_140_s_0_280=3.13e-04 mcm2m1_cc_w_0_140_s_0_280=7.97e-11 mcm2m1_cf_w_0_140_s_0_280=3.33e-11
+  mcm2m1_ca_w_0_140_s_0_350=3.13e-04 mcm2m1_cc_w_0_140_s_0_350=6.51e-11 mcm2m1_cf_w_0_140_s_0_350=4.03e-11
+  mcm2m1_ca_w_0_140_s_0_420=3.13e-04 mcm2m1_cc_w_0_140_s_0_420=5.34e-11 mcm2m1_cf_w_0_140_s_0_420=4.63e-11
+  mcm2m1_ca_w_0_140_s_0_560=3.13e-04 mcm2m1_cc_w_0_140_s_0_560=3.83e-11 mcm2m1_cf_w_0_140_s_0_560=5.53e-11
+  mcm2m1_ca_w_0_140_s_0_840=3.13e-04 mcm2m1_cc_w_0_140_s_0_840=2.34e-11 mcm2m1_cf_w_0_140_s_0_840=6.69e-11
+  mcm2m1_ca_w_0_140_s_1_540=3.13e-04 mcm2m1_cc_w_0_140_s_1_540=1.00e-11 mcm2m1_cf_w_0_140_s_1_540=7.99e-11
+  mcm2m1_ca_w_0_140_s_3_500=3.13e-04 mcm2m1_cc_w_0_140_s_3_500=2.75e-12 mcm2m1_cf_w_0_140_s_3_500=8.84e-11
+  mcm2m1_ca_w_1_120_s_0_140=3.13e-04 mcm2m1_cc_w_1_120_s_0_140=1.29e-10 mcm2m1_cf_w_1_120_s_0_140=1.45e-11
+  mcm2m1_ca_w_1_120_s_0_175=3.13e-04 mcm2m1_cc_w_1_120_s_0_175=1.21e-10 mcm2m1_cf_w_1_120_s_0_175=1.99e-11
+  mcm2m1_ca_w_1_120_s_0_210=3.13e-04 mcm2m1_cc_w_1_120_s_0_210=1.12e-10 mcm2m1_cf_w_1_120_s_0_210=2.47e-11
+  mcm2m1_ca_w_1_120_s_0_280=3.13e-04 mcm2m1_cc_w_1_120_s_0_280=9.35e-11 mcm2m1_cf_w_1_120_s_0_280=3.32e-11
+  mcm2m1_ca_w_1_120_s_0_350=3.13e-04 mcm2m1_cc_w_1_120_s_0_350=7.84e-11 mcm2m1_cf_w_1_120_s_0_350=4.03e-11
+  mcm2m1_ca_w_1_120_s_0_420=3.13e-04 mcm2m1_cc_w_1_120_s_0_420=6.60e-11 mcm2m1_cf_w_1_120_s_0_420=4.61e-11
+  mcm2m1_ca_w_1_120_s_0_560=3.13e-04 mcm2m1_cc_w_1_120_s_0_560=4.95e-11 mcm2m1_cf_w_1_120_s_0_560=5.53e-11
+  mcm2m1_ca_w_1_120_s_0_840=3.13e-04 mcm2m1_cc_w_1_120_s_0_840=3.28e-11 mcm2m1_cf_w_1_120_s_0_840=6.71e-11
+  mcm2m1_ca_w_1_120_s_1_540=3.13e-04 mcm2m1_cc_w_1_120_s_1_540=1.70e-11 mcm2m1_cf_w_1_120_s_1_540=8.15e-11
+  mcm2m1_ca_w_1_120_s_3_500=3.13e-04 mcm2m1_cc_w_1_120_s_3_500=5.90e-12 mcm2m1_cf_w_1_120_s_3_500=9.31e-11
+  mcm3f_ca_w_0_300_s_0_300=1.63e-05 mcm3f_cc_w_0_300_s_0_300=1.24e-10 mcm3f_cf_w_0_300_s_0_300=2.03e-12
+  mcm3f_ca_w_0_300_s_0_360=1.63e-05 mcm3f_cc_w_0_300_s_0_360=1.14e-10 mcm3f_cf_w_0_300_s_0_360=2.50e-12
+  mcm3f_ca_w_0_300_s_0_450=1.63e-05 mcm3f_cc_w_0_300_s_0_450=1.02e-10 mcm3f_cf_w_0_300_s_0_450=3.22e-12
+  mcm3f_ca_w_0_300_s_0_600=1.63e-05 mcm3f_cc_w_0_300_s_0_600=8.58e-11 mcm3f_cf_w_0_300_s_0_600=4.38e-12
+  mcm3f_ca_w_0_300_s_0_800=1.63e-05 mcm3f_cc_w_0_300_s_0_800=7.13e-11 mcm3f_cf_w_0_300_s_0_800=5.81e-12
+  mcm3f_ca_w_0_300_s_1_000=1.63e-05 mcm3f_cc_w_0_300_s_1_000=6.06e-11 mcm3f_cf_w_0_300_s_1_000=7.23e-12
+  mcm3f_ca_w_0_300_s_1_200=1.63e-05 mcm3f_cc_w_0_300_s_1_200=5.25e-11 mcm3f_cf_w_0_300_s_1_200=8.58e-12
+  mcm3f_ca_w_0_300_s_2_100=1.63e-05 mcm3f_cc_w_0_300_s_2_100=3.33e-11 mcm3f_cf_w_0_300_s_2_100=1.43e-11
+  mcm3f_ca_w_0_300_s_3_300=1.63e-05 mcm3f_cc_w_0_300_s_3_300=2.24e-11 mcm3f_cf_w_0_300_s_3_300=1.99e-11
+  mcm3f_ca_w_0_300_s_9_000=1.63e-05 mcm3f_cc_w_0_300_s_9_000=6.33e-12 mcm3f_cf_w_0_300_s_9_000=3.26e-11
+  mcm3f_ca_w_2_400_s_0_300=1.63e-05 mcm3f_cc_w_2_400_s_0_300=1.48e-10 mcm3f_cf_w_2_400_s_0_300=2.08e-12
+  mcm3f_ca_w_2_400_s_0_360=1.63e-05 mcm3f_cc_w_2_400_s_0_360=1.37e-10 mcm3f_cf_w_2_400_s_0_360=2.55e-12
+  mcm3f_ca_w_2_400_s_0_450=1.63e-05 mcm3f_cc_w_2_400_s_0_450=1.23e-10 mcm3f_cf_w_2_400_s_0_450=3.25e-12
+  mcm3f_ca_w_2_400_s_0_600=1.63e-05 mcm3f_cc_w_2_400_s_0_600=1.05e-10 mcm3f_cf_w_2_400_s_0_600=4.40e-12
+  mcm3f_ca_w_2_400_s_0_800=1.63e-05 mcm3f_cc_w_2_400_s_0_800=8.77e-11 mcm3f_cf_w_2_400_s_0_800=5.88e-12
+  mcm3f_ca_w_2_400_s_1_000=1.63e-05 mcm3f_cc_w_2_400_s_1_000=7.53e-11 mcm3f_cf_w_2_400_s_1_000=7.34e-12
+  mcm3f_ca_w_2_400_s_1_200=1.63e-05 mcm3f_cc_w_2_400_s_1_200=6.62e-11 mcm3f_cf_w_2_400_s_1_200=8.72e-12
+  mcm3f_ca_w_2_400_s_2_100=1.63e-05 mcm3f_cc_w_2_400_s_2_100=4.39e-11 mcm3f_cf_w_2_400_s_2_100=1.44e-11
+  mcm3f_ca_w_2_400_s_3_300=1.63e-05 mcm3f_cc_w_2_400_s_3_300=3.04e-11 mcm3f_cf_w_2_400_s_3_300=2.05e-11
+  mcm3f_ca_w_2_400_s_9_000=1.63e-05 mcm3f_cc_w_2_400_s_9_000=1.01e-11 mcm3f_cf_w_2_400_s_9_000=3.54e-11
+  mcm3d_ca_w_0_300_s_0_300=1.81e-05 mcm3d_cc_w_0_300_s_0_300=1.23e-10 mcm3d_cf_w_0_300_s_0_300=2.24e-12
+  mcm3d_ca_w_0_300_s_0_360=1.81e-05 mcm3d_cc_w_0_300_s_0_360=1.14e-10 mcm3d_cf_w_0_300_s_0_360=2.76e-12
+  mcm3d_ca_w_0_300_s_0_450=1.81e-05 mcm3d_cc_w_0_300_s_0_450=1.01e-10 mcm3d_cf_w_0_300_s_0_450=3.56e-12
+  mcm3d_ca_w_0_300_s_0_600=1.81e-05 mcm3d_cc_w_0_300_s_0_600=8.53e-11 mcm3d_cf_w_0_300_s_0_600=4.83e-12
+  mcm3d_ca_w_0_300_s_0_800=1.81e-05 mcm3d_cc_w_0_300_s_0_800=7.06e-11 mcm3d_cf_w_0_300_s_0_800=6.40e-12
+  mcm3d_ca_w_0_300_s_1_000=1.81e-05 mcm3d_cc_w_0_300_s_1_000=5.98e-11 mcm3d_cf_w_0_300_s_1_000=7.96e-12
+  mcm3d_ca_w_0_300_s_1_200=1.81e-05 mcm3d_cc_w_0_300_s_1_200=5.17e-11 mcm3d_cf_w_0_300_s_1_200=9.43e-12
+  mcm3d_ca_w_0_300_s_2_100=1.81e-05 mcm3d_cc_w_0_300_s_2_100=3.24e-11 mcm3d_cf_w_0_300_s_2_100=1.56e-11
+  mcm3d_ca_w_0_300_s_3_300=1.81e-05 mcm3d_cc_w_0_300_s_3_300=2.15e-11 mcm3d_cf_w_0_300_s_3_300=2.15e-11
+  mcm3d_ca_w_0_300_s_9_000=1.81e-05 mcm3d_cc_w_0_300_s_9_000=5.90e-12 mcm3d_cf_w_0_300_s_9_000=3.41e-11
+  mcm3d_ca_w_2_400_s_0_300=1.81e-05 mcm3d_cc_w_2_400_s_0_300=1.46e-10 mcm3d_cf_w_2_400_s_0_300=2.31e-12
+  mcm3d_ca_w_2_400_s_0_360=1.81e-05 mcm3d_cc_w_2_400_s_0_360=1.36e-10 mcm3d_cf_w_2_400_s_0_360=2.83e-12
+  mcm3d_ca_w_2_400_s_0_450=1.81e-05 mcm3d_cc_w_2_400_s_0_450=1.22e-10 mcm3d_cf_w_2_400_s_0_450=3.60e-12
+  mcm3d_ca_w_2_400_s_0_600=1.81e-05 mcm3d_cc_w_2_400_s_0_600=1.04e-10 mcm3d_cf_w_2_400_s_0_600=4.87e-12
+  mcm3d_ca_w_2_400_s_0_800=1.81e-05 mcm3d_cc_w_2_400_s_0_800=8.66e-11 mcm3d_cf_w_2_400_s_0_800=6.49e-12
+  mcm3d_ca_w_2_400_s_1_000=1.81e-05 mcm3d_cc_w_2_400_s_1_000=7.42e-11 mcm3d_cf_w_2_400_s_1_000=8.08e-12
+  mcm3d_ca_w_2_400_s_1_200=1.81e-05 mcm3d_cc_w_2_400_s_1_200=6.50e-11 mcm3d_cf_w_2_400_s_1_200=9.58e-12
+  mcm3d_ca_w_2_400_s_2_100=1.81e-05 mcm3d_cc_w_2_400_s_2_100=4.28e-11 mcm3d_cf_w_2_400_s_2_100=1.56e-11
+  mcm3d_ca_w_2_400_s_3_300=1.81e-05 mcm3d_cc_w_2_400_s_3_300=2.94e-11 mcm3d_cf_w_2_400_s_3_300=2.21e-11
+  mcm3d_ca_w_2_400_s_9_000=1.81e-05 mcm3d_cc_w_2_400_s_9_000=9.50e-12 mcm3d_cf_w_2_400_s_9_000=3.72e-11
+  mcm3p1_ca_w_0_300_s_0_300=2.13e-05 mcm3p1_cc_w_0_300_s_0_300=1.23e-10 mcm3p1_cf_w_0_300_s_0_300=2.64e-12
+  mcm3p1_ca_w_0_300_s_0_360=2.13e-05 mcm3p1_cc_w_0_300_s_0_360=1.13e-10 mcm3p1_cf_w_0_300_s_0_360=3.25e-12
+  mcm3p1_ca_w_0_300_s_0_450=2.13e-05 mcm3p1_cc_w_0_300_s_0_450=1.00e-10 mcm3p1_cf_w_0_300_s_0_450=4.17e-12
+  mcm3p1_ca_w_0_300_s_0_600=2.13e-05 mcm3p1_cc_w_0_300_s_0_600=8.43e-11 mcm3p1_cf_w_0_300_s_0_600=5.64e-12
+  mcm3p1_ca_w_0_300_s_0_800=2.13e-05 mcm3p1_cc_w_0_300_s_0_800=6.93e-11 mcm3p1_cf_w_0_300_s_0_800=7.46e-12
+  mcm3p1_ca_w_0_300_s_1_000=2.13e-05 mcm3p1_cc_w_0_300_s_1_000=5.86e-11 mcm3p1_cf_w_0_300_s_1_000=9.26e-12
+  mcm3p1_ca_w_0_300_s_1_200=2.13e-05 mcm3p1_cc_w_0_300_s_1_200=5.04e-11 mcm3p1_cf_w_0_300_s_1_200=1.09e-11
+  mcm3p1_ca_w_0_300_s_2_100=2.13e-05 mcm3p1_cc_w_0_300_s_2_100=3.10e-11 mcm3p1_cf_w_0_300_s_2_100=1.79e-11
+  mcm3p1_ca_w_0_300_s_3_300=2.13e-05 mcm3p1_cc_w_0_300_s_3_300=2.01e-11 mcm3p1_cf_w_0_300_s_3_300=2.41e-11
+  mcm3p1_ca_w_0_300_s_9_000=2.13e-05 mcm3p1_cc_w_0_300_s_9_000=5.22e-12 mcm3p1_cf_w_0_300_s_9_000=3.65e-11
+  mcm3p1_ca_w_2_400_s_0_300=2.13e-05 mcm3p1_cc_w_2_400_s_0_300=1.45e-10 mcm3p1_cf_w_2_400_s_0_300=2.74e-12
+  mcm3p1_ca_w_2_400_s_0_360=2.13e-05 mcm3p1_cc_w_2_400_s_0_360=1.34e-10 mcm3p1_cf_w_2_400_s_0_360=3.33e-12
+  mcm3p1_ca_w_2_400_s_0_450=2.13e-05 mcm3p1_cc_w_2_400_s_0_450=1.20e-10 mcm3p1_cf_w_2_400_s_0_450=4.23e-12
+  mcm3p1_ca_w_2_400_s_0_600=2.13e-05 mcm3p1_cc_w_2_400_s_0_600=1.02e-10 mcm3p1_cf_w_2_400_s_0_600=5.70e-12
+  mcm3p1_ca_w_2_400_s_0_800=2.13e-05 mcm3p1_cc_w_2_400_s_0_800=8.48e-11 mcm3p1_cf_w_2_400_s_0_800=7.58e-12
+  mcm3p1_ca_w_2_400_s_1_000=2.13e-05 mcm3p1_cc_w_2_400_s_1_000=7.24e-11 mcm3p1_cf_w_2_400_s_1_000=9.42e-12
+  mcm3p1_ca_w_2_400_s_1_200=2.13e-05 mcm3p1_cc_w_2_400_s_1_200=6.32e-11 mcm3p1_cf_w_2_400_s_1_200=1.11e-11
+  mcm3p1_ca_w_2_400_s_2_100=2.13e-05 mcm3p1_cc_w_2_400_s_2_100=4.11e-11 mcm3p1_cf_w_2_400_s_2_100=1.79e-11
+  mcm3p1_ca_w_2_400_s_3_300=2.13e-05 mcm3p1_cc_w_2_400_s_3_300=2.78e-11 mcm3p1_cf_w_2_400_s_3_300=2.48e-11
+  mcm3p1_ca_w_2_400_s_9_000=2.13e-05 mcm3p1_cc_w_2_400_s_9_000=8.65e-12 mcm3p1_cf_w_2_400_s_9_000=3.99e-11
+  mcm3l1_ca_w_0_300_s_0_300=2.63e-05 mcm3l1_cc_w_0_300_s_0_300=1.22e-10 mcm3l1_cf_w_0_300_s_0_300=3.23e-12
+  mcm3l1_ca_w_0_300_s_0_360=2.63e-05 mcm3l1_cc_w_0_300_s_0_360=1.11e-10 mcm3l1_cf_w_0_300_s_0_360=3.97e-12
+  mcm3l1_ca_w_0_300_s_0_450=2.63e-05 mcm3l1_cc_w_0_300_s_0_450=9.88e-11 mcm3l1_cf_w_0_300_s_0_450=5.08e-12
+  mcm3l1_ca_w_0_300_s_0_600=2.63e-05 mcm3l1_cc_w_0_300_s_0_600=8.28e-11 mcm3l1_cf_w_0_300_s_0_600=6.85e-12
+  mcm3l1_ca_w_0_300_s_0_800=2.63e-05 mcm3l1_cc_w_0_300_s_0_800=6.77e-11 mcm3l1_cf_w_0_300_s_0_800=9.04e-12
+  mcm3l1_ca_w_0_300_s_1_000=2.63e-05 mcm3l1_cc_w_0_300_s_1_000=5.68e-11 mcm3l1_cf_w_0_300_s_1_000=1.12e-11
+  mcm3l1_ca_w_0_300_s_1_200=2.63e-05 mcm3l1_cc_w_0_300_s_1_200=4.88e-11 mcm3l1_cf_w_0_300_s_1_200=1.31e-11
+  mcm3l1_ca_w_0_300_s_2_100=2.63e-05 mcm3l1_cc_w_0_300_s_2_100=2.91e-11 mcm3l1_cf_w_0_300_s_2_100=2.10e-11
+  mcm3l1_ca_w_0_300_s_3_300=2.63e-05 mcm3l1_cc_w_0_300_s_3_300=1.84e-11 mcm3l1_cf_w_0_300_s_3_300=2.77e-11
+  mcm3l1_ca_w_0_300_s_9_000=2.63e-05 mcm3l1_cc_w_0_300_s_9_000=4.48e-12 mcm3l1_cf_w_0_300_s_9_000=3.97e-11
+  mcm3l1_ca_w_2_400_s_0_300=2.63e-05 mcm3l1_cc_w_2_400_s_0_300=1.42e-10 mcm3l1_cf_w_2_400_s_0_300=3.27e-12
+  mcm3l1_ca_w_2_400_s_0_360=2.63e-05 mcm3l1_cc_w_2_400_s_0_360=1.31e-10 mcm3l1_cf_w_2_400_s_0_360=4.01e-12
+  mcm3l1_ca_w_2_400_s_0_450=2.63e-05 mcm3l1_cc_w_2_400_s_0_450=1.17e-10 mcm3l1_cf_w_2_400_s_0_450=5.11e-12
+  mcm3l1_ca_w_2_400_s_0_600=2.63e-05 mcm3l1_cc_w_2_400_s_0_600=9.97e-11 mcm3l1_cf_w_2_400_s_0_600=6.87e-12
+  mcm3l1_ca_w_2_400_s_0_800=2.63e-05 mcm3l1_cc_w_2_400_s_0_800=8.26e-11 mcm3l1_cf_w_2_400_s_0_800=9.12e-12
+  mcm3l1_ca_w_2_400_s_1_000=2.63e-05 mcm3l1_cc_w_2_400_s_1_000=7.03e-11 mcm3l1_cf_w_2_400_s_1_000=1.13e-11
+  mcm3l1_ca_w_2_400_s_1_200=2.63e-05 mcm3l1_cc_w_2_400_s_1_200=6.11e-11 mcm3l1_cf_w_2_400_s_1_200=1.33e-11
+  mcm3l1_ca_w_2_400_s_2_100=2.63e-05 mcm3l1_cc_w_2_400_s_2_100=3.91e-11 mcm3l1_cf_w_2_400_s_2_100=2.10e-11
+  mcm3l1_ca_w_2_400_s_3_300=2.63e-05 mcm3l1_cc_w_2_400_s_3_300=2.59e-11 mcm3l1_cf_w_2_400_s_3_300=2.85e-11
+  mcm3l1_ca_w_2_400_s_9_000=2.63e-05 mcm3l1_cc_w_2_400_s_9_000=7.75e-12 mcm3l1_cf_w_2_400_s_9_000=4.34e-11
+  mcm3m1_ca_w_0_300_s_0_300=4.52e-05 mcm3m1_cc_w_0_300_s_0_300=1.18e-10 mcm3m1_cf_w_0_300_s_0_300=5.43e-12
+  mcm3m1_ca_w_0_300_s_0_360=4.52e-05 mcm3m1_cc_w_0_300_s_0_360=1.07e-10 mcm3m1_cf_w_0_300_s_0_360=6.65e-12
+  mcm3m1_ca_w_0_300_s_0_450=4.52e-05 mcm3m1_cc_w_0_300_s_0_450=9.46e-11 mcm3m1_cf_w_0_300_s_0_450=8.43e-12
+  mcm3m1_ca_w_0_300_s_0_600=4.52e-05 mcm3m1_cc_w_0_300_s_0_600=7.83e-11 mcm3m1_cf_w_0_300_s_0_600=1.12e-11
+  mcm3m1_ca_w_0_300_s_0_800=4.52e-05 mcm3m1_cc_w_0_300_s_0_800=6.31e-11 mcm3m1_cf_w_0_300_s_0_800=1.46e-11
+  mcm3m1_ca_w_0_300_s_1_000=4.52e-05 mcm3m1_cc_w_0_300_s_1_000=5.19e-11 mcm3m1_cf_w_0_300_s_1_000=1.77e-11
+  mcm3m1_ca_w_0_300_s_1_200=4.52e-05 mcm3m1_cc_w_0_300_s_1_200=4.38e-11 mcm3m1_cf_w_0_300_s_1_200=2.04e-11
+  mcm3m1_ca_w_0_300_s_2_100=4.52e-05 mcm3m1_cc_w_0_300_s_2_100=2.45e-11 mcm3m1_cf_w_0_300_s_2_100=3.05e-11
+  mcm3m1_ca_w_0_300_s_3_300=4.52e-05 mcm3m1_cc_w_0_300_s_3_300=1.46e-11 mcm3m1_cf_w_0_300_s_3_300=3.79e-11
+  mcm3m1_ca_w_0_300_s_9_000=4.52e-05 mcm3m1_cc_w_0_300_s_9_000=3.20e-12 mcm3m1_cf_w_0_300_s_9_000=4.83e-11
+  mcm3m1_ca_w_2_400_s_0_300=4.52e-05 mcm3m1_cc_w_2_400_s_0_300=1.36e-10 mcm3m1_cf_w_2_400_s_0_300=5.43e-12
+  mcm3m1_ca_w_2_400_s_0_360=4.52e-05 mcm3m1_cc_w_2_400_s_0_360=1.25e-10 mcm3m1_cf_w_2_400_s_0_360=6.65e-12
+  mcm3m1_ca_w_2_400_s_0_450=4.52e-05 mcm3m1_cc_w_2_400_s_0_450=1.11e-10 mcm3m1_cf_w_2_400_s_0_450=8.42e-12
+  mcm3m1_ca_w_2_400_s_0_600=4.52e-05 mcm3m1_cc_w_2_400_s_0_600=9.39e-11 mcm3m1_cf_w_2_400_s_0_600=1.12e-11
+  mcm3m1_ca_w_2_400_s_0_800=4.52e-05 mcm3m1_cc_w_2_400_s_0_800=7.68e-11 mcm3m1_cf_w_2_400_s_0_800=1.46e-11
+  mcm3m1_ca_w_2_400_s_1_000=4.52e-05 mcm3m1_cc_w_2_400_s_1_000=6.45e-11 mcm3m1_cf_w_2_400_s_1_000=1.77e-11
+  mcm3m1_ca_w_2_400_s_1_200=4.52e-05 mcm3m1_cc_w_2_400_s_1_200=5.56e-11 mcm3m1_cf_w_2_400_s_1_200=2.05e-11
+  mcm3m1_ca_w_2_400_s_2_100=4.52e-05 mcm3m1_cc_w_2_400_s_2_100=3.43e-11 mcm3m1_cf_w_2_400_s_2_100=3.04e-11
+  mcm3m1_ca_w_2_400_s_3_300=4.52e-05 mcm3m1_cc_w_2_400_s_3_300=2.20e-11 mcm3m1_cf_w_2_400_s_3_300=3.88e-11
+  mcm3m1_ca_w_2_400_s_9_000=4.52e-05 mcm3m1_cc_w_2_400_s_9_000=6.05e-12 mcm3m1_cf_w_2_400_s_9_000=5.29e-11
+  mcm3m2_ca_w_0_300_s_0_300=1.31e-04 mcm3m2_cc_w_0_300_s_0_300=1.07e-10 mcm3m2_cf_w_0_300_s_0_300=1.44e-11
+  mcm3m2_ca_w_0_300_s_0_360=1.31e-04 mcm3m2_cc_w_0_300_s_0_360=9.72e-11 mcm3m2_cf_w_0_300_s_0_360=1.72e-11
+  mcm3m2_ca_w_0_300_s_0_450=1.31e-04 mcm3m2_cc_w_0_300_s_0_450=8.43e-11 mcm3m2_cf_w_0_300_s_0_450=2.11e-11
+  mcm3m2_ca_w_0_300_s_0_600=1.31e-04 mcm3m2_cc_w_0_300_s_0_600=6.83e-11 mcm3m2_cf_w_0_300_s_0_600=2.66e-11
+  mcm3m2_ca_w_0_300_s_0_800=1.31e-04 mcm3m2_cc_w_0_300_s_0_800=5.36e-11 mcm3m2_cf_w_0_300_s_0_800=3.24e-11
+  mcm3m2_ca_w_0_300_s_1_000=1.31e-04 mcm3m2_cc_w_0_300_s_1_000=4.32e-11 mcm3m2_cf_w_0_300_s_1_000=3.72e-11
+  mcm3m2_ca_w_0_300_s_1_200=1.31e-04 mcm3m2_cc_w_0_300_s_1_200=3.55e-11 mcm3m2_cf_w_0_300_s_1_200=4.11e-11
+  mcm3m2_ca_w_0_300_s_2_100=1.31e-04 mcm3m2_cc_w_0_300_s_2_100=1.80e-11 mcm3m2_cf_w_0_300_s_2_100=5.31e-11
+  mcm3m2_ca_w_0_300_s_3_300=1.31e-04 mcm3m2_cc_w_0_300_s_3_300=1.01e-11 mcm3m2_cf_w_0_300_s_3_300=6.00e-11
+  mcm3m2_ca_w_0_300_s_9_000=1.31e-04 mcm3m2_cc_w_0_300_s_9_000=2.10e-12 mcm3m2_cf_w_0_300_s_9_000=6.77e-11
+  mcm3m2_ca_w_2_400_s_0_300=1.31e-04 mcm3m2_cc_w_2_400_s_0_300=1.25e-10 mcm3m2_cf_w_2_400_s_0_300=1.43e-11
+  mcm3m2_ca_w_2_400_s_0_360=1.31e-04 mcm3m2_cc_w_2_400_s_0_360=1.14e-10 mcm3m2_cf_w_2_400_s_0_360=1.72e-11
+  mcm3m2_ca_w_2_400_s_0_450=1.31e-04 mcm3m2_cc_w_2_400_s_0_450=1.01e-10 mcm3m2_cf_w_2_400_s_0_450=2.10e-11
+  mcm3m2_ca_w_2_400_s_0_600=1.31e-04 mcm3m2_cc_w_2_400_s_0_600=8.32e-11 mcm3m2_cf_w_2_400_s_0_600=2.65e-11
+  mcm3m2_ca_w_2_400_s_0_800=1.31e-04 mcm3m2_cc_w_2_400_s_0_800=6.71e-11 mcm3m2_cf_w_2_400_s_0_800=3.24e-11
+  mcm3m2_ca_w_2_400_s_1_000=1.31e-04 mcm3m2_cc_w_2_400_s_1_000=5.56e-11 mcm3m2_cf_w_2_400_s_1_000=3.72e-11
+  mcm3m2_ca_w_2_400_s_1_200=1.31e-04 mcm3m2_cc_w_2_400_s_1_200=4.73e-11 mcm3m2_cf_w_2_400_s_1_200=4.11e-11
+  mcm3m2_ca_w_2_400_s_2_100=1.31e-04 mcm3m2_cc_w_2_400_s_2_100=2.80e-11 mcm3m2_cf_w_2_400_s_2_100=5.30e-11
+  mcm3m2_ca_w_2_400_s_3_300=1.31e-04 mcm3m2_cc_w_2_400_s_3_300=1.74e-11 mcm3m2_cf_w_2_400_s_3_300=6.16e-11
+  mcm3m2_ca_w_2_400_s_9_000=1.31e-04 mcm3m2_cc_w_2_400_s_9_000=4.55e-12 mcm3m2_cf_w_2_400_s_9_000=7.38e-11
+  mcm4f_ca_w_0_300_s_0_300=1.07e-05 mcm4f_cc_w_0_300_s_0_300=1.27e-10 mcm4f_cf_w_0_300_s_0_300=1.34e-12
+  mcm4f_ca_w_0_300_s_0_360=1.07e-05 mcm4f_cc_w_0_300_s_0_360=1.18e-10 mcm4f_cf_w_0_300_s_0_360=1.65e-12
+  mcm4f_ca_w_0_300_s_0_450=1.07e-05 mcm4f_cc_w_0_300_s_0_450=1.05e-10 mcm4f_cf_w_0_300_s_0_450=2.14e-12
+  mcm4f_ca_w_0_300_s_0_600=1.07e-05 mcm4f_cc_w_0_300_s_0_600=9.01e-11 mcm4f_cf_w_0_300_s_0_600=2.93e-12
+  mcm4f_ca_w_0_300_s_0_800=1.07e-05 mcm4f_cc_w_0_300_s_0_800=7.59e-11 mcm4f_cf_w_0_300_s_0_800=3.88e-12
+  mcm4f_ca_w_0_300_s_1_000=1.07e-05 mcm4f_cc_w_0_300_s_1_000=6.54e-11 mcm4f_cf_w_0_300_s_1_000=4.86e-12
+  mcm4f_ca_w_0_300_s_1_200=1.07e-05 mcm4f_cc_w_0_300_s_1_200=5.77e-11 mcm4f_cf_w_0_300_s_1_200=5.81e-12
+  mcm4f_ca_w_0_300_s_2_100=1.07e-05 mcm4f_cc_w_0_300_s_2_100=3.87e-11 mcm4f_cf_w_0_300_s_2_100=9.97e-12
+  mcm4f_ca_w_0_300_s_3_300=1.07e-05 mcm4f_cc_w_0_300_s_3_300=2.73e-11 mcm4f_cf_w_0_300_s_3_300=1.43e-11
+  mcm4f_ca_w_0_300_s_9_000=1.07e-05 mcm4f_cc_w_0_300_s_9_000=9.06e-12 mcm4f_cf_w_0_300_s_9_000=2.67e-11
+  mcm4f_ca_w_2_400_s_0_300=1.07e-05 mcm4f_cc_w_2_400_s_0_300=1.56e-10 mcm4f_cf_w_2_400_s_0_300=1.37e-12
+  mcm4f_ca_w_2_400_s_0_360=1.07e-05 mcm4f_cc_w_2_400_s_0_360=1.45e-10 mcm4f_cf_w_2_400_s_0_360=1.68e-12
+  mcm4f_ca_w_2_400_s_0_450=1.07e-05 mcm4f_cc_w_2_400_s_0_450=1.31e-10 mcm4f_cf_w_2_400_s_0_450=2.15e-12
+  mcm4f_ca_w_2_400_s_0_600=1.07e-05 mcm4f_cc_w_2_400_s_0_600=1.14e-10 mcm4f_cf_w_2_400_s_0_600=2.92e-12
+  mcm4f_ca_w_2_400_s_0_800=1.07e-05 mcm4f_cc_w_2_400_s_0_800=9.60e-11 mcm4f_cf_w_2_400_s_0_800=3.92e-12
+  mcm4f_ca_w_2_400_s_1_000=1.07e-05 mcm4f_cc_w_2_400_s_1_000=8.34e-11 mcm4f_cf_w_2_400_s_1_000=4.92e-12
+  mcm4f_ca_w_2_400_s_1_200=1.07e-05 mcm4f_cc_w_2_400_s_1_200=7.40e-11 mcm4f_cf_w_2_400_s_1_200=5.88e-12
+  mcm4f_ca_w_2_400_s_2_100=1.07e-05 mcm4f_cc_w_2_400_s_2_100=5.05e-11 mcm4f_cf_w_2_400_s_2_100=9.95e-12
+  mcm4f_ca_w_2_400_s_3_300=1.07e-05 mcm4f_cc_w_2_400_s_3_300=3.61e-11 mcm4f_cf_w_2_400_s_3_300=1.47e-11
+  mcm4f_ca_w_2_400_s_9_000=1.07e-05 mcm4f_cc_w_2_400_s_9_000=1.32e-11 mcm4f_cf_w_2_400_s_9_000=2.89e-11
+  mcm4d_ca_w_0_300_s_0_300=1.14e-05 mcm4d_cc_w_0_300_s_0_300=1.27e-10 mcm4d_cf_w_0_300_s_0_300=1.43e-12
+  mcm4d_ca_w_0_300_s_0_360=1.14e-05 mcm4d_cc_w_0_300_s_0_360=1.17e-10 mcm4d_cf_w_0_300_s_0_360=1.77e-12
+  mcm4d_ca_w_0_300_s_0_450=1.14e-05 mcm4d_cc_w_0_300_s_0_450=1.05e-10 mcm4d_cf_w_0_300_s_0_450=2.28e-12
+  mcm4d_ca_w_0_300_s_0_600=1.14e-05 mcm4d_cc_w_0_300_s_0_600=8.98e-11 mcm4d_cf_w_0_300_s_0_600=3.13e-12
+  mcm4d_ca_w_0_300_s_0_800=1.14e-05 mcm4d_cc_w_0_300_s_0_800=7.56e-11 mcm4d_cf_w_0_300_s_0_800=4.14e-12
+  mcm4d_ca_w_0_300_s_1_000=1.14e-05 mcm4d_cc_w_0_300_s_1_000=6.51e-11 mcm4d_cf_w_0_300_s_1_000=5.18e-12
+  mcm4d_ca_w_0_300_s_1_200=1.14e-05 mcm4d_cc_w_0_300_s_1_200=5.73e-11 mcm4d_cf_w_0_300_s_1_200=6.19e-12
+  mcm4d_ca_w_0_300_s_2_100=1.14e-05 mcm4d_cc_w_0_300_s_2_100=3.82e-11 mcm4d_cf_w_0_300_s_2_100=1.06e-11
+  mcm4d_ca_w_0_300_s_3_300=1.14e-05 mcm4d_cc_w_0_300_s_3_300=2.68e-11 mcm4d_cf_w_0_300_s_3_300=1.52e-11
+  mcm4d_ca_w_0_300_s_9_000=1.14e-05 mcm4d_cc_w_0_300_s_9_000=8.65e-12 mcm4d_cf_w_0_300_s_9_000=2.77e-11
+  mcm4d_ca_w_2_400_s_0_300=1.14e-05 mcm4d_cc_w_2_400_s_0_300=1.56e-10 mcm4d_cf_w_2_400_s_0_300=1.46e-12
+  mcm4d_ca_w_2_400_s_0_360=1.14e-05 mcm4d_cc_w_2_400_s_0_360=1.45e-10 mcm4d_cf_w_2_400_s_0_360=1.80e-12
+  mcm4d_ca_w_2_400_s_0_450=1.14e-05 mcm4d_cc_w_2_400_s_0_450=1.31e-10 mcm4d_cf_w_2_400_s_0_450=2.30e-12
+  mcm4d_ca_w_2_400_s_0_600=1.14e-05 mcm4d_cc_w_2_400_s_0_600=1.13e-10 mcm4d_cf_w_2_400_s_0_600=3.12e-12
+  mcm4d_ca_w_2_400_s_0_800=1.14e-05 mcm4d_cc_w_2_400_s_0_800=9.54e-11 mcm4d_cf_w_2_400_s_0_800=4.19e-12
+  mcm4d_ca_w_2_400_s_1_000=1.14e-05 mcm4d_cc_w_2_400_s_1_000=8.28e-11 mcm4d_cf_w_2_400_s_1_000=5.24e-12
+  mcm4d_ca_w_2_400_s_1_200=1.14e-05 mcm4d_cc_w_2_400_s_1_200=7.33e-11 mcm4d_cf_w_2_400_s_1_200=6.27e-12
+  mcm4d_ca_w_2_400_s_2_100=1.14e-05 mcm4d_cc_w_2_400_s_2_100=4.98e-11 mcm4d_cf_w_2_400_s_2_100=1.06e-11
+  mcm4d_ca_w_2_400_s_3_300=1.14e-05 mcm4d_cc_w_2_400_s_3_300=3.54e-11 mcm4d_cf_w_2_400_s_3_300=1.56e-11
+  mcm4d_ca_w_2_400_s_9_000=1.14e-05 mcm4d_cc_w_2_400_s_9_000=1.26e-11 mcm4d_cf_w_2_400_s_9_000=3.00e-11
+  mcm4p1_ca_w_0_300_s_0_300=1.26e-05 mcm4p1_cc_w_0_300_s_0_300=1.27e-10 mcm4p1_cf_w_0_300_s_0_300=1.58e-12
+  mcm4p1_ca_w_0_300_s_0_360=1.26e-05 mcm4p1_cc_w_0_300_s_0_360=1.17e-10 mcm4p1_cf_w_0_300_s_0_360=1.96e-12
+  mcm4p1_ca_w_0_300_s_0_450=1.26e-05 mcm4p1_cc_w_0_300_s_0_450=1.05e-10 mcm4p1_cf_w_0_300_s_0_450=2.52e-12
+  mcm4p1_ca_w_0_300_s_0_600=1.26e-05 mcm4p1_cc_w_0_300_s_0_600=8.94e-11 mcm4p1_cf_w_0_300_s_0_600=3.45e-12
+  mcm4p1_ca_w_0_300_s_0_800=1.26e-05 mcm4p1_cc_w_0_300_s_0_800=7.51e-11 mcm4p1_cf_w_0_300_s_0_800=4.57e-12
+  mcm4p1_ca_w_0_300_s_1_000=1.26e-05 mcm4p1_cc_w_0_300_s_1_000=6.45e-11 mcm4p1_cf_w_0_300_s_1_000=5.70e-12
+  mcm4p1_ca_w_0_300_s_1_200=1.26e-05 mcm4p1_cc_w_0_300_s_1_200=5.67e-11 mcm4p1_cf_w_0_300_s_1_200=6.81e-12
+  mcm4p1_ca_w_0_300_s_2_100=1.26e-05 mcm4p1_cc_w_0_300_s_2_100=3.74e-11 mcm4p1_cf_w_0_300_s_2_100=1.15e-11
+  mcm4p1_ca_w_0_300_s_3_300=1.26e-05 mcm4p1_cc_w_0_300_s_3_300=2.59e-11 mcm4p1_cf_w_0_300_s_3_300=1.65e-11
+  mcm4p1_ca_w_0_300_s_9_000=1.26e-05 mcm4p1_cc_w_0_300_s_9_000=8.02e-12 mcm4p1_cf_w_0_300_s_9_000=2.92e-11
+  mcm4p1_ca_w_2_400_s_0_300=1.26e-05 mcm4p1_cc_w_2_400_s_0_300=1.55e-10 mcm4p1_cf_w_2_400_s_0_300=1.63e-12
+  mcm4p1_ca_w_2_400_s_0_360=1.26e-05 mcm4p1_cc_w_2_400_s_0_360=1.44e-10 mcm4p1_cf_w_2_400_s_0_360=2.00e-12
+  mcm4p1_ca_w_2_400_s_0_450=1.26e-05 mcm4p1_cc_w_2_400_s_0_450=1.30e-10 mcm4p1_cf_w_2_400_s_0_450=2.55e-12
+  mcm4p1_ca_w_2_400_s_0_600=1.26e-05 mcm4p1_cc_w_2_400_s_0_600=1.12e-10 mcm4p1_cf_w_2_400_s_0_600=3.46e-12
+  mcm4p1_ca_w_2_400_s_0_800=1.26e-05 mcm4p1_cc_w_2_400_s_0_800=9.44e-11 mcm4p1_cf_w_2_400_s_0_800=4.62e-12
+  mcm4p1_ca_w_2_400_s_1_000=1.26e-05 mcm4p1_cc_w_2_400_s_1_000=8.18e-11 mcm4p1_cf_w_2_400_s_1_000=5.79e-12
+  mcm4p1_ca_w_2_400_s_1_200=1.26e-05 mcm4p1_cc_w_2_400_s_1_200=7.23e-11 mcm4p1_cf_w_2_400_s_1_200=6.91e-12
+  mcm4p1_ca_w_2_400_s_2_100=1.26e-05 mcm4p1_cc_w_2_400_s_2_100=4.88e-11 mcm4p1_cf_w_2_400_s_2_100=1.16e-11
+  mcm4p1_ca_w_2_400_s_3_300=1.26e-05 mcm4p1_cc_w_2_400_s_3_300=3.44e-11 mcm4p1_cf_w_2_400_s_3_300=1.69e-11
+  mcm4p1_ca_w_2_400_s_9_000=1.26e-05 mcm4p1_cc_w_2_400_s_9_000=1.19e-11 mcm4p1_cf_w_2_400_s_9_000=3.18e-11
+  mcm4l1_ca_w_0_300_s_0_300=1.43e-05 mcm4l1_cc_w_0_300_s_0_300=1.26e-10 mcm4l1_cf_w_0_300_s_0_300=1.77e-12
+  mcm4l1_ca_w_0_300_s_0_360=1.43e-05 mcm4l1_cc_w_0_300_s_0_360=1.17e-10 mcm4l1_cf_w_0_300_s_0_360=2.19e-12
+  mcm4l1_ca_w_0_300_s_0_450=1.43e-05 mcm4l1_cc_w_0_300_s_0_450=1.04e-10 mcm4l1_cf_w_0_300_s_0_450=2.82e-12
+  mcm4l1_ca_w_0_300_s_0_600=1.43e-05 mcm4l1_cc_w_0_300_s_0_600=8.89e-11 mcm4l1_cf_w_0_300_s_0_600=3.86e-12
+  mcm4l1_ca_w_0_300_s_0_800=1.43e-05 mcm4l1_cc_w_0_300_s_0_800=7.45e-11 mcm4l1_cf_w_0_300_s_0_800=5.11e-12
+  mcm4l1_ca_w_0_300_s_1_000=1.43e-05 mcm4l1_cc_w_0_300_s_1_000=6.38e-11 mcm4l1_cf_w_0_300_s_1_000=6.37e-12
+  mcm4l1_ca_w_0_300_s_1_200=1.43e-05 mcm4l1_cc_w_0_300_s_1_200=5.59e-11 mcm4l1_cf_w_0_300_s_1_200=7.60e-12
+  mcm4l1_ca_w_0_300_s_2_100=1.43e-05 mcm4l1_cc_w_0_300_s_2_100=3.64e-11 mcm4l1_cf_w_0_300_s_2_100=1.28e-11
+  mcm4l1_ca_w_0_300_s_3_300=1.43e-05 mcm4l1_cc_w_0_300_s_3_300=2.49e-11 mcm4l1_cf_w_0_300_s_3_300=1.80e-11
+  mcm4l1_ca_w_0_300_s_9_000=1.43e-05 mcm4l1_cc_w_0_300_s_9_000=7.33e-12 mcm4l1_cf_w_0_300_s_9_000=3.10e-11
+  mcm4l1_ca_w_2_400_s_0_300=1.43e-05 mcm4l1_cc_w_2_400_s_0_300=1.54e-10 mcm4l1_cf_w_2_400_s_0_300=1.79e-12
+  mcm4l1_ca_w_2_400_s_0_360=1.43e-05 mcm4l1_cc_w_2_400_s_0_360=1.43e-10 mcm4l1_cf_w_2_400_s_0_360=2.20e-12
+  mcm4l1_ca_w_2_400_s_0_450=1.43e-05 mcm4l1_cc_w_2_400_s_0_450=1.29e-10 mcm4l1_cf_w_2_400_s_0_450=2.82e-12
+  mcm4l1_ca_w_2_400_s_0_600=1.43e-05 mcm4l1_cc_w_2_400_s_0_600=1.11e-10 mcm4l1_cf_w_2_400_s_0_600=3.84e-12
+  mcm4l1_ca_w_2_400_s_0_800=1.43e-05 mcm4l1_cc_w_2_400_s_0_800=9.32e-11 mcm4l1_cf_w_2_400_s_0_800=5.15e-12
+  mcm4l1_ca_w_2_400_s_1_000=1.43e-05 mcm4l1_cc_w_2_400_s_1_000=8.05e-11 mcm4l1_cf_w_2_400_s_1_000=6.43e-12
+  mcm4l1_ca_w_2_400_s_1_200=1.43e-05 mcm4l1_cc_w_2_400_s_1_200=7.11e-11 mcm4l1_cf_w_2_400_s_1_200=7.67e-12
+  mcm4l1_ca_w_2_400_s_2_100=1.43e-05 mcm4l1_cc_w_2_400_s_2_100=4.77e-11 mcm4l1_cf_w_2_400_s_2_100=1.28e-11
+  mcm4l1_ca_w_2_400_s_3_300=1.43e-05 mcm4l1_cc_w_2_400_s_3_300=3.32e-11 mcm4l1_cf_w_2_400_s_3_300=1.85e-11
+  mcm4l1_ca_w_2_400_s_9_000=1.43e-05 mcm4l1_cc_w_2_400_s_9_000=1.11e-11 mcm4l1_cf_w_2_400_s_9_000=3.37e-11
+  mcm4m1_ca_w_0_300_s_0_300=1.85e-05 mcm4m1_cc_w_0_300_s_0_300=1.25e-10 mcm4m1_cf_w_0_300_s_0_300=2.28e-12
+  mcm4m1_ca_w_0_300_s_0_360=1.85e-05 mcm4m1_cc_w_0_300_s_0_360=1.16e-10 mcm4m1_cf_w_0_300_s_0_360=2.81e-12
+  mcm4m1_ca_w_0_300_s_0_450=1.85e-05 mcm4m1_cc_w_0_300_s_0_450=1.03e-10 mcm4m1_cf_w_0_300_s_0_450=3.62e-12
+  mcm4m1_ca_w_0_300_s_0_600=1.85e-05 mcm4m1_cc_w_0_300_s_0_600=8.73e-11 mcm4m1_cf_w_0_300_s_0_600=4.92e-12
+  mcm4m1_ca_w_0_300_s_0_800=1.85e-05 mcm4m1_cc_w_0_300_s_0_800=7.29e-11 mcm4m1_cf_w_0_300_s_0_800=6.51e-12
+  mcm4m1_ca_w_0_300_s_1_000=1.85e-05 mcm4m1_cc_w_0_300_s_1_000=6.21e-11 mcm4m1_cf_w_0_300_s_1_000=8.10e-12
+  mcm4m1_ca_w_0_300_s_1_200=1.85e-05 mcm4m1_cc_w_0_300_s_1_200=5.40e-11 mcm4m1_cf_w_0_300_s_1_200=9.59e-12
+  mcm4m1_ca_w_0_300_s_2_100=1.85e-05 mcm4m1_cc_w_0_300_s_2_100=3.42e-11 mcm4m1_cf_w_0_300_s_2_100=1.58e-11
+  mcm4m1_ca_w_0_300_s_3_300=1.85e-05 mcm4m1_cc_w_0_300_s_3_300=2.27e-11 mcm4m1_cf_w_0_300_s_3_300=2.19e-11
+  mcm4m1_ca_w_0_300_s_9_000=1.85e-05 mcm4m1_cc_w_0_300_s_9_000=6.13e-12 mcm4m1_cf_w_0_300_s_9_000=3.49e-11
+  mcm4m1_ca_w_2_400_s_0_300=1.85e-05 mcm4m1_cc_w_2_400_s_0_300=1.51e-10 mcm4m1_cf_w_2_400_s_0_300=2.28e-12
+  mcm4m1_ca_w_2_400_s_0_360=1.85e-05 mcm4m1_cc_w_2_400_s_0_360=1.40e-10 mcm4m1_cf_w_2_400_s_0_360=2.82e-12
+  mcm4m1_ca_w_2_400_s_0_450=1.85e-05 mcm4m1_cc_w_2_400_s_0_450=1.26e-10 mcm4m1_cf_w_2_400_s_0_450=3.60e-12
+  mcm4m1_ca_w_2_400_s_0_600=1.85e-05 mcm4m1_cc_w_2_400_s_0_600=1.08e-10 mcm4m1_cf_w_2_400_s_0_600=4.89e-12
+  mcm4m1_ca_w_2_400_s_0_800=1.85e-05 mcm4m1_cc_w_2_400_s_0_800=9.06e-11 mcm4m1_cf_w_2_400_s_0_800=6.54e-12
+  mcm4m1_ca_w_2_400_s_1_000=1.85e-05 mcm4m1_cc_w_2_400_s_1_000=7.79e-11 mcm4m1_cf_w_2_400_s_1_000=8.15e-12
+  mcm4m1_ca_w_2_400_s_1_200=1.85e-05 mcm4m1_cc_w_2_400_s_1_200=6.84e-11 mcm4m1_cf_w_2_400_s_1_200=9.67e-12
+  mcm4m1_ca_w_2_400_s_2_100=1.85e-05 mcm4m1_cc_w_2_400_s_2_100=4.50e-11 mcm4m1_cf_w_2_400_s_2_100=1.58e-11
+  mcm4m1_ca_w_2_400_s_3_300=1.85e-05 mcm4m1_cc_w_2_400_s_3_300=3.07e-11 mcm4m1_cf_w_2_400_s_3_300=2.25e-11
+  mcm4m1_ca_w_2_400_s_9_000=1.85e-05 mcm4m1_cc_w_2_400_s_9_000=9.60e-12 mcm4m1_cf_w_2_400_s_9_000=3.81e-11
+  mcm4m2_ca_w_0_300_s_0_300=2.52e-05 mcm4m2_cc_w_0_300_s_0_300=1.24e-10 mcm4m2_cf_w_0_300_s_0_300=3.09e-12
+  mcm4m2_ca_w_0_300_s_0_360=2.52e-05 mcm4m2_cc_w_0_300_s_0_360=1.13e-10 mcm4m2_cf_w_0_300_s_0_360=3.81e-12
+  mcm4m2_ca_w_0_300_s_0_450=2.52e-05 mcm4m2_cc_w_0_300_s_0_450=1.01e-10 mcm4m2_cf_w_0_300_s_0_450=4.87e-12
+  mcm4m2_ca_w_0_300_s_0_600=2.52e-05 mcm4m2_cc_w_0_300_s_0_600=8.53e-11 mcm4m2_cf_w_0_300_s_0_600=6.59e-12
+  mcm4m2_ca_w_0_300_s_0_800=2.52e-05 mcm4m2_cc_w_0_300_s_0_800=7.05e-11 mcm4m2_cf_w_0_300_s_0_800=8.69e-12
+  mcm4m2_ca_w_0_300_s_1_000=2.52e-05 mcm4m2_cc_w_0_300_s_1_000=5.97e-11 mcm4m2_cf_w_0_300_s_1_000=1.08e-11
+  mcm4m2_ca_w_0_300_s_1_200=2.52e-05 mcm4m2_cc_w_0_300_s_1_200=5.15e-11 mcm4m2_cf_w_0_300_s_1_200=1.27e-11
+  mcm4m2_ca_w_0_300_s_2_100=2.52e-05 mcm4m2_cc_w_0_300_s_2_100=3.15e-11 mcm4m2_cf_w_0_300_s_2_100=2.03e-11
+  mcm4m2_ca_w_0_300_s_3_300=2.52e-05 mcm4m2_cc_w_0_300_s_3_300=2.01e-11 mcm4m2_cf_w_0_300_s_3_300=2.71e-11
+  mcm4m2_ca_w_0_300_s_9_000=2.52e-05 mcm4m2_cc_w_0_300_s_9_000=4.87e-12 mcm4m2_cf_w_0_300_s_9_000=3.99e-11
+  mcm4m2_ca_w_2_400_s_0_300=2.52e-05 mcm4m2_cc_w_2_400_s_0_300=1.48e-10 mcm4m2_cf_w_2_400_s_0_300=3.10e-12
+  mcm4m2_ca_w_2_400_s_0_360=2.52e-05 mcm4m2_cc_w_2_400_s_0_360=1.37e-10 mcm4m2_cf_w_2_400_s_0_360=3.81e-12
+  mcm4m2_ca_w_2_400_s_0_450=2.52e-05 mcm4m2_cc_w_2_400_s_0_450=1.23e-10 mcm4m2_cf_w_2_400_s_0_450=4.86e-12
+  mcm4m2_ca_w_2_400_s_0_600=2.52e-05 mcm4m2_cc_w_2_400_s_0_600=1.05e-10 mcm4m2_cf_w_2_400_s_0_600=6.57e-12
+  mcm4m2_ca_w_2_400_s_0_800=2.52e-05 mcm4m2_cc_w_2_400_s_0_800=8.72e-11 mcm4m2_cf_w_2_400_s_0_800=8.73e-12
+  mcm4m2_ca_w_2_400_s_1_000=2.52e-05 mcm4m2_cc_w_2_400_s_1_000=7.45e-11 mcm4m2_cf_w_2_400_s_1_000=1.08e-11
+  mcm4m2_ca_w_2_400_s_1_200=2.52e-05 mcm4m2_cc_w_2_400_s_1_200=6.51e-11 mcm4m2_cf_w_2_400_s_1_200=1.27e-11
+  mcm4m2_ca_w_2_400_s_2_100=2.52e-05 mcm4m2_cc_w_2_400_s_2_100=4.19e-11 mcm4m2_cf_w_2_400_s_2_100=2.03e-11
+  mcm4m2_ca_w_2_400_s_3_300=2.52e-05 mcm4m2_cc_w_2_400_s_3_300=2.79e-11 mcm4m2_cf_w_2_400_s_3_300=2.78e-11
+  mcm4m2_ca_w_2_400_s_9_000=2.52e-05 mcm4m2_cc_w_2_400_s_9_000=8.10e-12 mcm4m2_cf_w_2_400_s_9_000=4.36e-11
+  mcm4m3_ca_w_0_300_s_0_300=1.91e-04 mcm4m3_cc_w_0_300_s_0_300=1.05e-10 mcm4m3_cf_w_0_300_s_0_300=1.96e-11
+  mcm4m3_ca_w_0_300_s_0_360=1.91e-04 mcm4m3_cc_w_0_300_s_0_360=9.56e-11 mcm4m3_cf_w_0_300_s_0_360=2.31e-11
+  mcm4m3_ca_w_0_300_s_0_450=1.91e-04 mcm4m3_cc_w_0_300_s_0_450=8.29e-11 mcm4m3_cf_w_0_300_s_0_450=2.78e-11
+  mcm4m3_ca_w_0_300_s_0_600=1.91e-04 mcm4m3_cc_w_0_300_s_0_600=6.76e-11 mcm4m3_cf_w_0_300_s_0_600=3.42e-11
+  mcm4m3_ca_w_0_300_s_0_800=1.91e-04 mcm4m3_cc_w_0_300_s_0_800=5.35e-11 mcm4m3_cf_w_0_300_s_0_800=4.07e-11
+  mcm4m3_ca_w_0_300_s_1_000=1.91e-04 mcm4m3_cc_w_0_300_s_1_000=4.33e-11 mcm4m3_cf_w_0_300_s_1_000=4.56e-11
+  mcm4m3_ca_w_0_300_s_1_200=1.91e-04 mcm4m3_cc_w_0_300_s_1_200=3.59e-11 mcm4m3_cf_w_0_300_s_1_200=4.97e-11
+  mcm4m3_ca_w_0_300_s_2_100=1.91e-04 mcm4m3_cc_w_0_300_s_2_100=1.86e-11 mcm4m3_cf_w_0_300_s_2_100=6.19e-11
+  mcm4m3_ca_w_0_300_s_3_300=1.91e-04 mcm4m3_cc_w_0_300_s_3_300=1.05e-11 mcm4m3_cf_w_0_300_s_3_300=6.90e-11
+  mcm4m3_ca_w_0_300_s_9_000=1.91e-04 mcm4m3_cc_w_0_300_s_9_000=2.00e-12 mcm4m3_cf_w_0_300_s_9_000=7.72e-11
+  mcm4m3_ca_w_2_400_s_0_300=1.91e-04 mcm4m3_cc_w_2_400_s_0_300=1.26e-10 mcm4m3_cf_w_2_400_s_0_300=1.96e-11
+  mcm4m3_ca_w_2_400_s_0_360=1.91e-04 mcm4m3_cc_w_2_400_s_0_360=1.15e-10 mcm4m3_cf_w_2_400_s_0_360=2.31e-11
+  mcm4m3_ca_w_2_400_s_0_450=1.91e-04 mcm4m3_cc_w_2_400_s_0_450=1.02e-10 mcm4m3_cf_w_2_400_s_0_450=2.78e-11
+  mcm4m3_ca_w_2_400_s_0_600=1.91e-04 mcm4m3_cc_w_2_400_s_0_600=8.47e-11 mcm4m3_cf_w_2_400_s_0_600=3.41e-11
+  mcm4m3_ca_w_2_400_s_0_800=1.91e-04 mcm4m3_cc_w_2_400_s_0_800=6.87e-11 mcm4m3_cf_w_2_400_s_0_800=4.06e-11
+  mcm4m3_ca_w_2_400_s_1_000=1.91e-04 mcm4m3_cc_w_2_400_s_1_000=5.73e-11 mcm4m3_cf_w_2_400_s_1_000=4.58e-11
+  mcm4m3_ca_w_2_400_s_1_200=1.91e-04 mcm4m3_cc_w_2_400_s_1_200=4.89e-11 mcm4m3_cf_w_2_400_s_1_200=4.99e-11
+  mcm4m3_ca_w_2_400_s_2_100=1.91e-04 mcm4m3_cc_w_2_400_s_2_100=2.91e-11 mcm4m3_cf_w_2_400_s_2_100=6.21e-11
+  mcm4m3_ca_w_2_400_s_3_300=1.91e-04 mcm4m3_cc_w_2_400_s_3_300=1.78e-11 mcm4m3_cf_w_2_400_s_3_300=7.11e-11
+  mcm4m3_ca_w_2_400_s_9_000=1.91e-04 mcm4m3_cc_w_2_400_s_9_000=4.30e-12 mcm4m3_cf_w_2_400_s_9_000=8.40e-11
+  mcm5f_ca_w_1_600_s_1_600=7.76e-06 mcm5f_cc_w_1_600_s_1_600=8.87e-11 mcm5f_cf_w_1_600_s_1_600=5.58e-12
+  mcm5f_ca_w_1_600_s_1_700=7.76e-06 mcm5f_cc_w_1_600_s_1_700=8.37e-11 mcm5f_cf_w_1_600_s_1_700=5.94e-12
+  mcm5f_ca_w_1_600_s_1_900=7.76e-06 mcm5f_cc_w_1_600_s_1_900=7.54e-11 mcm5f_cf_w_1_600_s_1_900=6.64e-12
+  mcm5f_ca_w_1_600_s_2_000=7.76e-06 mcm5f_cc_w_1_600_s_2_000=7.20e-11 mcm5f_cf_w_1_600_s_2_000=7.00e-12
+  mcm5f_ca_w_1_600_s_2_400=7.76e-06 mcm5f_cc_w_1_600_s_2_400=6.13e-11 mcm5f_cf_w_1_600_s_2_400=8.37e-12
+  mcm5f_ca_w_1_600_s_2_800=7.76e-06 mcm5f_cc_w_1_600_s_2_800=5.36e-11 mcm5f_cf_w_1_600_s_2_800=9.71e-12
+  mcm5f_ca_w_1_600_s_3_200=7.76e-06 mcm5f_cc_w_1_600_s_3_200=4.77e-11 mcm5f_cf_w_1_600_s_3_200=1.10e-11
+  mcm5f_ca_w_1_600_s_4_800=7.76e-06 mcm5f_cc_w_1_600_s_4_800=3.33e-11 mcm5f_cf_w_1_600_s_4_800=1.57e-11
+  mcm5f_ca_w_1_600_s_10_000=7.76e-06 mcm5f_cc_w_1_600_s_10_000=1.52e-11 mcm5f_cf_w_1_600_s_10_000=2.64e-11
+  mcm5f_ca_w_1_600_s_12_000=7.76e-06 mcm5f_cc_w_1_600_s_12_000=1.20e-11 mcm5f_cf_w_1_600_s_12_000=2.89e-11
+  mcm5f_ca_w_4_000_s_1_600=7.76e-06 mcm5f_cc_w_4_000_s_1_600=9.55e-11 mcm5f_cf_w_4_000_s_1_600=5.59e-12
+  mcm5f_ca_w_4_000_s_1_700=7.76e-06 mcm5f_cc_w_4_000_s_1_700=9.04e-11 mcm5f_cf_w_4_000_s_1_700=5.95e-12
+  mcm5f_ca_w_4_000_s_1_900=7.76e-06 mcm5f_cc_w_4_000_s_1_900=8.19e-11 mcm5f_cf_w_4_000_s_1_900=6.66e-12
+  mcm5f_ca_w_4_000_s_2_000=7.76e-06 mcm5f_cc_w_4_000_s_2_000=7.82e-11 mcm5f_cf_w_4_000_s_2_000=7.01e-12
+  mcm5f_ca_w_4_000_s_2_400=7.76e-06 mcm5f_cc_w_4_000_s_2_400=6.71e-11 mcm5f_cf_w_4_000_s_2_400=8.39e-12
+  mcm5f_ca_w_4_000_s_2_800=7.76e-06 mcm5f_cc_w_4_000_s_2_800=5.89e-11 mcm5f_cf_w_4_000_s_2_800=9.73e-12
+  mcm5f_ca_w_4_000_s_3_200=7.76e-06 mcm5f_cc_w_4_000_s_3_200=5.27e-11 mcm5f_cf_w_4_000_s_3_200=1.10e-11
+  mcm5f_ca_w_4_000_s_4_800=7.76e-06 mcm5f_cc_w_4_000_s_4_800=3.73e-11 mcm5f_cf_w_4_000_s_4_800=1.58e-11
+  mcm5f_ca_w_4_000_s_10_000=7.76e-06 mcm5f_cc_w_4_000_s_10_000=1.78e-11 mcm5f_cf_w_4_000_s_10_000=2.68e-11
+  mcm5f_ca_w_4_000_s_12_000=7.76e-06 mcm5f_cc_w_4_000_s_12_000=1.43e-11 mcm5f_cf_w_4_000_s_12_000=2.95e-11
+  mcm5d_ca_w_1_600_s_1_600=8.14e-06 mcm5d_cc_w_1_600_s_1_600=8.83e-11 mcm5d_cf_w_1_600_s_1_600=5.85e-12
+  mcm5d_ca_w_1_600_s_1_700=8.14e-06 mcm5d_cc_w_1_600_s_1_700=8.33e-11 mcm5d_cf_w_1_600_s_1_700=6.22e-12
+  mcm5d_ca_w_1_600_s_1_900=8.14e-06 mcm5d_cc_w_1_600_s_1_900=7.50e-11 mcm5d_cf_w_1_600_s_1_900=6.96e-12
+  mcm5d_ca_w_1_600_s_2_000=8.14e-06 mcm5d_cc_w_1_600_s_2_000=7.16e-11 mcm5d_cf_w_1_600_s_2_000=7.32e-12
+  mcm5d_ca_w_1_600_s_2_400=8.14e-06 mcm5d_cc_w_1_600_s_2_400=6.08e-11 mcm5d_cf_w_1_600_s_2_400=8.76e-12
+  mcm5d_ca_w_1_600_s_2_800=8.14e-06 mcm5d_cc_w_1_600_s_2_800=5.31e-11 mcm5d_cf_w_1_600_s_2_800=1.02e-11
+  mcm5d_ca_w_1_600_s_3_200=8.14e-06 mcm5d_cc_w_1_600_s_3_200=4.73e-11 mcm5d_cf_w_1_600_s_3_200=1.15e-11
+  mcm5d_ca_w_1_600_s_4_800=8.14e-06 mcm5d_cc_w_1_600_s_4_800=3.28e-11 mcm5d_cf_w_1_600_s_4_800=1.64e-11
+  mcm5d_ca_w_1_600_s_10_000=8.14e-06 mcm5d_cc_w_1_600_s_10_000=1.48e-11 mcm5d_cf_w_1_600_s_10_000=2.72e-11
+  mcm5d_ca_w_1_600_s_12_000=8.14e-06 mcm5d_cc_w_1_600_s_12_000=1.16e-11 mcm5d_cf_w_1_600_s_12_000=2.98e-11
+  mcm5d_ca_w_4_000_s_1_600=8.14e-06 mcm5d_cc_w_4_000_s_1_600=9.51e-11 mcm5d_cf_w_4_000_s_1_600=5.85e-12
+  mcm5d_ca_w_4_000_s_1_700=8.14e-06 mcm5d_cc_w_4_000_s_1_700=8.98e-11 mcm5d_cf_w_4_000_s_1_700=6.22e-12
+  mcm5d_ca_w_4_000_s_1_900=8.14e-06 mcm5d_cc_w_4_000_s_1_900=8.14e-11 mcm5d_cf_w_4_000_s_1_900=6.97e-12
+  mcm5d_ca_w_4_000_s_2_000=8.14e-06 mcm5d_cc_w_4_000_s_2_000=7.77e-11 mcm5d_cf_w_4_000_s_2_000=7.33e-12
+  mcm5d_ca_w_4_000_s_2_400=8.14e-06 mcm5d_cc_w_4_000_s_2_400=6.65e-11 mcm5d_cf_w_4_000_s_2_400=8.77e-12
+  mcm5d_ca_w_4_000_s_2_800=8.14e-06 mcm5d_cc_w_4_000_s_2_800=5.84e-11 mcm5d_cf_w_4_000_s_2_800=1.02e-11
+  mcm5d_ca_w_4_000_s_3_200=8.14e-06 mcm5d_cc_w_4_000_s_3_200=5.22e-11 mcm5d_cf_w_4_000_s_3_200=1.15e-11
+  mcm5d_ca_w_4_000_s_4_800=8.14e-06 mcm5d_cc_w_4_000_s_4_800=3.68e-11 mcm5d_cf_w_4_000_s_4_800=1.64e-11
+  mcm5d_ca_w_4_000_s_10_000=8.14e-06 mcm5d_cc_w_4_000_s_10_000=1.74e-11 mcm5d_cf_w_4_000_s_10_000=2.76e-11
+  mcm5d_ca_w_4_000_s_12_000=8.14e-06 mcm5d_cc_w_4_000_s_12_000=1.40e-11 mcm5d_cf_w_4_000_s_12_000=3.04e-11
+  mcm5p1_ca_w_1_600_s_1_600=8.74e-06 mcm5p1_cc_w_1_600_s_1_600=8.77e-11 mcm5p1_cf_w_1_600_s_1_600=6.26e-12
+  mcm5p1_ca_w_1_600_s_1_700=8.74e-06 mcm5p1_cc_w_1_600_s_1_700=8.27e-11 mcm5p1_cf_w_1_600_s_1_700=6.66e-12
+  mcm5p1_ca_w_1_600_s_1_900=8.74e-06 mcm5p1_cc_w_1_600_s_1_900=7.43e-11 mcm5p1_cf_w_1_600_s_1_900=7.44e-12
+  mcm5p1_ca_w_1_600_s_2_000=8.74e-06 mcm5p1_cc_w_1_600_s_2_000=7.10e-11 mcm5p1_cf_w_1_600_s_2_000=7.83e-12
+  mcm5p1_ca_w_1_600_s_2_400=8.74e-06 mcm5p1_cc_w_1_600_s_2_400=6.02e-11 mcm5p1_cf_w_1_600_s_2_400=9.36e-12
+  mcm5p1_ca_w_1_600_s_2_800=8.74e-06 mcm5p1_cc_w_1_600_s_2_800=5.24e-11 mcm5p1_cf_w_1_600_s_2_800=1.08e-11
+  mcm5p1_ca_w_1_600_s_3_200=8.74e-06 mcm5p1_cc_w_1_600_s_3_200=4.66e-11 mcm5p1_cf_w_1_600_s_3_200=1.22e-11
+  mcm5p1_ca_w_1_600_s_4_800=8.74e-06 mcm5p1_cc_w_1_600_s_4_800=3.21e-11 mcm5p1_cf_w_1_600_s_4_800=1.74e-11
+  mcm5p1_ca_w_1_600_s_10_000=8.74e-06 mcm5p1_cc_w_1_600_s_10_000=1.42e-11 mcm5p1_cf_w_1_600_s_10_000=2.85e-11
+  mcm5p1_ca_w_1_600_s_12_000=8.74e-06 mcm5p1_cc_w_1_600_s_12_000=1.11e-11 mcm5p1_cf_w_1_600_s_12_000=3.11e-11
+  mcm5p1_ca_w_4_000_s_1_600=8.74e-06 mcm5p1_cc_w_4_000_s_1_600=9.42e-11 mcm5p1_cf_w_4_000_s_1_600=6.27e-12
+  mcm5p1_ca_w_4_000_s_1_700=8.74e-06 mcm5p1_cc_w_4_000_s_1_700=8.90e-11 mcm5p1_cf_w_4_000_s_1_700=6.67e-12
+  mcm5p1_ca_w_4_000_s_1_900=8.74e-06 mcm5p1_cc_w_4_000_s_1_900=8.06e-11 mcm5p1_cf_w_4_000_s_1_900=7.46e-12
+  mcm5p1_ca_w_4_000_s_2_000=8.74e-06 mcm5p1_cc_w_4_000_s_2_000=7.70e-11 mcm5p1_cf_w_4_000_s_2_000=7.85e-12
+  mcm5p1_ca_w_4_000_s_2_400=8.74e-06 mcm5p1_cc_w_4_000_s_2_400=6.58e-11 mcm5p1_cf_w_4_000_s_2_400=9.39e-12
+  mcm5p1_ca_w_4_000_s_2_800=8.74e-06 mcm5p1_cc_w_4_000_s_2_800=5.76e-11 mcm5p1_cf_w_4_000_s_2_800=1.09e-11
+  mcm5p1_ca_w_4_000_s_3_200=8.74e-06 mcm5p1_cc_w_4_000_s_3_200=5.14e-11 mcm5p1_cf_w_4_000_s_3_200=1.23e-11
+  mcm5p1_ca_w_4_000_s_4_800=8.74e-06 mcm5p1_cc_w_4_000_s_4_800=3.60e-11 mcm5p1_cf_w_4_000_s_4_800=1.74e-11
+  mcm5p1_ca_w_4_000_s_10_000=8.74e-06 mcm5p1_cc_w_4_000_s_10_000=1.68e-11 mcm5p1_cf_w_4_000_s_10_000=2.90e-11
+  mcm5p1_ca_w_4_000_s_12_000=8.74e-06 mcm5p1_cc_w_4_000_s_12_000=1.34e-11 mcm5p1_cf_w_4_000_s_12_000=3.17e-11
+  mcm5l1_ca_w_1_600_s_1_600=9.48e-06 mcm5l1_cc_w_1_600_s_1_600=8.70e-11 mcm5l1_cf_w_1_600_s_1_600=6.75e-12
+  mcm5l1_ca_w_1_600_s_1_700=9.48e-06 mcm5l1_cc_w_1_600_s_1_700=8.20e-11 mcm5l1_cf_w_1_600_s_1_700=7.18e-12
+  mcm5l1_ca_w_1_600_s_1_900=9.48e-06 mcm5l1_cc_w_1_600_s_1_900=7.36e-11 mcm5l1_cf_w_1_600_s_1_900=8.02e-12
+  mcm5l1_ca_w_1_600_s_2_000=9.48e-06 mcm5l1_cc_w_1_600_s_2_000=7.03e-11 mcm5l1_cf_w_1_600_s_2_000=8.44e-12
+  mcm5l1_ca_w_1_600_s_2_400=9.48e-06 mcm5l1_cc_w_1_600_s_2_400=5.95e-11 mcm5l1_cf_w_1_600_s_2_400=1.01e-11
+  mcm5l1_ca_w_1_600_s_2_800=9.48e-06 mcm5l1_cc_w_1_600_s_2_800=5.17e-11 mcm5l1_cf_w_1_600_s_2_800=1.16e-11
+  mcm5l1_ca_w_1_600_s_3_200=9.48e-06 mcm5l1_cc_w_1_600_s_3_200=4.58e-11 mcm5l1_cf_w_1_600_s_3_200=1.31e-11
+  mcm5l1_ca_w_1_600_s_4_800=9.48e-06 mcm5l1_cc_w_1_600_s_4_800=3.13e-11 mcm5l1_cf_w_1_600_s_4_800=1.86e-11
+  mcm5l1_ca_w_1_600_s_10_000=9.48e-06 mcm5l1_cc_w_1_600_s_10_000=1.35e-11 mcm5l1_cf_w_1_600_s_10_000=3.00e-11
+  mcm5l1_ca_w_1_600_s_12_000=9.48e-06 mcm5l1_cc_w_1_600_s_12_000=1.05e-11 mcm5l1_cf_w_1_600_s_12_000=3.25e-11
+  mcm5l1_ca_w_4_000_s_1_600=9.48e-06 mcm5l1_cc_w_4_000_s_1_600=9.34e-11 mcm5l1_cf_w_4_000_s_1_600=6.76e-12
+  mcm5l1_ca_w_4_000_s_1_700=9.48e-06 mcm5l1_cc_w_4_000_s_1_700=8.82e-11 mcm5l1_cf_w_4_000_s_1_700=7.19e-12
+  mcm5l1_ca_w_4_000_s_1_900=9.48e-06 mcm5l1_cc_w_4_000_s_1_900=7.98e-11 mcm5l1_cf_w_4_000_s_1_900=8.03e-12
+  mcm5l1_ca_w_4_000_s_2_000=9.48e-06 mcm5l1_cc_w_4_000_s_2_000=7.62e-11 mcm5l1_cf_w_4_000_s_2_000=8.45e-12
+  mcm5l1_ca_w_4_000_s_2_400=9.48e-06 mcm5l1_cc_w_4_000_s_2_400=6.49e-11 mcm5l1_cf_w_4_000_s_2_400=1.01e-11
+  mcm5l1_ca_w_4_000_s_2_800=9.48e-06 mcm5l1_cc_w_4_000_s_2_800=5.68e-11 mcm5l1_cf_w_4_000_s_2_800=1.17e-11
+  mcm5l1_ca_w_4_000_s_3_200=9.48e-06 mcm5l1_cc_w_4_000_s_3_200=5.05e-11 mcm5l1_cf_w_4_000_s_3_200=1.32e-11
+  mcm5l1_ca_w_4_000_s_4_800=9.48e-06 mcm5l1_cc_w_4_000_s_4_800=3.52e-11 mcm5l1_cf_w_4_000_s_4_800=1.86e-11
+  mcm5l1_ca_w_4_000_s_10_000=9.48e-06 mcm5l1_cc_w_4_000_s_10_000=1.61e-11 mcm5l1_cf_w_4_000_s_10_000=3.05e-11
+  mcm5l1_ca_w_4_000_s_12_000=9.48e-06 mcm5l1_cc_w_4_000_s_12_000=1.28e-11 mcm5l1_cf_w_4_000_s_12_000=3.32e-11
+  mcm5m1_ca_w_1_600_s_1_600=1.12e-05 mcm5m1_cc_w_1_600_s_1_600=8.53e-11 mcm5m1_cf_w_1_600_s_1_600=7.88e-12
+  mcm5m1_ca_w_1_600_s_1_700=1.12e-05 mcm5m1_cc_w_1_600_s_1_700=8.03e-11 mcm5m1_cf_w_1_600_s_1_700=8.37e-12
+  mcm5m1_ca_w_1_600_s_1_900=1.12e-05 mcm5m1_cc_w_1_600_s_1_900=7.21e-11 mcm5m1_cf_w_1_600_s_1_900=9.34e-12
+  mcm5m1_ca_w_1_600_s_2_000=1.12e-05 mcm5m1_cc_w_1_600_s_2_000=6.87e-11 mcm5m1_cf_w_1_600_s_2_000=9.83e-12
+  mcm5m1_ca_w_1_600_s_2_400=1.12e-05 mcm5m1_cc_w_1_600_s_2_400=5.79e-11 mcm5m1_cf_w_1_600_s_2_400=1.17e-11
+  mcm5m1_ca_w_1_600_s_2_800=1.12e-05 mcm5m1_cc_w_1_600_s_2_800=5.01e-11 mcm5m1_cf_w_1_600_s_2_800=1.35e-11
+  mcm5m1_ca_w_1_600_s_3_200=1.12e-05 mcm5m1_cc_w_1_600_s_3_200=4.42e-11 mcm5m1_cf_w_1_600_s_3_200=1.52e-11
+  mcm5m1_ca_w_1_600_s_4_800=1.12e-05 mcm5m1_cc_w_1_600_s_4_800=2.97e-11 mcm5m1_cf_w_1_600_s_4_800=2.12e-11
+  mcm5m1_ca_w_1_600_s_10_000=1.12e-05 mcm5m1_cc_w_1_600_s_10_000=1.23e-11 mcm5m1_cf_w_1_600_s_10_000=3.31e-11
+  mcm5m1_ca_w_1_600_s_12_000=1.12e-05 mcm5m1_cc_w_1_600_s_12_000=9.39e-12 mcm5m1_cf_w_1_600_s_12_000=3.56e-11
+  mcm5m1_ca_w_4_000_s_1_600=1.12e-05 mcm5m1_cc_w_4_000_s_1_600=9.17e-11 mcm5m1_cf_w_4_000_s_1_600=7.88e-12
+  mcm5m1_ca_w_4_000_s_1_700=1.12e-05 mcm5m1_cc_w_4_000_s_1_700=8.65e-11 mcm5m1_cf_w_4_000_s_1_700=8.37e-12
+  mcm5m1_ca_w_4_000_s_1_900=1.12e-05 mcm5m1_cc_w_4_000_s_1_900=7.81e-11 mcm5m1_cf_w_4_000_s_1_900=9.35e-12
+  mcm5m1_ca_w_4_000_s_2_000=1.12e-05 mcm5m1_cc_w_4_000_s_2_000=7.44e-11 mcm5m1_cf_w_4_000_s_2_000=9.83e-12
+  mcm5m1_ca_w_4_000_s_2_400=1.12e-05 mcm5m1_cc_w_4_000_s_2_400=6.32e-11 mcm5m1_cf_w_4_000_s_2_400=1.17e-11
+  mcm5m1_ca_w_4_000_s_2_800=1.12e-05 mcm5m1_cc_w_4_000_s_2_800=5.51e-11 mcm5m1_cf_w_4_000_s_2_800=1.35e-11
+  mcm5m1_ca_w_4_000_s_3_200=1.12e-05 mcm5m1_cc_w_4_000_s_3_200=4.88e-11 mcm5m1_cf_w_4_000_s_3_200=1.52e-11
+  mcm5m1_ca_w_4_000_s_4_800=1.12e-05 mcm5m1_cc_w_4_000_s_4_800=3.36e-11 mcm5m1_cf_w_4_000_s_4_800=2.13e-11
+  mcm5m1_ca_w_4_000_s_10_000=1.12e-05 mcm5m1_cc_w_4_000_s_10_000=1.49e-11 mcm5m1_cf_w_4_000_s_10_000=3.36e-11
+  mcm5m1_ca_w_4_000_s_12_000=1.12e-05 mcm5m1_cc_w_4_000_s_12_000=1.16e-11 mcm5m1_cf_w_4_000_s_12_000=3.63e-11
+  mcm5m2_ca_w_1_600_s_1_600=1.33e-05 mcm5m2_cc_w_1_600_s_1_600=8.36e-11 mcm5m2_cf_w_1_600_s_1_600=9.30e-12
+  mcm5m2_ca_w_1_600_s_1_700=1.33e-05 mcm5m2_cc_w_1_600_s_1_700=7.85e-11 mcm5m2_cf_w_1_600_s_1_700=9.87e-12
+  mcm5m2_ca_w_1_600_s_1_900=1.33e-05 mcm5m2_cc_w_1_600_s_1_900=7.03e-11 mcm5m2_cf_w_1_600_s_1_900=1.10e-11
+  mcm5m2_ca_w_1_600_s_2_000=1.33e-05 mcm5m2_cc_w_1_600_s_2_000=6.70e-11 mcm5m2_cf_w_1_600_s_2_000=1.16e-11
+  mcm5m2_ca_w_1_600_s_2_400=1.33e-05 mcm5m2_cc_w_1_600_s_2_400=5.61e-11 mcm5m2_cf_w_1_600_s_2_400=1.37e-11
+  mcm5m2_ca_w_1_600_s_2_800=1.33e-05 mcm5m2_cc_w_1_600_s_2_800=4.83e-11 mcm5m2_cf_w_1_600_s_2_800=1.58e-11
+  mcm5m2_ca_w_1_600_s_3_200=1.33e-05 mcm5m2_cc_w_1_600_s_3_200=4.24e-11 mcm5m2_cf_w_1_600_s_3_200=1.77e-11
+  mcm5m2_ca_w_1_600_s_4_800=1.33e-05 mcm5m2_cc_w_1_600_s_4_800=2.79e-11 mcm5m2_cf_w_1_600_s_4_800=2.43e-11
+  mcm5m2_ca_w_1_600_s_10_000=1.33e-05 mcm5m2_cc_w_1_600_s_10_000=1.11e-11 mcm5m2_cf_w_1_600_s_10_000=3.66e-11
+  mcm5m2_ca_w_1_600_s_12_000=1.33e-05 mcm5m2_cc_w_1_600_s_12_000=8.35e-12 mcm5m2_cf_w_1_600_s_12_000=3.90e-11
+  mcm5m2_ca_w_4_000_s_1_600=1.33e-05 mcm5m2_cc_w_4_000_s_1_600=8.98e-11 mcm5m2_cf_w_4_000_s_1_600=9.30e-12
+  mcm5m2_ca_w_4_000_s_1_700=1.33e-05 mcm5m2_cc_w_4_000_s_1_700=8.46e-11 mcm5m2_cf_w_4_000_s_1_700=9.88e-12
+  mcm5m2_ca_w_4_000_s_1_900=1.33e-05 mcm5m2_cc_w_4_000_s_1_900=7.61e-11 mcm5m2_cf_w_4_000_s_1_900=1.10e-11
+  mcm5m2_ca_w_4_000_s_2_000=1.33e-05 mcm5m2_cc_w_4_000_s_2_000=7.26e-11 mcm5m2_cf_w_4_000_s_2_000=1.16e-11
+  mcm5m2_ca_w_4_000_s_2_400=1.33e-05 mcm5m2_cc_w_4_000_s_2_400=6.12e-11 mcm5m2_cf_w_4_000_s_2_400=1.37e-11
+  mcm5m2_ca_w_4_000_s_2_800=1.33e-05 mcm5m2_cc_w_4_000_s_2_800=5.32e-11 mcm5m2_cf_w_4_000_s_2_800=1.58e-11
+  mcm5m2_ca_w_4_000_s_3_200=1.33e-05 mcm5m2_cc_w_4_000_s_3_200=4.70e-11 mcm5m2_cf_w_4_000_s_3_200=1.77e-11
+  mcm5m2_ca_w_4_000_s_4_800=1.33e-05 mcm5m2_cc_w_4_000_s_4_800=3.17e-11 mcm5m2_cf_w_4_000_s_4_800=2.44e-11
+  mcm5m2_ca_w_4_000_s_10_000=1.33e-05 mcm5m2_cc_w_4_000_s_10_000=1.36e-11 mcm5m2_cf_w_4_000_s_10_000=3.72e-11
+  mcm5m2_ca_w_4_000_s_12_000=1.33e-05 mcm5m2_cc_w_4_000_s_12_000=1.06e-11 mcm5m2_cf_w_4_000_s_12_000=3.98e-11
+  mcm5m3_ca_w_1_600_s_1_600=2.46e-05 mcm5m3_cc_w_1_600_s_1_600=7.71e-11 mcm5m3_cf_w_1_600_s_1_600=1.62e-11
+  mcm5m3_ca_w_1_600_s_1_700=2.46e-05 mcm5m3_cc_w_1_600_s_1_700=7.21e-11 mcm5m3_cf_w_1_600_s_1_700=1.72e-11
+  mcm5m3_ca_w_1_600_s_1_900=2.46e-05 mcm5m3_cc_w_1_600_s_1_900=6.41e-11 mcm5m3_cf_w_1_600_s_1_900=1.90e-11
+  mcm5m3_ca_w_1_600_s_2_000=2.46e-05 mcm5m3_cc_w_1_600_s_2_000=6.05e-11 mcm5m3_cf_w_1_600_s_2_000=1.99e-11
+  mcm5m3_ca_w_1_600_s_2_400=2.46e-05 mcm5m3_cc_w_1_600_s_2_400=4.97e-11 mcm5m3_cf_w_1_600_s_2_400=2.32e-11
+  mcm5m3_ca_w_1_600_s_2_800=2.46e-05 mcm5m3_cc_w_1_600_s_2_800=4.20e-11 mcm5m3_cf_w_1_600_s_2_800=2.62e-11
+  mcm5m3_ca_w_1_600_s_3_200=2.46e-05 mcm5m3_cc_w_1_600_s_3_200=3.62e-11 mcm5m3_cf_w_1_600_s_3_200=2.89e-11
+  mcm5m3_ca_w_1_600_s_4_800=2.46e-05 mcm5m3_cc_w_1_600_s_4_800=2.24e-11 mcm5m3_cf_w_1_600_s_4_800=3.74e-11
+  mcm5m3_ca_w_1_600_s_10_000=2.46e-05 mcm5m3_cc_w_1_600_s_10_000=7.70e-12 mcm5m3_cf_w_1_600_s_10_000=4.95e-11
+  mcm5m3_ca_w_1_600_s_12_000=2.46e-05 mcm5m3_cc_w_1_600_s_12_000=5.75e-12 mcm5m3_cf_w_1_600_s_12_000=5.15e-11
+  mcm5m3_ca_w_4_000_s_1_600=2.46e-05 mcm5m3_cc_w_4_000_s_1_600=8.32e-11 mcm5m3_cf_w_4_000_s_1_600=1.62e-11
+  mcm5m3_ca_w_4_000_s_1_700=2.46e-05 mcm5m3_cc_w_4_000_s_1_700=7.80e-11 mcm5m3_cf_w_4_000_s_1_700=1.72e-11
+  mcm5m3_ca_w_4_000_s_1_900=2.46e-05 mcm5m3_cc_w_4_000_s_1_900=6.95e-11 mcm5m3_cf_w_4_000_s_1_900=1.90e-11
+  mcm5m3_ca_w_4_000_s_2_000=2.46e-05 mcm5m3_cc_w_4_000_s_2_000=6.59e-11 mcm5m3_cf_w_4_000_s_2_000=1.99e-11
+  mcm5m3_ca_w_4_000_s_2_400=2.46e-05 mcm5m3_cc_w_4_000_s_2_400=5.47e-11 mcm5m3_cf_w_4_000_s_2_400=2.32e-11
+  mcm5m3_ca_w_4_000_s_2_800=2.46e-05 mcm5m3_cc_w_4_000_s_2_800=4.67e-11 mcm5m3_cf_w_4_000_s_2_800=2.62e-11
+  mcm5m3_ca_w_4_000_s_3_200=2.46e-05 mcm5m3_cc_w_4_000_s_3_200=4.06e-11 mcm5m3_cf_w_4_000_s_3_200=2.90e-11
+  mcm5m3_ca_w_4_000_s_4_800=2.46e-05 mcm5m3_cc_w_4_000_s_4_800=2.61e-11 mcm5m3_cf_w_4_000_s_4_800=3.75e-11
+  mcm5m3_ca_w_4_000_s_10_000=2.46e-05 mcm5m3_cc_w_4_000_s_10_000=1.01e-11 mcm5m3_cf_w_4_000_s_10_000=5.05e-11
+  mcm5m3_ca_w_4_000_s_12_000=2.46e-05 mcm5m3_cc_w_4_000_s_12_000=7.75e-12 mcm5m3_cf_w_4_000_s_12_000=5.28e-11
+  mcm5m4_ca_w_1_600_s_1_600=1.15e-04 mcm5m4_cc_w_1_600_s_1_600=6.12e-11 mcm5m4_cf_w_1_600_s_1_600=5.18e-11
+  mcm5m4_ca_w_1_600_s_1_700=1.15e-04 mcm5m4_cc_w_1_600_s_1_700=5.65e-11 mcm5m4_cf_w_1_600_s_1_700=5.38e-11
+  mcm5m4_ca_w_1_600_s_1_900=1.15e-04 mcm5m4_cc_w_1_600_s_1_900=4.86e-11 mcm5m4_cf_w_1_600_s_1_900=5.73e-11
+  mcm5m4_ca_w_1_600_s_2_000=1.15e-04 mcm5m4_cc_w_1_600_s_2_000=4.54e-11 mcm5m4_cf_w_1_600_s_2_000=5.89e-11
+  mcm5m4_ca_w_1_600_s_2_400=1.15e-04 mcm5m4_cc_w_1_600_s_2_400=3.57e-11 mcm5m4_cf_w_1_600_s_2_400=6.45e-11
+  mcm5m4_ca_w_1_600_s_2_800=1.15e-04 mcm5m4_cc_w_1_600_s_2_800=2.90e-11 mcm5m4_cf_w_1_600_s_2_800=6.89e-11
+  mcm5m4_ca_w_1_600_s_3_200=1.15e-04 mcm5m4_cc_w_1_600_s_3_200=2.42e-11 mcm5m4_cf_w_1_600_s_3_200=7.24e-11
+  mcm5m4_ca_w_1_600_s_4_800=1.15e-04 mcm5m4_cc_w_1_600_s_4_800=1.36e-11 mcm5m4_cf_w_1_600_s_4_800=8.11e-11
+  mcm5m4_ca_w_1_600_s_10_000=1.15e-04 mcm5m4_cc_w_1_600_s_10_000=4.30e-12 mcm5m4_cf_w_1_600_s_10_000=9.00e-11
+  mcm5m4_ca_w_1_600_s_12_000=1.15e-04 mcm5m4_cc_w_1_600_s_12_000=3.15e-12 mcm5m4_cf_w_1_600_s_12_000=9.12e-11
+  mcm5m4_ca_w_4_000_s_1_600=1.15e-04 mcm5m4_cc_w_4_000_s_1_600=6.72e-11 mcm5m4_cf_w_4_000_s_1_600=5.18e-11
+  mcm5m4_ca_w_4_000_s_1_700=1.15e-04 mcm5m4_cc_w_4_000_s_1_700=6.21e-11 mcm5m4_cf_w_4_000_s_1_700=5.38e-11
+  mcm5m4_ca_w_4_000_s_1_900=1.15e-04 mcm5m4_cc_w_4_000_s_1_900=5.42e-11 mcm5m4_cf_w_4_000_s_1_900=5.73e-11
+  mcm5m4_ca_w_4_000_s_2_000=1.15e-04 mcm5m4_cc_w_4_000_s_2_000=5.08e-11 mcm5m4_cf_w_4_000_s_2_000=5.89e-11
+  mcm5m4_ca_w_4_000_s_2_400=1.15e-04 mcm5m4_cc_w_4_000_s_2_400=4.07e-11 mcm5m4_cf_w_4_000_s_2_400=6.45e-11
+  mcm5m4_ca_w_4_000_s_2_800=1.15e-04 mcm5m4_cc_w_4_000_s_2_800=3.38e-11 mcm5m4_cf_w_4_000_s_2_800=6.89e-11
+  mcm5m4_ca_w_4_000_s_3_200=1.15e-04 mcm5m4_cc_w_4_000_s_3_200=2.88e-11 mcm5m4_cf_w_4_000_s_3_200=7.25e-11
+  mcm5m4_ca_w_4_000_s_4_800=1.15e-04 mcm5m4_cc_w_4_000_s_4_800=1.75e-11 mcm5m4_cf_w_4_000_s_4_800=8.16e-11
+  mcm5m4_ca_w_4_000_s_10_000=1.15e-04 mcm5m4_cc_w_4_000_s_10_000=6.45e-12 mcm5m4_cf_w_4_000_s_10_000=9.19e-11
+  mcm5m4_ca_w_4_000_s_12_000=1.15e-04 mcm5m4_cc_w_4_000_s_12_000=4.95e-12 mcm5m4_cf_w_4_000_s_12_000=9.35e-11
+  mcrdlf_ca_w_10_000_s_5_000=3.49e-06 mcrdlf_cc_w_10_000_s_5_000=6.98e-11 mcrdlf_cf_w_10_000_s_5_000=6.48e-12
+  mcrdlf_ca_w_10_000_s_8_000=3.49e-06 mcrdlf_cc_w_10_000_s_8_000=4.70e-11 mcrdlf_cf_w_10_000_s_8_000=1.06e-11
+  mcrdlf_ca_w_10_000_s_10_000=3.49e-06 mcrdlf_cc_w_10_000_s_10_000=3.90e-11 mcrdlf_cf_w_10_000_s_10_000=1.31e-11
+  mcrdlf_ca_w_10_000_s_12_000=3.49e-06 mcrdlf_cc_w_10_000_s_12_000=3.35e-11 mcrdlf_cf_w_10_000_s_12_000=1.53e-11
+  mcrdlf_ca_w_10_000_s_30_000=3.49e-06 mcrdlf_cc_w_10_000_s_30_000=1.37e-11 mcrdlf_cf_w_10_000_s_30_000=2.79e-11
+  mcrdlf_ca_w_40_000_s_5_000=3.49e-06 mcrdlf_cc_w_40_000_s_5_000=8.13e-11 mcrdlf_cf_w_40_000_s_5_000=6.54e-12
+  mcrdlf_ca_w_40_000_s_8_000=3.49e-06 mcrdlf_cc_w_40_000_s_8_000=5.74e-11 mcrdlf_cf_w_40_000_s_8_000=1.07e-11
+  mcrdlf_ca_w_40_000_s_10_000=3.49e-06 mcrdlf_cc_w_40_000_s_10_000=4.89e-11 mcrdlf_cf_w_40_000_s_10_000=1.31e-11
+  mcrdlf_ca_w_40_000_s_12_000=3.49e-06 mcrdlf_cc_w_40_000_s_12_000=4.29e-11 mcrdlf_cf_w_40_000_s_12_000=1.54e-11
+  mcrdlf_ca_w_40_000_s_30_000=3.49e-06 mcrdlf_cc_w_40_000_s_30_000=2.08e-11 mcrdlf_cf_w_40_000_s_30_000=2.85e-11
+  mcrdld_ca_w_10_000_s_5_000=3.57e-06 mcrdld_cc_w_10_000_s_5_000=6.95e-11 mcrdld_cf_w_10_000_s_5_000=6.61e-12
+  mcrdld_ca_w_10_000_s_8_000=3.57e-06 mcrdld_cc_w_10_000_s_8_000=4.68e-11 mcrdld_cf_w_10_000_s_8_000=1.08e-11
+  mcrdld_ca_w_10_000_s_10_000=3.57e-06 mcrdld_cc_w_10_000_s_10_000=3.89e-11 mcrdld_cf_w_10_000_s_10_000=1.33e-11
+  mcrdld_ca_w_10_000_s_12_000=3.57e-06 mcrdld_cc_w_10_000_s_12_000=3.33e-11 mcrdld_cf_w_10_000_s_12_000=1.55e-11
+  mcrdld_ca_w_10_000_s_30_000=3.57e-06 mcrdld_cc_w_10_000_s_30_000=1.35e-11 mcrdld_cf_w_10_000_s_30_000=2.82e-11
+  mcrdld_ca_w_40_000_s_5_000=3.57e-06 mcrdld_cc_w_40_000_s_5_000=8.11e-11 mcrdld_cf_w_40_000_s_5_000=6.67e-12
+  mcrdld_ca_w_40_000_s_8_000=3.57e-06 mcrdld_cc_w_40_000_s_8_000=5.72e-11 mcrdld_cf_w_40_000_s_8_000=1.09e-11
+  mcrdld_ca_w_40_000_s_10_000=3.57e-06 mcrdld_cc_w_40_000_s_10_000=4.88e-11 mcrdld_cf_w_40_000_s_10_000=1.34e-11
+  mcrdld_ca_w_40_000_s_12_000=3.57e-06 mcrdld_cc_w_40_000_s_12_000=4.27e-11 mcrdld_cf_w_40_000_s_12_000=1.56e-11
+  mcrdld_ca_w_40_000_s_30_000=3.57e-06 mcrdld_cc_w_40_000_s_30_000=2.06e-11 mcrdld_cf_w_40_000_s_30_000=2.88e-11
+  mcrdlp1_ca_w_10_000_s_5_000=3.67e-06 mcrdlp1_cc_w_10_000_s_5_000=6.92e-11 mcrdlp1_cf_w_10_000_s_5_000=6.80e-12
+  mcrdlp1_ca_w_10_000_s_8_000=3.67e-06 mcrdlp1_cc_w_10_000_s_8_000=4.65e-11 mcrdlp1_cf_w_10_000_s_8_000=1.11e-11
+  mcrdlp1_ca_w_10_000_s_10_000=3.67e-06 mcrdlp1_cc_w_10_000_s_10_000=3.86e-11 mcrdlp1_cf_w_10_000_s_10_000=1.36e-11
+  mcrdlp1_ca_w_10_000_s_12_000=3.67e-06 mcrdlp1_cc_w_10_000_s_12_000=3.30e-11 mcrdlp1_cf_w_10_000_s_12_000=1.59e-11
+  mcrdlp1_ca_w_10_000_s_30_000=3.67e-06 mcrdlp1_cc_w_10_000_s_30_000=1.33e-11 mcrdlp1_cf_w_10_000_s_30_000=2.86e-11
+  mcrdlp1_ca_w_40_000_s_5_000=3.67e-06 mcrdlp1_cc_w_40_000_s_5_000=8.07e-11 mcrdlp1_cf_w_40_000_s_5_000=6.87e-12
+  mcrdlp1_ca_w_40_000_s_8_000=3.67e-06 mcrdlp1_cc_w_40_000_s_8_000=5.70e-11 mcrdlp1_cf_w_40_000_s_8_000=1.12e-11
+  mcrdlp1_ca_w_40_000_s_10_000=3.67e-06 mcrdlp1_cc_w_40_000_s_10_000=4.84e-11 mcrdlp1_cf_w_40_000_s_10_000=1.37e-11
+  mcrdlp1_ca_w_40_000_s_12_000=3.67e-06 mcrdlp1_cc_w_40_000_s_12_000=4.25e-11 mcrdlp1_cf_w_40_000_s_12_000=1.60e-11
+  mcrdlp1_ca_w_40_000_s_30_000=3.67e-06 mcrdlp1_cc_w_40_000_s_30_000=2.05e-11 mcrdlp1_cf_w_40_000_s_30_000=2.92e-11
+  mcrdll1_ca_w_10_000_s_5_000=3.80e-06 mcrdll1_cc_w_10_000_s_5_000=6.89e-11 mcrdll1_cf_w_10_000_s_5_000=7.00e-12
+  mcrdll1_ca_w_10_000_s_8_000=3.80e-06 mcrdll1_cc_w_10_000_s_8_000=4.62e-11 mcrdll1_cf_w_10_000_s_8_000=1.14e-11
+  mcrdll1_ca_w_10_000_s_10_000=3.80e-06 mcrdll1_cc_w_10_000_s_10_000=3.82e-11 mcrdll1_cf_w_10_000_s_10_000=1.40e-11
+  mcrdll1_ca_w_10_000_s_12_000=3.80e-06 mcrdll1_cc_w_10_000_s_12_000=3.27e-11 mcrdll1_cf_w_10_000_s_12_000=1.63e-11
+  mcrdll1_ca_w_10_000_s_30_000=3.80e-06 mcrdll1_cc_w_10_000_s_30_000=1.31e-11 mcrdll1_cf_w_10_000_s_30_000=2.91e-11
+  mcrdll1_ca_w_40_000_s_5_000=3.80e-06 mcrdll1_cc_w_40_000_s_5_000=8.04e-11 mcrdll1_cf_w_40_000_s_5_000=7.06e-12
+  mcrdll1_ca_w_40_000_s_8_000=3.80e-06 mcrdll1_cc_w_40_000_s_8_000=5.66e-11 mcrdll1_cf_w_40_000_s_8_000=1.15e-11
+  mcrdll1_ca_w_40_000_s_10_000=3.80e-06 mcrdll1_cc_w_40_000_s_10_000=4.81e-11 mcrdll1_cf_w_40_000_s_10_000=1.40e-11
+  mcrdll1_ca_w_40_000_s_12_000=3.80e-06 mcrdll1_cc_w_40_000_s_12_000=4.22e-11 mcrdll1_cf_w_40_000_s_12_000=1.64e-11
+  mcrdll1_ca_w_40_000_s_30_000=3.80e-06 mcrdll1_cc_w_40_000_s_30_000=2.03e-11 mcrdll1_cf_w_40_000_s_30_000=2.97e-11
+  mcrdlm1_ca_w_10_000_s_5_000=4.04e-06 mcrdlm1_cc_w_10_000_s_5_000=6.83e-11 mcrdlm1_cf_w_10_000_s_5_000=7.40e-12
+  mcrdlm1_ca_w_10_000_s_8_000=4.04e-06 mcrdlm1_cc_w_10_000_s_8_000=4.55e-11 mcrdlm1_cf_w_10_000_s_8_000=1.20e-11
+  mcrdlm1_ca_w_10_000_s_10_000=4.04e-06 mcrdlm1_cc_w_10_000_s_10_000=3.77e-11 mcrdlm1_cf_w_10_000_s_10_000=1.47e-11
+  mcrdlm1_ca_w_10_000_s_12_000=4.04e-06 mcrdlm1_cc_w_10_000_s_12_000=3.22e-11 mcrdlm1_cf_w_10_000_s_12_000=1.70e-11
+  mcrdlm1_ca_w_10_000_s_30_000=4.04e-06 mcrdlm1_cc_w_10_000_s_30_000=1.28e-11 mcrdlm1_cf_w_10_000_s_30_000=2.99e-11
+  mcrdlm1_ca_w_40_000_s_5_000=4.04e-06 mcrdlm1_cc_w_40_000_s_5_000=7.98e-11 mcrdlm1_cf_w_40_000_s_5_000=7.44e-12
+  mcrdlm1_ca_w_40_000_s_8_000=4.04e-06 mcrdlm1_cc_w_40_000_s_8_000=5.60e-11 mcrdlm1_cf_w_40_000_s_8_000=1.20e-11
+  mcrdlm1_ca_w_40_000_s_10_000=4.04e-06 mcrdlm1_cc_w_40_000_s_10_000=4.75e-11 mcrdlm1_cf_w_40_000_s_10_000=1.47e-11
+  mcrdlm1_ca_w_40_000_s_12_000=4.04e-06 mcrdlm1_cc_w_40_000_s_12_000=4.16e-11 mcrdlm1_cf_w_40_000_s_12_000=1.71e-11
+  mcrdlm1_ca_w_40_000_s_30_000=4.04e-06 mcrdlm1_cc_w_40_000_s_30_000=1.99e-11 mcrdlm1_cf_w_40_000_s_30_000=3.06e-11
+  mcrdlm2_ca_w_10_000_s_5_000=4.29e-06 mcrdlm2_cc_w_10_000_s_5_000=6.76e-11 mcrdlm2_cf_w_10_000_s_5_000=7.82e-12
+  mcrdlm2_ca_w_10_000_s_8_000=4.29e-06 mcrdlm2_cc_w_10_000_s_8_000=4.49e-11 mcrdlm2_cf_w_10_000_s_8_000=1.26e-11
+  mcrdlm2_ca_w_10_000_s_10_000=4.29e-06 mcrdlm2_cc_w_10_000_s_10_000=3.71e-11 mcrdlm2_cf_w_10_000_s_10_000=1.54e-11
+  mcrdlm2_ca_w_10_000_s_12_000=4.29e-06 mcrdlm2_cc_w_10_000_s_12_000=3.16e-11 mcrdlm2_cf_w_10_000_s_12_000=1.78e-11
+  mcrdlm2_ca_w_10_000_s_30_000=4.29e-06 mcrdlm2_cc_w_10_000_s_30_000=1.24e-11 mcrdlm2_cf_w_10_000_s_30_000=3.08e-11
+  mcrdlm2_ca_w_40_000_s_5_000=4.29e-06 mcrdlm2_cc_w_40_000_s_5_000=7.91e-11 mcrdlm2_cf_w_40_000_s_5_000=7.86e-12
+  mcrdlm2_ca_w_40_000_s_8_000=4.29e-06 mcrdlm2_cc_w_40_000_s_8_000=5.54e-11 mcrdlm2_cf_w_40_000_s_8_000=1.27e-11
+  mcrdlm2_ca_w_40_000_s_10_000=4.29e-06 mcrdlm2_cc_w_40_000_s_10_000=4.70e-11 mcrdlm2_cf_w_40_000_s_10_000=1.54e-11
+  mcrdlm2_ca_w_40_000_s_12_000=4.29e-06 mcrdlm2_cc_w_40_000_s_12_000=4.11e-11 mcrdlm2_cf_w_40_000_s_12_000=1.79e-11
+  mcrdlm2_ca_w_40_000_s_30_000=4.29e-06 mcrdlm2_cc_w_40_000_s_30_000=1.96e-11 mcrdlm2_cf_w_40_000_s_30_000=3.15e-11
+  mcrdlm3_ca_w_10_000_s_5_000=5.04e-06 mcrdlm3_cc_w_10_000_s_5_000=6.60e-11 mcrdlm3_cf_w_10_000_s_5_000=9.01e-12
+  mcrdlm3_ca_w_10_000_s_8_000=5.04e-06 mcrdlm3_cc_w_10_000_s_8_000=4.34e-11 mcrdlm3_cf_w_10_000_s_8_000=1.43e-11
+  mcrdlm3_ca_w_10_000_s_10_000=5.04e-06 mcrdlm3_cc_w_10_000_s_10_000=3.57e-11 mcrdlm3_cf_w_10_000_s_10_000=1.73e-11
+  mcrdlm3_ca_w_10_000_s_12_000=5.04e-06 mcrdlm3_cc_w_10_000_s_12_000=3.03e-11 mcrdlm3_cf_w_10_000_s_12_000=1.99e-11
+  mcrdlm3_ca_w_10_000_s_30_000=5.04e-06 mcrdlm3_cc_w_10_000_s_30_000=1.17e-11 mcrdlm3_cf_w_10_000_s_30_000=3.31e-11
+  mcrdlm3_ca_w_40_000_s_5_000=5.04e-06 mcrdlm3_cc_w_40_000_s_5_000=7.76e-11 mcrdlm3_cf_w_40_000_s_5_000=9.02e-12
+  mcrdlm3_ca_w_40_000_s_8_000=5.04e-06 mcrdlm3_cc_w_40_000_s_8_000=5.39e-11 mcrdlm3_cf_w_40_000_s_8_000=1.44e-11
+  mcrdlm3_ca_w_40_000_s_10_000=5.04e-06 mcrdlm3_cc_w_40_000_s_10_000=4.56e-11 mcrdlm3_cf_w_40_000_s_10_000=1.74e-11
+  mcrdlm3_ca_w_40_000_s_12_000=5.04e-06 mcrdlm3_cc_w_40_000_s_12_000=3.98e-11 mcrdlm3_cf_w_40_000_s_12_000=2.00e-11
+  mcrdlm3_ca_w_40_000_s_30_000=5.04e-06 mcrdlm3_cc_w_40_000_s_30_000=1.88e-11 mcrdlm3_cf_w_40_000_s_30_000=3.40e-11
+  mcrdlm4_ca_w_10_000_s_5_000=6.01e-06 mcrdlm4_cc_w_10_000_s_5_000=6.43e-11 mcrdlm4_cf_w_10_000_s_5_000=1.05e-11
+  mcrdlm4_ca_w_10_000_s_8_000=6.01e-06 mcrdlm4_cc_w_10_000_s_8_000=4.19e-11 mcrdlm4_cf_w_10_000_s_8_000=1.64e-11
+  mcrdlm4_ca_w_10_000_s_10_000=6.01e-06 mcrdlm4_cc_w_10_000_s_10_000=3.42e-11 mcrdlm4_cf_w_10_000_s_10_000=1.96e-11
+  mcrdlm4_ca_w_10_000_s_12_000=6.01e-06 mcrdlm4_cc_w_10_000_s_12_000=2.89e-11 mcrdlm4_cf_w_10_000_s_12_000=2.24e-11
+  mcrdlm4_ca_w_10_000_s_30_000=6.01e-06 mcrdlm4_cc_w_10_000_s_30_000=1.09e-11 mcrdlm4_cf_w_10_000_s_30_000=3.56e-11
+  mcrdlm4_ca_w_40_000_s_5_000=6.01e-06 mcrdlm4_cc_w_40_000_s_5_000=7.59e-11 mcrdlm4_cf_w_40_000_s_5_000=1.04e-11
+  mcrdlm4_ca_w_40_000_s_8_000=6.01e-06 mcrdlm4_cc_w_40_000_s_8_000=5.23e-11 mcrdlm4_cf_w_40_000_s_8_000=1.64e-11
+  mcrdlm4_ca_w_40_000_s_10_000=6.01e-06 mcrdlm4_cc_w_40_000_s_10_000=4.41e-11 mcrdlm4_cf_w_40_000_s_10_000=1.96e-11
+  mcrdlm4_ca_w_40_000_s_12_000=6.01e-06 mcrdlm4_cc_w_40_000_s_12_000=3.85e-11 mcrdlm4_cf_w_40_000_s_12_000=2.24e-11
+  mcrdlm4_ca_w_40_000_s_30_000=6.01e-06 mcrdlm4_cc_w_40_000_s_30_000=1.80e-11 mcrdlm4_cf_w_40_000_s_30_000=3.66e-11
+  mcrdlm5_ca_w_10_000_s_5_000=8.81e-06 mcrdlm5_cc_w_10_000_s_5_000=6.08e-11 mcrdlm5_cf_w_10_000_s_5_000=1.43e-11
+  mcrdlm5_ca_w_10_000_s_8_000=8.81e-06 mcrdlm5_cc_w_10_000_s_8_000=3.88e-11 mcrdlm5_cf_w_10_000_s_8_000=2.15e-11
+  mcrdlm5_ca_w_10_000_s_10_000=8.81e-06 mcrdlm5_cc_w_10_000_s_10_000=3.14e-11 mcrdlm5_cf_w_10_000_s_10_000=2.51e-11
+  mcrdlm5_ca_w_10_000_s_12_000=8.81e-06 mcrdlm5_cc_w_10_000_s_12_000=2.64e-11 mcrdlm5_cf_w_10_000_s_12_000=2.81e-11
+  mcrdlm5_ca_w_10_000_s_30_000=8.81e-06 mcrdlm5_cc_w_10_000_s_30_000=9.60e-12 mcrdlm5_cf_w_10_000_s_30_000=4.13e-11
+  mcrdlm5_ca_w_40_000_s_5_000=8.81e-06 mcrdlm5_cc_w_40_000_s_5_000=7.24e-11 mcrdlm5_cf_w_40_000_s_5_000=1.42e-11
+  mcrdlm5_ca_w_40_000_s_8_000=8.81e-06 mcrdlm5_cc_w_40_000_s_8_000=4.93e-11 mcrdlm5_cf_w_40_000_s_8_000=2.15e-11
+  mcrdlm5_ca_w_40_000_s_10_000=8.81e-06 mcrdlm5_cc_w_40_000_s_10_000=4.14e-11 mcrdlm5_cf_w_40_000_s_10_000=2.51e-11
+  mcrdlm5_ca_w_40_000_s_12_000=8.81e-06 mcrdlm5_cc_w_40_000_s_12_000=3.59e-11 mcrdlm5_cf_w_40_000_s_12_000=2.81e-11
+  mcrdlm5_ca_w_40_000_s_30_000=8.81e-06 mcrdlm5_cc_w_40_000_s_30_000=1.67e-11 mcrdlm5_cf_w_40_000_s_30_000=4.25e-11
+  mcl1p1f_ca_w_0_150_s_0_210=3.29e-04 mcl1p1f_cc_w_0_150_s_0_210=6.99e-11 mcl1p1f_cf_w_0_150_s_0_210=2.72e-11
+  mcl1p1f_ca_w_0_150_s_0_263=3.29e-04 mcl1p1f_cc_w_0_150_s_0_263=4.97e-11 mcl1p1f_cf_w_0_150_s_0_263=3.31e-11
+  mcl1p1f_ca_w_0_150_s_0_315=3.29e-04 mcl1p1f_cc_w_0_150_s_0_315=3.70e-11 mcl1p1f_cf_w_0_150_s_0_315=3.82e-11
+  mcl1p1f_ca_w_0_150_s_0_420=3.29e-04 mcl1p1f_cc_w_0_150_s_0_420=2.18e-11 mcl1p1f_cf_w_0_150_s_0_420=4.66e-11
+  mcl1p1f_ca_w_0_150_s_0_525=3.29e-04 mcl1p1f_cc_w_0_150_s_0_525=1.33e-11 mcl1p1f_cf_w_0_150_s_0_525=5.27e-11
+  mcl1p1f_ca_w_0_150_s_0_630=3.29e-04 mcl1p1f_cc_w_0_150_s_0_630=8.23e-12 mcl1p1f_cf_w_0_150_s_0_630=5.66e-11
+  mcl1p1f_ca_w_0_150_s_0_840=3.29e-04 mcl1p1f_cc_w_0_150_s_0_840=3.19e-12 mcl1p1f_cf_w_0_150_s_0_840=6.13e-11
+  mcl1p1f_ca_w_0_150_s_1_260=3.29e-04 mcl1p1f_cc_w_0_150_s_1_260=6.20e-13 mcl1p1f_cf_w_0_150_s_1_260=6.37e-11
+  mcl1p1f_ca_w_0_150_s_2_310=3.29e-04 mcl1p1f_cc_w_0_150_s_2_310=5.00e-14 mcl1p1f_cf_w_0_150_s_2_310=6.42e-11
+  mcl1p1f_ca_w_0_150_s_5_250=3.29e-04 mcl1p1f_cc_w_0_150_s_5_250=2.50e-14 mcl1p1f_cf_w_0_150_s_5_250=6.43e-11
+  mcl1p1f_ca_w_1_200_s_0_210=3.29e-04 mcl1p1f_cc_w_1_200_s_0_210=7.07e-11 mcl1p1f_cf_w_1_200_s_0_210=2.70e-11
+  mcl1p1f_ca_w_1_200_s_0_263=3.29e-04 mcl1p1f_cc_w_1_200_s_0_263=5.01e-11 mcl1p1f_cf_w_1_200_s_0_263=3.28e-11
+  mcl1p1f_ca_w_1_200_s_0_315=3.29e-04 mcl1p1f_cc_w_1_200_s_0_315=3.75e-11 mcl1p1f_cf_w_1_200_s_0_315=3.80e-11
+  mcl1p1f_ca_w_1_200_s_0_420=3.29e-04 mcl1p1f_cc_w_1_200_s_0_420=2.21e-11 mcl1p1f_cf_w_1_200_s_0_420=4.64e-11
+  mcl1p1f_ca_w_1_200_s_0_525=3.29e-04 mcl1p1f_cc_w_1_200_s_0_525=1.35e-11 mcl1p1f_cf_w_1_200_s_0_525=5.25e-11
+  mcl1p1f_ca_w_1_200_s_0_630=3.29e-04 mcl1p1f_cc_w_1_200_s_0_630=8.35e-12 mcl1p1f_cf_w_1_200_s_0_630=5.67e-11
+  mcl1p1f_ca_w_1_200_s_0_840=3.29e-04 mcl1p1f_cc_w_1_200_s_0_840=3.25e-12 mcl1p1f_cf_w_1_200_s_0_840=6.12e-11
+  mcl1p1f_ca_w_1_200_s_1_260=3.29e-04 mcl1p1f_cc_w_1_200_s_1_260=5.50e-13 mcl1p1f_cf_w_1_200_s_1_260=6.39e-11
+  mcl1p1f_ca_w_1_200_s_2_310=3.29e-04 mcl1p1f_cc_w_1_200_s_2_310=5.00e-14 mcl1p1f_cf_w_1_200_s_2_310=6.44e-11
+  mcl1p1f_ca_w_1_200_s_5_250=3.29e-04 mcl1p1f_cc_w_1_200_s_5_250=0.00e+00 mcl1p1f_cf_w_1_200_s_5_250=6.44e-11
+  mcm1p1f_ca_w_0_150_s_0_210=2.29e-04 mcm1p1f_cc_w_0_150_s_0_210=7.90e-11 mcm1p1f_cf_w_0_150_s_0_210=1.98e-11
+  mcm1p1f_ca_w_0_150_s_0_263=2.29e-04 mcm1p1f_cc_w_0_150_s_0_263=5.87e-11 mcm1p1f_cf_w_0_150_s_0_263=2.43e-11
+  mcm1p1f_ca_w_0_150_s_0_315=2.29e-04 mcm1p1f_cc_w_0_150_s_0_315=4.58e-11 mcm1p1f_cf_w_0_150_s_0_315=2.85e-11
+  mcm1p1f_ca_w_0_150_s_0_420=2.29e-04 mcm1p1f_cc_w_0_150_s_0_420=3.00e-11 mcm1p1f_cf_w_0_150_s_0_420=3.57e-11
+  mcm1p1f_ca_w_0_150_s_0_525=2.29e-04 mcm1p1f_cc_w_0_150_s_0_525=2.05e-11 mcm1p1f_cf_w_0_150_s_0_525=4.14e-11
+  mcm1p1f_ca_w_0_150_s_0_630=2.29e-04 mcm1p1f_cc_w_0_150_s_0_630=1.43e-11 mcm1p1f_cf_w_0_150_s_0_630=4.57e-11
+  mcm1p1f_ca_w_0_150_s_0_840=2.29e-04 mcm1p1f_cc_w_0_150_s_0_840=7.29e-12 mcm1p1f_cf_w_0_150_s_0_840=5.15e-11
+  mcm1p1f_ca_w_0_150_s_1_260=2.29e-04 mcm1p1f_cc_w_0_150_s_1_260=2.00e-12 mcm1p1f_cf_w_0_150_s_1_260=5.64e-11
+  mcm1p1f_ca_w_0_150_s_2_310=2.29e-04 mcm1p1f_cc_w_0_150_s_2_310=1.15e-13 mcm1p1f_cf_w_0_150_s_2_310=5.82e-11
+  mcm1p1f_ca_w_0_150_s_5_250=2.29e-04 mcm1p1f_cc_w_0_150_s_5_250=0.00e+00 mcm1p1f_cf_w_0_150_s_5_250=5.84e-11
+  mcm1p1f_ca_w_1_200_s_0_210=2.29e-04 mcm1p1f_cc_w_1_200_s_0_210=8.24e-11 mcm1p1f_cf_w_1_200_s_0_210=1.96e-11
+  mcm1p1f_ca_w_1_200_s_0_263=2.29e-04 mcm1p1f_cc_w_1_200_s_0_263=6.13e-11 mcm1p1f_cf_w_1_200_s_0_263=2.42e-11
+  mcm1p1f_ca_w_1_200_s_0_315=2.29e-04 mcm1p1f_cc_w_1_200_s_0_315=4.80e-11 mcm1p1f_cf_w_1_200_s_0_315=2.83e-11
+  mcm1p1f_ca_w_1_200_s_0_420=2.29e-04 mcm1p1f_cc_w_1_200_s_0_420=3.16e-11 mcm1p1f_cf_w_1_200_s_0_420=3.56e-11
+  mcm1p1f_ca_w_1_200_s_0_525=2.29e-04 mcm1p1f_cc_w_1_200_s_0_525=2.18e-11 mcm1p1f_cf_w_1_200_s_0_525=4.14e-11
+  mcm1p1f_ca_w_1_200_s_0_630=2.29e-04 mcm1p1f_cc_w_1_200_s_0_630=1.54e-11 mcm1p1f_cf_w_1_200_s_0_630=4.59e-11
+  mcm1p1f_ca_w_1_200_s_0_840=2.29e-04 mcm1p1f_cc_w_1_200_s_0_840=7.90e-12 mcm1p1f_cf_w_1_200_s_0_840=5.20e-11
+  mcm1p1f_ca_w_1_200_s_1_260=2.29e-04 mcm1p1f_cc_w_1_200_s_1_260=2.20e-12 mcm1p1f_cf_w_1_200_s_1_260=5.72e-11
+  mcm1p1f_ca_w_1_200_s_2_310=2.29e-04 mcm1p1f_cc_w_1_200_s_2_310=1.50e-13 mcm1p1f_cf_w_1_200_s_2_310=5.92e-11
+  mcm1p1f_ca_w_1_200_s_5_250=2.29e-04 mcm1p1f_cc_w_1_200_s_5_250=5.00e-14 mcm1p1f_cf_w_1_200_s_5_250=5.94e-11
+  mcm2p1f_ca_w_0_150_s_0_210=1.91e-04 mcm2p1f_cc_w_0_150_s_0_210=8.41e-11 mcm2p1f_cf_w_0_150_s_0_210=1.66e-11
+  mcm2p1f_ca_w_0_150_s_0_263=1.91e-04 mcm2p1f_cc_w_0_150_s_0_263=6.40e-11 mcm2p1f_cf_w_0_150_s_0_263=2.04e-11
+  mcm2p1f_ca_w_0_150_s_0_315=1.91e-04 mcm2p1f_cc_w_0_150_s_0_315=5.13e-11 mcm2p1f_cf_w_0_150_s_0_315=2.39e-11
+  mcm2p1f_ca_w_0_150_s_0_420=1.91e-04 mcm2p1f_cc_w_0_150_s_0_420=3.58e-11 mcm2p1f_cf_w_0_150_s_0_420=3.02e-11
+  mcm2p1f_ca_w_0_150_s_0_525=1.91e-04 mcm2p1f_cc_w_0_150_s_0_525=2.62e-11 mcm2p1f_cf_w_0_150_s_0_525=3.53e-11
+  mcm2p1f_ca_w_0_150_s_0_630=1.91e-04 mcm2p1f_cc_w_0_150_s_0_630=1.97e-11 mcm2p1f_cf_w_0_150_s_0_630=3.94e-11
+  mcm2p1f_ca_w_0_150_s_0_840=1.91e-04 mcm2p1f_cc_w_0_150_s_0_840=1.19e-11 mcm2p1f_cf_w_0_150_s_0_840=4.54e-11
+  mcm2p1f_ca_w_0_150_s_1_260=1.91e-04 mcm2p1f_cc_w_0_150_s_1_260=4.69e-12 mcm2p1f_cf_w_0_150_s_1_260=5.15e-11
+  mcm2p1f_ca_w_0_150_s_2_310=1.91e-04 mcm2p1f_cc_w_0_150_s_2_310=5.60e-13 mcm2p1f_cf_w_0_150_s_2_310=5.54e-11
+  mcm2p1f_ca_w_0_150_s_5_250=1.91e-04 mcm2p1f_cc_w_0_150_s_5_250=0.00e+00 mcm2p1f_cf_w_0_150_s_5_250=5.60e-11
+  mcm2p1f_ca_w_1_200_s_0_210=1.91e-04 mcm2p1f_cc_w_1_200_s_0_210=9.14e-11 mcm2p1f_cf_w_1_200_s_0_210=1.64e-11
+  mcm2p1f_ca_w_1_200_s_0_263=1.91e-04 mcm2p1f_cc_w_1_200_s_0_263=7.02e-11 mcm2p1f_cf_w_1_200_s_0_263=2.04e-11
+  mcm2p1f_ca_w_1_200_s_0_315=1.91e-04 mcm2p1f_cc_w_1_200_s_0_315=5.69e-11 mcm2p1f_cf_w_1_200_s_0_315=2.39e-11
+  mcm2p1f_ca_w_1_200_s_0_420=1.91e-04 mcm2p1f_cc_w_1_200_s_0_420=4.00e-11 mcm2p1f_cf_w_1_200_s_0_420=3.02e-11
+  mcm2p1f_ca_w_1_200_s_0_525=1.91e-04 mcm2p1f_cc_w_1_200_s_0_525=2.98e-11 mcm2p1f_cf_w_1_200_s_0_525=3.54e-11
+  mcm2p1f_ca_w_1_200_s_0_630=1.91e-04 mcm2p1f_cc_w_1_200_s_0_630=2.28e-11 mcm2p1f_cf_w_1_200_s_0_630=3.97e-11
+  mcm2p1f_ca_w_1_200_s_0_840=1.91e-04 mcm2p1f_cc_w_1_200_s_0_840=1.40e-11 mcm2p1f_cf_w_1_200_s_0_840=4.61e-11
+  mcm2p1f_ca_w_1_200_s_1_260=1.91e-04 mcm2p1f_cc_w_1_200_s_1_260=5.78e-12 mcm2p1f_cf_w_1_200_s_1_260=5.31e-11
+  mcm2p1f_ca_w_1_200_s_2_310=1.91e-04 mcm2p1f_cc_w_1_200_s_2_310=7.10e-13 mcm2p1f_cf_w_1_200_s_2_310=5.78e-11
+  mcm2p1f_ca_w_1_200_s_5_250=1.91e-04 mcm2p1f_cc_w_1_200_s_5_250=0.00e+00 mcm2p1f_cf_w_1_200_s_5_250=5.86e-11
+  mcm3p1f_ca_w_0_150_s_0_210=1.76e-04 mcm3p1f_cc_w_0_150_s_0_210=8.60e-11 mcm3p1f_cf_w_0_150_s_0_210=1.53e-11
+  mcm3p1f_ca_w_0_150_s_0_263=1.76e-04 mcm3p1f_cc_w_0_150_s_0_263=6.62e-11 mcm3p1f_cf_w_0_150_s_0_263=1.88e-11
+  mcm3p1f_ca_w_0_150_s_0_315=1.76e-04 mcm3p1f_cc_w_0_150_s_0_315=5.39e-11 mcm3p1f_cf_w_0_150_s_0_315=2.20e-11
+  mcm3p1f_ca_w_0_150_s_0_420=1.76e-04 mcm3p1f_cc_w_0_150_s_0_420=3.85e-11 mcm3p1f_cf_w_0_150_s_0_420=2.79e-11
+  mcm3p1f_ca_w_0_150_s_0_525=1.76e-04 mcm3p1f_cc_w_0_150_s_0_525=2.92e-11 mcm3p1f_cf_w_0_150_s_0_525=3.26e-11
+  mcm3p1f_ca_w_0_150_s_0_630=1.76e-04 mcm3p1f_cc_w_0_150_s_0_630=2.27e-11 mcm3p1f_cf_w_0_150_s_0_630=3.65e-11
+  mcm3p1f_ca_w_0_150_s_0_840=1.76e-04 mcm3p1f_cc_w_0_150_s_0_840=1.46e-11 mcm3p1f_cf_w_0_150_s_0_840=4.24e-11
+  mcm3p1f_ca_w_0_150_s_1_260=1.76e-04 mcm3p1f_cc_w_0_150_s_1_260=6.70e-12 mcm3p1f_cf_w_0_150_s_1_260=4.90e-11
+  mcm3p1f_ca_w_0_150_s_2_310=1.76e-04 mcm3p1f_cc_w_0_150_s_2_310=1.33e-12 mcm3p1f_cf_w_0_150_s_2_310=5.39e-11
+  mcm3p1f_ca_w_0_150_s_5_250=1.76e-04 mcm3p1f_cc_w_0_150_s_5_250=7.50e-14 mcm3p1f_cf_w_0_150_s_5_250=5.52e-11
+  mcm3p1f_ca_w_1_200_s_0_210=1.76e-04 mcm3p1f_cc_w_1_200_s_0_210=9.66e-11 mcm3p1f_cf_w_1_200_s_0_210=1.52e-11
+  mcm3p1f_ca_w_1_200_s_0_263=1.76e-04 mcm3p1f_cc_w_1_200_s_0_263=7.55e-11 mcm3p1f_cf_w_1_200_s_0_263=1.88e-11
+  mcm3p1f_ca_w_1_200_s_0_315=1.76e-04 mcm3p1f_cc_w_1_200_s_0_315=6.22e-11 mcm3p1f_cf_w_1_200_s_0_315=2.20e-11
+  mcm3p1f_ca_w_1_200_s_0_420=1.76e-04 mcm3p1f_cc_w_1_200_s_0_420=4.54e-11 mcm3p1f_cf_w_1_200_s_0_420=2.78e-11
+  mcm3p1f_ca_w_1_200_s_0_525=1.76e-04 mcm3p1f_cc_w_1_200_s_0_525=3.50e-11 mcm3p1f_cf_w_1_200_s_0_525=3.27e-11
+  mcm3p1f_ca_w_1_200_s_0_630=1.76e-04 mcm3p1f_cc_w_1_200_s_0_630=2.78e-11 mcm3p1f_cf_w_1_200_s_0_630=3.68e-11
+  mcm3p1f_ca_w_1_200_s_0_840=1.76e-04 mcm3p1f_cc_w_1_200_s_0_840=1.86e-11 mcm3p1f_cf_w_1_200_s_0_840=4.31e-11
+  mcm3p1f_ca_w_1_200_s_1_260=1.76e-04 mcm3p1f_cc_w_1_200_s_1_260=9.21e-12 mcm3p1f_cf_w_1_200_s_1_260=5.06e-11
+  mcm3p1f_ca_w_1_200_s_2_310=1.76e-04 mcm3p1f_cc_w_1_200_s_2_310=1.92e-12 mcm3p1f_cf_w_1_200_s_2_310=5.73e-11
+  mcm3p1f_ca_w_1_200_s_5_250=1.76e-04 mcm3p1f_cc_w_1_200_s_5_250=7.50e-14 mcm3p1f_cf_w_1_200_s_5_250=5.92e-11
+  mcm4p1f_ca_w_0_150_s_0_210=1.67e-04 mcm4p1f_cc_w_0_150_s_0_210=8.73e-11 mcm4p1f_cf_w_0_150_s_0_210=1.45e-11
+  mcm4p1f_ca_w_0_150_s_0_263=1.67e-04 mcm4p1f_cc_w_0_150_s_0_263=6.76e-11 mcm4p1f_cf_w_0_150_s_0_263=1.78e-11
+  mcm4p1f_ca_w_0_150_s_0_315=1.67e-04 mcm4p1f_cc_w_0_150_s_0_315=5.55e-11 mcm4p1f_cf_w_0_150_s_0_315=2.09e-11
+  mcm4p1f_ca_w_0_150_s_0_420=1.67e-04 mcm4p1f_cc_w_0_150_s_0_420=4.03e-11 mcm4p1f_cf_w_0_150_s_0_420=2.64e-11
+  mcm4p1f_ca_w_0_150_s_0_525=1.67e-04 mcm4p1f_cc_w_0_150_s_0_525=3.11e-11 mcm4p1f_cf_w_0_150_s_0_525=3.09e-11
+  mcm4p1f_ca_w_0_150_s_0_630=1.67e-04 mcm4p1f_cc_w_0_150_s_0_630=2.48e-11 mcm4p1f_cf_w_0_150_s_0_630=3.46e-11
+  mcm4p1f_ca_w_0_150_s_0_840=1.67e-04 mcm4p1f_cc_w_0_150_s_0_840=1.67e-11 mcm4p1f_cf_w_0_150_s_0_840=4.04e-11
+  mcm4p1f_ca_w_0_150_s_1_260=1.67e-04 mcm4p1f_cc_w_0_150_s_1_260=8.46e-12 mcm4p1f_cf_w_0_150_s_1_260=4.73e-11
+  mcm4p1f_ca_w_0_150_s_2_310=1.67e-04 mcm4p1f_cc_w_0_150_s_2_310=2.23e-12 mcm4p1f_cf_w_0_150_s_2_310=5.29e-11
+  mcm4p1f_ca_w_0_150_s_5_250=1.67e-04 mcm4p1f_cc_w_0_150_s_5_250=1.60e-13 mcm4p1f_cf_w_0_150_s_5_250=5.49e-11
+  mcm4p1f_ca_w_1_200_s_0_210=1.67e-04 mcm4p1f_cc_w_1_200_s_0_210=1.01e-10 mcm4p1f_cf_w_1_200_s_0_210=1.45e-11
+  mcm4p1f_ca_w_1_200_s_0_263=1.67e-04 mcm4p1f_cc_w_1_200_s_0_263=7.96e-11 mcm4p1f_cf_w_1_200_s_0_263=1.78e-11
+  mcm4p1f_ca_w_1_200_s_0_315=1.67e-04 mcm4p1f_cc_w_1_200_s_0_315=6.64e-11 mcm4p1f_cf_w_1_200_s_0_315=2.09e-11
+  mcm4p1f_ca_w_1_200_s_0_420=1.67e-04 mcm4p1f_cc_w_1_200_s_0_420=4.96e-11 mcm4p1f_cf_w_1_200_s_0_420=2.63e-11
+  mcm4p1f_ca_w_1_200_s_0_525=1.67e-04 mcm4p1f_cc_w_1_200_s_0_525=3.93e-11 mcm4p1f_cf_w_1_200_s_0_525=3.10e-11
+  mcm4p1f_ca_w_1_200_s_0_630=1.67e-04 mcm4p1f_cc_w_1_200_s_0_630=3.21e-11 mcm4p1f_cf_w_1_200_s_0_630=3.49e-11
+  mcm4p1f_ca_w_1_200_s_0_840=1.67e-04 mcm4p1f_cc_w_1_200_s_0_840=2.27e-11 mcm4p1f_cf_w_1_200_s_0_840=4.10e-11
+  mcm4p1f_ca_w_1_200_s_1_260=1.67e-04 mcm4p1f_cc_w_1_200_s_1_260=1.27e-11 mcm4p1f_cf_w_1_200_s_1_260=4.88e-11
+  mcm4p1f_ca_w_1_200_s_2_310=1.67e-04 mcm4p1f_cc_w_1_200_s_2_310=3.78e-12 mcm4p1f_cf_w_1_200_s_2_310=5.68e-11
+  mcm4p1f_ca_w_1_200_s_5_250=1.67e-04 mcm4p1f_cc_w_1_200_s_5_250=2.40e-13 mcm4p1f_cf_w_1_200_s_5_250=6.03e-11
+  mcm5p1f_ca_w_0_150_s_0_210=1.64e-04 mcm5p1f_cc_w_0_150_s_0_210=8.78e-11 mcm5p1f_cf_w_0_150_s_0_210=1.42e-11
+  mcm5p1f_ca_w_0_150_s_0_263=1.64e-04 mcm5p1f_cc_w_0_150_s_0_263=6.82e-11 mcm5p1f_cf_w_0_150_s_0_263=1.74e-11
+  mcm5p1f_ca_w_0_150_s_0_315=1.64e-04 mcm5p1f_cc_w_0_150_s_0_315=5.62e-11 mcm5p1f_cf_w_0_150_s_0_315=2.03e-11
+  mcm5p1f_ca_w_0_150_s_0_420=1.64e-04 mcm5p1f_cc_w_0_150_s_0_420=4.11e-11 mcm5p1f_cf_w_0_150_s_0_420=2.57e-11
+  mcm5p1f_ca_w_0_150_s_0_525=1.64e-04 mcm5p1f_cc_w_0_150_s_0_525=3.21e-11 mcm5p1f_cf_w_0_150_s_0_525=3.01e-11
+  mcm5p1f_ca_w_0_150_s_0_630=1.64e-04 mcm5p1f_cc_w_0_150_s_0_630=2.59e-11 mcm5p1f_cf_w_0_150_s_0_630=3.37e-11
+  mcm5p1f_ca_w_0_150_s_0_840=1.64e-04 mcm5p1f_cc_w_0_150_s_0_840=1.78e-11 mcm5p1f_cf_w_0_150_s_0_840=3.94e-11
+  mcm5p1f_ca_w_0_150_s_1_260=1.64e-04 mcm5p1f_cc_w_0_150_s_1_260=9.36e-12 mcm5p1f_cf_w_0_150_s_1_260=4.65e-11
+  mcm5p1f_ca_w_0_150_s_2_310=1.64e-04 mcm5p1f_cc_w_0_150_s_2_310=2.86e-12 mcm5p1f_cf_w_0_150_s_2_310=5.23e-11
+  mcm5p1f_ca_w_0_150_s_5_250=1.64e-04 mcm5p1f_cc_w_0_150_s_5_250=2.66e-13 mcm5p1f_cf_w_0_150_s_5_250=5.48e-11
+  mcm5p1f_ca_w_1_200_s_0_210=1.64e-04 mcm5p1f_cc_w_1_200_s_0_210=1.03e-10 mcm5p1f_cf_w_1_200_s_0_210=1.41e-11
+  mcm5p1f_ca_w_1_200_s_0_263=1.64e-04 mcm5p1f_cc_w_1_200_s_0_263=8.18e-11 mcm5p1f_cf_w_1_200_s_0_263=1.74e-11
+  mcm5p1f_ca_w_1_200_s_0_315=1.64e-04 mcm5p1f_cc_w_1_200_s_0_315=6.87e-11 mcm5p1f_cf_w_1_200_s_0_315=2.03e-11
+  mcm5p1f_ca_w_1_200_s_0_420=1.64e-04 mcm5p1f_cc_w_1_200_s_0_420=5.20e-11 mcm5p1f_cf_w_1_200_s_0_420=2.56e-11
+  mcm5p1f_ca_w_1_200_s_0_525=1.64e-04 mcm5p1f_cc_w_1_200_s_0_525=4.17e-11 mcm5p1f_cf_w_1_200_s_0_525=3.02e-11
+  mcm5p1f_ca_w_1_200_s_0_630=1.64e-04 mcm5p1f_cc_w_1_200_s_0_630=3.46e-11 mcm5p1f_cf_w_1_200_s_0_630=3.40e-11
+  mcm5p1f_ca_w_1_200_s_0_840=1.64e-04 mcm5p1f_cc_w_1_200_s_0_840=2.51e-11 mcm5p1f_cf_w_1_200_s_0_840=4.00e-11
+  mcm5p1f_ca_w_1_200_s_1_260=1.64e-04 mcm5p1f_cc_w_1_200_s_1_260=1.48e-11 mcm5p1f_cf_w_1_200_s_1_260=4.78e-11
+  mcm5p1f_ca_w_1_200_s_2_310=1.64e-04 mcm5p1f_cc_w_1_200_s_2_310=5.24e-12 mcm5p1f_cf_w_1_200_s_2_310=5.64e-11
+  mcm5p1f_ca_w_1_200_s_5_250=1.64e-04 mcm5p1f_cc_w_1_200_s_5_250=5.65e-13 mcm5p1f_cf_w_1_200_s_5_250=6.09e-11
+  mcrdlp1f_ca_w_0_150_s_0_210=1.58e-04 mcrdlp1f_cc_w_0_150_s_0_210=8.86e-11 mcrdlp1f_cf_w_0_150_s_0_210=1.37e-11
+  mcrdlp1f_ca_w_0_150_s_0_263=1.58e-04 mcrdlp1f_cc_w_0_150_s_0_263=6.90e-11 mcrdlp1f_cf_w_0_150_s_0_263=1.67e-11
+  mcrdlp1f_ca_w_0_150_s_0_315=1.58e-04 mcrdlp1f_cc_w_0_150_s_0_315=5.72e-11 mcrdlp1f_cf_w_0_150_s_0_315=1.96e-11
+  mcrdlp1f_ca_w_0_150_s_0_420=1.58e-04 mcrdlp1f_cc_w_0_150_s_0_420=4.22e-11 mcrdlp1f_cf_w_0_150_s_0_420=2.48e-11
+  mcrdlp1f_ca_w_0_150_s_0_525=1.58e-04 mcrdlp1f_cc_w_0_150_s_0_525=3.34e-11 mcrdlp1f_cf_w_0_150_s_0_525=2.90e-11
+  mcrdlp1f_ca_w_0_150_s_0_630=1.58e-04 mcrdlp1f_cc_w_0_150_s_0_630=2.73e-11 mcrdlp1f_cf_w_0_150_s_0_630=3.25e-11
+  mcrdlp1f_ca_w_0_150_s_0_840=1.58e-04 mcrdlp1f_cc_w_0_150_s_0_840=1.93e-11 mcrdlp1f_cf_w_0_150_s_0_840=3.81e-11
+  mcrdlp1f_ca_w_0_150_s_1_260=1.58e-04 mcrdlp1f_cc_w_0_150_s_1_260=1.06e-11 mcrdlp1f_cf_w_0_150_s_1_260=4.53e-11
+  mcrdlp1f_ca_w_0_150_s_2_310=1.58e-04 mcrdlp1f_cc_w_0_150_s_2_310=3.93e-12 mcrdlp1f_cf_w_0_150_s_2_310=5.13e-11
+  mcrdlp1f_ca_w_0_150_s_5_250=1.58e-04 mcrdlp1f_cc_w_0_150_s_5_250=7.38e-13 mcrdlp1f_cf_w_0_150_s_5_250=5.45e-11
+  mcrdlp1f_ca_w_1_200_s_0_210=1.58e-04 mcrdlp1f_cc_w_1_200_s_0_210=1.06e-10 mcrdlp1f_cf_w_1_200_s_0_210=1.36e-11
+  mcrdlp1f_ca_w_1_200_s_0_263=1.58e-04 mcrdlp1f_cc_w_1_200_s_0_263=8.49e-11 mcrdlp1f_cf_w_1_200_s_0_263=1.67e-11
+  mcrdlp1f_ca_w_1_200_s_0_315=1.58e-04 mcrdlp1f_cc_w_1_200_s_0_315=7.18e-11 mcrdlp1f_cf_w_1_200_s_0_315=1.96e-11
+  mcrdlp1f_ca_w_1_200_s_0_420=1.58e-04 mcrdlp1f_cc_w_1_200_s_0_420=5.53e-11 mcrdlp1f_cf_w_1_200_s_0_420=2.47e-11
+  mcrdlp1f_ca_w_1_200_s_0_525=1.58e-04 mcrdlp1f_cc_w_1_200_s_0_525=4.51e-11 mcrdlp1f_cf_w_1_200_s_0_525=2.91e-11
+  mcrdlp1f_ca_w_1_200_s_0_630=1.58e-04 mcrdlp1f_cc_w_1_200_s_0_630=3.80e-11 mcrdlp1f_cf_w_1_200_s_0_630=3.27e-11
+  mcrdlp1f_ca_w_1_200_s_0_840=1.58e-04 mcrdlp1f_cc_w_1_200_s_0_840=2.87e-11 mcrdlp1f_cf_w_1_200_s_0_840=3.86e-11
+  mcrdlp1f_ca_w_1_200_s_1_260=1.58e-04 mcrdlp1f_cc_w_1_200_s_1_260=1.84e-11 mcrdlp1f_cf_w_1_200_s_1_260=4.65e-11
+  mcrdlp1f_ca_w_1_200_s_2_310=1.58e-04 mcrdlp1f_cc_w_1_200_s_2_310=7.89e-12 mcrdlp1f_cf_w_1_200_s_2_310=5.57e-11
+  mcrdlp1f_ca_w_1_200_s_5_250=1.58e-04 mcrdlp1f_cc_w_1_200_s_5_250=1.72e-12 mcrdlp1f_cf_w_1_200_s_5_250=6.16e-11
+  mcm1l1f_ca_w_0_170_s_0_180=2.66e-04 mcm1l1f_cc_w_0_170_s_0_180=7.99e-11 mcm1l1f_cf_w_0_170_s_0_180=1.76e-11
+  mcm1l1f_ca_w_0_170_s_0_225=2.66e-04 mcm1l1f_cc_w_0_170_s_0_225=6.04e-11 mcm1l1f_cf_w_0_170_s_0_225=2.19e-11
+  mcm1l1f_ca_w_0_170_s_0_270=2.66e-04 mcm1l1f_cc_w_0_170_s_0_270=4.79e-11 mcm1l1f_cf_w_0_170_s_0_270=2.58e-11
+  mcm1l1f_ca_w_0_170_s_0_360=2.66e-04 mcm1l1f_cc_w_0_170_s_0_360=3.23e-11 mcm1l1f_cf_w_0_170_s_0_360=3.27e-11
+  mcm1l1f_ca_w_0_170_s_0_450=2.66e-04 mcm1l1f_cc_w_0_170_s_0_450=2.29e-11 mcm1l1f_cf_w_0_170_s_0_450=3.82e-11
+  mcm1l1f_ca_w_0_170_s_0_540=2.66e-04 mcm1l1f_cc_w_0_170_s_0_540=1.66e-11 mcm1l1f_cf_w_0_170_s_0_540=4.25e-11
+  mcm1l1f_ca_w_0_170_s_0_720=2.66e-04 mcm1l1f_cc_w_0_170_s_0_720=9.06e-12 mcm1l1f_cf_w_0_170_s_0_720=4.85e-11
+  mcm1l1f_ca_w_0_170_s_1_080=2.66e-04 mcm1l1f_cc_w_0_170_s_1_080=2.90e-12 mcm1l1f_cf_w_0_170_s_1_080=5.41e-11
+  mcm1l1f_ca_w_0_170_s_1_980=2.66e-04 mcm1l1f_cc_w_0_170_s_1_980=2.40e-13 mcm1l1f_cf_w_0_170_s_1_980=5.67e-11
+  mcm1l1f_ca_w_0_170_s_4_500=2.66e-04 mcm1l1f_cc_w_0_170_s_4_500=0.00e+00 mcm1l1f_cf_w_0_170_s_4_500=5.69e-11
+  mcm1l1f_ca_w_1_360_s_0_180=2.66e-04 mcm1l1f_cc_w_1_360_s_0_180=8.29e-11 mcm1l1f_cf_w_1_360_s_0_180=1.74e-11
+  mcm1l1f_ca_w_1_360_s_0_225=2.66e-04 mcm1l1f_cc_w_1_360_s_0_225=6.30e-11 mcm1l1f_cf_w_1_360_s_0_225=2.17e-11
+  mcm1l1f_ca_w_1_360_s_0_270=2.66e-04 mcm1l1f_cc_w_1_360_s_0_270=5.01e-11 mcm1l1f_cf_w_1_360_s_0_270=2.57e-11
+  mcm1l1f_ca_w_1_360_s_0_360=2.66e-04 mcm1l1f_cc_w_1_360_s_0_360=3.40e-11 mcm1l1f_cf_w_1_360_s_0_360=3.26e-11
+  mcm1l1f_ca_w_1_360_s_0_450=2.66e-04 mcm1l1f_cc_w_1_360_s_0_450=2.43e-11 mcm1l1f_cf_w_1_360_s_0_450=3.82e-11
+  mcm1l1f_ca_w_1_360_s_0_540=2.66e-04 mcm1l1f_cc_w_1_360_s_0_540=1.78e-11 mcm1l1f_cf_w_1_360_s_0_540=4.26e-11
+  mcm1l1f_ca_w_1_360_s_0_720=2.66e-04 mcm1l1f_cc_w_1_360_s_0_720=9.85e-12 mcm1l1f_cf_w_1_360_s_0_720=4.88e-11
+  mcm1l1f_ca_w_1_360_s_1_080=2.66e-04 mcm1l1f_cc_w_1_360_s_1_080=3.24e-12 mcm1l1f_cf_w_1_360_s_1_080=5.47e-11
+  mcm1l1f_ca_w_1_360_s_1_980=2.66e-04 mcm1l1f_cc_w_1_360_s_1_980=2.35e-13 mcm1l1f_cf_w_1_360_s_1_980=5.76e-11
+  mcm1l1f_ca_w_1_360_s_4_500=2.66e-04 mcm1l1f_cc_w_1_360_s_4_500=0.00e+00 mcm1l1f_cf_w_1_360_s_4_500=5.78e-11
+  mcm1l1d_ca_w_0_170_s_0_180=2.87e-04 mcm1l1d_cc_w_0_170_s_0_180=7.74e-11 mcm1l1d_cf_w_0_170_s_0_180=1.90e-11
+  mcm1l1d_ca_w_0_170_s_0_225=2.87e-04 mcm1l1d_cc_w_0_170_s_0_225=5.78e-11 mcm1l1d_cf_w_0_170_s_0_225=2.37e-11
+  mcm1l1d_ca_w_0_170_s_0_270=2.87e-04 mcm1l1d_cc_w_0_170_s_0_270=4.51e-11 mcm1l1d_cf_w_0_170_s_0_270=2.79e-11
+  mcm1l1d_ca_w_0_170_s_0_360=2.87e-04 mcm1l1d_cc_w_0_170_s_0_360=2.95e-11 mcm1l1d_cf_w_0_170_s_0_360=3.53e-11
+  mcm1l1d_ca_w_0_170_s_0_450=2.87e-04 mcm1l1d_cc_w_0_170_s_0_450=2.02e-11 mcm1l1d_cf_w_0_170_s_0_450=4.10e-11
+  mcm1l1d_ca_w_0_170_s_0_540=2.87e-04 mcm1l1d_cc_w_0_170_s_0_540=1.40e-11 mcm1l1d_cf_w_0_170_s_0_540=4.55e-11
+  mcm1l1d_ca_w_0_170_s_0_720=2.87e-04 mcm1l1d_cc_w_0_170_s_0_720=7.08e-12 mcm1l1d_cf_w_0_170_s_0_720=5.13e-11
+  mcm1l1d_ca_w_0_170_s_1_080=2.87e-04 mcm1l1d_cc_w_0_170_s_1_080=1.86e-12 mcm1l1d_cf_w_0_170_s_1_080=5.62e-11
+  mcm1l1d_ca_w_0_170_s_1_980=2.87e-04 mcm1l1d_cc_w_0_170_s_1_980=1.15e-13 mcm1l1d_cf_w_0_170_s_1_980=5.79e-11
+  mcm1l1d_ca_w_0_170_s_4_500=2.87e-04 mcm1l1d_cc_w_0_170_s_4_500=4.00e-14 mcm1l1d_cf_w_0_170_s_4_500=5.79e-11
+  mcm1l1d_ca_w_1_360_s_0_180=2.87e-04 mcm1l1d_cc_w_1_360_s_0_180=7.92e-11 mcm1l1d_cf_w_1_360_s_0_180=1.88e-11
+  mcm1l1d_ca_w_1_360_s_0_225=2.87e-04 mcm1l1d_cc_w_1_360_s_0_225=5.94e-11 mcm1l1d_cf_w_1_360_s_0_225=2.35e-11
+  mcm1l1d_ca_w_1_360_s_0_270=2.87e-04 mcm1l1d_cc_w_1_360_s_0_270=4.65e-11 mcm1l1d_cf_w_1_360_s_0_270=2.77e-11
+  mcm1l1d_ca_w_1_360_s_0_360=2.87e-04 mcm1l1d_cc_w_1_360_s_0_360=3.05e-11 mcm1l1d_cf_w_1_360_s_0_360=3.51e-11
+  mcm1l1d_ca_w_1_360_s_0_450=2.87e-04 mcm1l1d_cc_w_1_360_s_0_450=2.11e-11 mcm1l1d_cf_w_1_360_s_0_450=4.09e-11
+  mcm1l1d_ca_w_1_360_s_0_540=2.87e-04 mcm1l1d_cc_w_1_360_s_0_540=1.47e-11 mcm1l1d_cf_w_1_360_s_0_540=4.54e-11
+  mcm1l1d_ca_w_1_360_s_0_720=2.87e-04 mcm1l1d_cc_w_1_360_s_0_720=7.40e-12 mcm1l1d_cf_w_1_360_s_0_720=5.13e-11
+  mcm1l1d_ca_w_1_360_s_1_080=2.87e-04 mcm1l1d_cc_w_1_360_s_1_080=1.95e-12 mcm1l1d_cf_w_1_360_s_1_080=5.63e-11
+  mcm1l1d_ca_w_1_360_s_1_980=2.87e-04 mcm1l1d_cc_w_1_360_s_1_980=1.50e-13 mcm1l1d_cf_w_1_360_s_1_980=5.81e-11
+  mcm1l1d_ca_w_1_360_s_4_500=2.87e-04 mcm1l1d_cc_w_1_360_s_4_500=2.58e-26 mcm1l1d_cf_w_1_360_s_4_500=5.82e-11
+  mcm1l1p1_ca_w_0_170_s_0_180=3.91e-04 mcm1l1p1_cc_w_0_170_s_0_180=6.95e-11 mcm1l1p1_cf_w_0_170_s_0_180=2.56e-11
+  mcm1l1p1_ca_w_0_170_s_0_225=3.91e-04 mcm1l1p1_cc_w_0_170_s_0_225=4.98e-11 mcm1l1p1_cf_w_0_170_s_0_225=3.19e-11
+  mcm1l1p1_ca_w_0_170_s_0_270=3.91e-04 mcm1l1p1_cc_w_0_170_s_0_270=3.72e-11 mcm1l1p1_cf_w_0_170_s_0_270=3.73e-11
+  mcm1l1p1_ca_w_0_170_s_0_360=3.91e-04 mcm1l1p1_cc_w_0_170_s_0_360=2.20e-11 mcm1l1p1_cf_w_0_170_s_0_360=4.62e-11
+  mcm1l1p1_ca_w_0_170_s_0_450=3.91e-04 mcm1l1p1_cc_w_0_170_s_0_450=1.34e-11 mcm1l1p1_cf_w_0_170_s_0_450=5.25e-11
+  mcm1l1p1_ca_w_0_170_s_0_540=3.91e-04 mcm1l1p1_cc_w_0_170_s_0_540=8.33e-12 mcm1l1p1_cf_w_0_170_s_0_540=5.68e-11
+  mcm1l1p1_ca_w_0_170_s_0_720=3.91e-04 mcm1l1p1_cc_w_0_170_s_0_720=3.23e-12 mcm1l1p1_cf_w_0_170_s_0_720=6.14e-11
+  mcm1l1p1_ca_w_0_170_s_1_080=3.91e-04 mcm1l1p1_cc_w_0_170_s_1_080=5.70e-13 mcm1l1p1_cf_w_0_170_s_1_080=6.40e-11
+  mcm1l1p1_ca_w_0_170_s_1_980=3.91e-04 mcm1l1p1_cc_w_0_170_s_1_980=1.00e-14 mcm1l1p1_cf_w_0_170_s_1_980=6.45e-11
+  mcm1l1p1_ca_w_0_170_s_4_500=3.91e-04 mcm1l1p1_cc_w_0_170_s_4_500=5.00e-15 mcm1l1p1_cf_w_0_170_s_4_500=6.44e-11
+  mcm1l1p1_ca_w_1_360_s_0_180=3.91e-04 mcm1l1p1_cc_w_1_360_s_0_180=6.99e-11 mcm1l1p1_cf_w_1_360_s_0_180=2.53e-11
+  mcm1l1p1_ca_w_1_360_s_0_225=3.91e-04 mcm1l1p1_cc_w_1_360_s_0_225=5.01e-11 mcm1l1p1_cf_w_1_360_s_0_225=3.14e-11
+  mcm1l1p1_ca_w_1_360_s_0_270=3.91e-04 mcm1l1p1_cc_w_1_360_s_0_270=3.75e-11 mcm1l1p1_cf_w_1_360_s_0_270=3.69e-11
+  mcm1l1p1_ca_w_1_360_s_0_360=3.91e-04 mcm1l1p1_cc_w_1_360_s_0_360=2.23e-11 mcm1l1p1_cf_w_1_360_s_0_360=4.58e-11
+  mcm1l1p1_ca_w_1_360_s_0_450=3.91e-04 mcm1l1p1_cc_w_1_360_s_0_450=1.36e-11 mcm1l1p1_cf_w_1_360_s_0_450=5.20e-11
+  mcm1l1p1_ca_w_1_360_s_0_540=3.91e-04 mcm1l1p1_cc_w_1_360_s_0_540=8.40e-12 mcm1l1p1_cf_w_1_360_s_0_540=5.64e-11
+  mcm1l1p1_ca_w_1_360_s_0_720=3.91e-04 mcm1l1p1_cc_w_1_360_s_0_720=3.30e-12 mcm1l1p1_cf_w_1_360_s_0_720=6.10e-11
+  mcm1l1p1_ca_w_1_360_s_1_080=3.91e-04 mcm1l1p1_cc_w_1_360_s_1_080=5.50e-13 mcm1l1p1_cf_w_1_360_s_1_080=6.37e-11
+  mcm1l1p1_ca_w_1_360_s_1_980=3.91e-04 mcm1l1p1_cc_w_1_360_s_1_980=5.00e-14 mcm1l1p1_cf_w_1_360_s_1_980=6.42e-11
+  mcm1l1p1_ca_w_1_360_s_4_500=3.91e-04 mcm1l1p1_cc_w_1_360_s_4_500=2.58e-26 mcm1l1p1_cf_w_1_360_s_4_500=6.41e-11
+  mcm2l1f_ca_w_0_170_s_0_180=1.02e-04 mcm2l1f_cc_w_0_170_s_0_180=9.39e-11 mcm2l1f_cf_w_0_170_s_0_180=7.27e-12
+  mcm2l1f_ca_w_0_170_s_0_225=1.02e-04 mcm2l1f_cc_w_0_170_s_0_225=7.42e-11 mcm2l1f_cf_w_0_170_s_0_225=9.38e-12
+  mcm2l1f_ca_w_0_170_s_0_270=1.02e-04 mcm2l1f_cc_w_0_170_s_0_270=6.17e-11 mcm2l1f_cf_w_0_170_s_0_270=1.14e-11
+  mcm2l1f_ca_w_0_170_s_0_360=1.02e-04 mcm2l1f_cc_w_0_170_s_0_360=4.56e-11 mcm2l1f_cf_w_0_170_s_0_360=1.53e-11
+  mcm2l1f_ca_w_0_170_s_0_450=1.02e-04 mcm2l1f_cc_w_0_170_s_0_450=3.55e-11 mcm2l1f_cf_w_0_170_s_0_450=1.89e-11
+  mcm2l1f_ca_w_0_170_s_0_540=1.02e-04 mcm2l1f_cc_w_0_170_s_0_540=2.84e-11 mcm2l1f_cf_w_0_170_s_0_540=2.21e-11
+  mcm2l1f_ca_w_0_170_s_0_720=1.02e-04 mcm2l1f_cc_w_0_170_s_0_720=1.89e-11 mcm2l1f_cf_w_0_170_s_0_720=2.74e-11
+  mcm2l1f_ca_w_0_170_s_1_080=1.02e-04 mcm2l1f_cc_w_0_170_s_1_080=8.93e-12 mcm2l1f_cf_w_0_170_s_1_080=3.46e-11
+  mcm2l1f_ca_w_0_170_s_1_980=1.02e-04 mcm2l1f_cc_w_0_170_s_1_980=1.50e-12 mcm2l1f_cf_w_0_170_s_1_980=4.13e-11
+  mcm2l1f_ca_w_0_170_s_4_500=1.02e-04 mcm2l1f_cc_w_0_170_s_4_500=1.00e-14 mcm2l1f_cf_w_0_170_s_4_500=4.27e-11
+  mcm2l1f_ca_w_1_360_s_0_180=1.02e-04 mcm2l1f_cc_w_1_360_s_0_180=9.95e-11 mcm2l1f_cf_w_1_360_s_0_180=7.24e-12
+  mcm2l1f_ca_w_1_360_s_0_225=1.02e-04 mcm2l1f_cc_w_1_360_s_0_225=7.90e-11 mcm2l1f_cf_w_1_360_s_0_225=9.34e-12
+  mcm2l1f_ca_w_1_360_s_0_270=1.02e-04 mcm2l1f_cc_w_1_360_s_0_270=6.58e-11 mcm2l1f_cf_w_1_360_s_0_270=1.14e-11
+  mcm2l1f_ca_w_1_360_s_0_360=1.02e-04 mcm2l1f_cc_w_1_360_s_0_360=4.88e-11 mcm2l1f_cf_w_1_360_s_0_360=1.53e-11
+  mcm2l1f_ca_w_1_360_s_0_450=1.02e-04 mcm2l1f_cc_w_1_360_s_0_450=3.81e-11 mcm2l1f_cf_w_1_360_s_0_450=1.89e-11
+  mcm2l1f_ca_w_1_360_s_0_540=1.02e-04 mcm2l1f_cc_w_1_360_s_0_540=3.04e-11 mcm2l1f_cf_w_1_360_s_0_540=2.22e-11
+  mcm2l1f_ca_w_1_360_s_0_720=1.02e-04 mcm2l1f_cc_w_1_360_s_0_720=2.03e-11 mcm2l1f_cf_w_1_360_s_0_720=2.77e-11
+  mcm2l1f_ca_w_1_360_s_1_080=1.02e-04 mcm2l1f_cc_w_1_360_s_1_080=9.70e-12 mcm2l1f_cf_w_1_360_s_1_080=3.54e-11
+  mcm2l1f_ca_w_1_360_s_1_980=1.02e-04 mcm2l1f_cc_w_1_360_s_1_980=1.65e-12 mcm2l1f_cf_w_1_360_s_1_980=4.25e-11
+  mcm2l1f_ca_w_1_360_s_4_500=1.02e-04 mcm2l1f_cc_w_1_360_s_4_500=1.00e-13 mcm2l1f_cf_w_1_360_s_4_500=4.41e-11
+  mcm2l1d_ca_w_0_170_s_0_180=1.23e-04 mcm2l1d_cc_w_0_170_s_0_180=9.12e-11 mcm2l1d_cf_w_0_170_s_0_180=8.72e-12
+  mcm2l1d_ca_w_0_170_s_0_225=1.23e-04 mcm2l1d_cc_w_0_170_s_0_225=7.15e-11 mcm2l1d_cf_w_0_170_s_0_225=1.12e-11
+  mcm2l1d_ca_w_0_170_s_0_270=1.23e-04 mcm2l1d_cc_w_0_170_s_0_270=5.88e-11 mcm2l1d_cf_w_0_170_s_0_270=1.37e-11
+  mcm2l1d_ca_w_0_170_s_0_360=1.23e-04 mcm2l1d_cc_w_0_170_s_0_360=4.26e-11 mcm2l1d_cf_w_0_170_s_0_360=1.82e-11
+  mcm2l1d_ca_w_0_170_s_0_450=1.23e-04 mcm2l1d_cc_w_0_170_s_0_450=3.24e-11 mcm2l1d_cf_w_0_170_s_0_450=2.23e-11
+  mcm2l1d_ca_w_0_170_s_0_540=1.23e-04 mcm2l1d_cc_w_0_170_s_0_540=2.53e-11 mcm2l1d_cf_w_0_170_s_0_540=2.59e-11
+  mcm2l1d_ca_w_0_170_s_0_720=1.23e-04 mcm2l1d_cc_w_0_170_s_0_720=1.61e-11 mcm2l1d_cf_w_0_170_s_0_720=3.17e-11
+  mcm2l1d_ca_w_0_170_s_1_080=1.23e-04 mcm2l1d_cc_w_0_170_s_1_080=6.80e-12 mcm2l1d_cf_w_0_170_s_1_080=3.89e-11
+  mcm2l1d_ca_w_0_170_s_1_980=1.23e-04 mcm2l1d_cc_w_0_170_s_1_980=9.10e-13 mcm2l1d_cf_w_0_170_s_1_980=4.44e-11
+  mcm2l1d_ca_w_0_170_s_4_500=1.23e-04 mcm2l1d_cc_w_0_170_s_4_500=0.00e+00 mcm2l1d_cf_w_0_170_s_4_500=4.52e-11
+  mcm2l1d_ca_w_1_360_s_0_180=1.23e-04 mcm2l1d_cc_w_1_360_s_0_180=9.56e-11 mcm2l1d_cf_w_1_360_s_0_180=8.70e-12
+  mcm2l1d_ca_w_1_360_s_0_225=1.23e-04 mcm2l1d_cc_w_1_360_s_0_225=7.52e-11 mcm2l1d_cf_w_1_360_s_0_225=1.12e-11
+  mcm2l1d_ca_w_1_360_s_0_270=1.23e-04 mcm2l1d_cc_w_1_360_s_0_270=6.20e-11 mcm2l1d_cf_w_1_360_s_0_270=1.36e-11
+  mcm2l1d_ca_w_1_360_s_0_360=1.23e-04 mcm2l1d_cc_w_1_360_s_0_360=4.50e-11 mcm2l1d_cf_w_1_360_s_0_360=1.82e-11
+  mcm2l1d_ca_w_1_360_s_0_450=1.23e-04 mcm2l1d_cc_w_1_360_s_0_450=3.43e-11 mcm2l1d_cf_w_1_360_s_0_450=2.23e-11
+  mcm2l1d_ca_w_1_360_s_0_540=1.23e-04 mcm2l1d_cc_w_1_360_s_0_540=2.68e-11 mcm2l1d_cf_w_1_360_s_0_540=2.60e-11
+  mcm2l1d_ca_w_1_360_s_0_720=1.23e-04 mcm2l1d_cc_w_1_360_s_0_720=1.71e-11 mcm2l1d_cf_w_1_360_s_0_720=3.20e-11
+  mcm2l1d_ca_w_1_360_s_1_080=1.23e-04 mcm2l1d_cc_w_1_360_s_1_080=7.35e-12 mcm2l1d_cf_w_1_360_s_1_080=3.95e-11
+  mcm2l1d_ca_w_1_360_s_1_980=1.23e-04 mcm2l1d_cc_w_1_360_s_1_980=1.00e-12 mcm2l1d_cf_w_1_360_s_1_980=4.54e-11
+  mcm2l1d_ca_w_1_360_s_4_500=1.23e-04 mcm2l1d_cc_w_1_360_s_4_500=5.00e-14 mcm2l1d_cf_w_1_360_s_4_500=4.63e-11
+  mcm2l1p1_ca_w_0_170_s_0_180=2.27e-04 mcm2l1p1_cc_w_0_170_s_0_180=8.33e-11 mcm2l1p1_cf_w_0_170_s_0_180=1.55e-11
+  mcm2l1p1_ca_w_0_170_s_0_225=2.27e-04 mcm2l1p1_cc_w_0_170_s_0_225=6.34e-11 mcm2l1p1_cf_w_0_170_s_0_225=1.97e-11
+  mcm2l1p1_ca_w_0_170_s_0_270=2.27e-04 mcm2l1p1_cc_w_0_170_s_0_270=5.05e-11 mcm2l1p1_cf_w_0_170_s_0_270=2.36e-11
+  mcm2l1p1_ca_w_0_170_s_0_360=2.27e-04 mcm2l1p1_cc_w_0_170_s_0_360=3.43e-11 mcm2l1p1_cf_w_0_170_s_0_360=3.06e-11
+  mcm2l1p1_ca_w_0_170_s_0_450=2.27e-04 mcm2l1p1_cc_w_0_170_s_0_450=2.44e-11 mcm2l1p1_cf_w_0_170_s_0_450=3.62e-11
+  mcm2l1p1_ca_w_0_170_s_0_540=2.27e-04 mcm2l1p1_cc_w_0_170_s_0_540=1.78e-11 mcm2l1p1_cf_w_0_170_s_0_540=4.07e-11
+  mcm2l1p1_ca_w_0_170_s_0_720=2.27e-04 mcm2l1p1_cc_w_0_170_s_0_720=9.74e-12 mcm2l1p1_cf_w_0_170_s_0_720=4.70e-11
+  mcm2l1p1_ca_w_0_170_s_1_080=2.27e-04 mcm2l1p1_cc_w_0_170_s_1_080=3.12e-12 mcm2l1p1_cf_w_0_170_s_1_080=5.30e-11
+  mcm2l1p1_ca_w_0_170_s_1_980=2.27e-04 mcm2l1p1_cc_w_0_170_s_1_980=2.65e-13 mcm2l1p1_cf_w_0_170_s_1_980=5.58e-11
+  mcm2l1p1_ca_w_0_170_s_4_500=2.27e-04 mcm2l1p1_cc_w_0_170_s_4_500=5.00e-15 mcm2l1p1_cf_w_0_170_s_4_500=5.60e-11
+  mcm2l1p1_ca_w_1_360_s_0_180=2.27e-04 mcm2l1p1_cc_w_1_360_s_0_180=8.66e-11 mcm2l1p1_cf_w_1_360_s_0_180=1.55e-11
+  mcm2l1p1_ca_w_1_360_s_0_225=2.27e-04 mcm2l1p1_cc_w_1_360_s_0_225=6.63e-11 mcm2l1p1_cf_w_1_360_s_0_225=1.96e-11
+  mcm2l1p1_ca_w_1_360_s_0_270=2.27e-04 mcm2l1p1_cc_w_1_360_s_0_270=5.29e-11 mcm2l1p1_cf_w_1_360_s_0_270=2.35e-11
+  mcm2l1p1_ca_w_1_360_s_0_360=2.27e-04 mcm2l1p1_cc_w_1_360_s_0_360=3.62e-11 mcm2l1p1_cf_w_1_360_s_0_360=3.05e-11
+  mcm2l1p1_ca_w_1_360_s_0_450=2.27e-04 mcm2l1p1_cc_w_1_360_s_0_450=2.59e-11 mcm2l1p1_cf_w_1_360_s_0_450=3.62e-11
+  mcm2l1p1_ca_w_1_360_s_0_540=2.27e-04 mcm2l1p1_cc_w_1_360_s_0_540=1.90e-11 mcm2l1p1_cf_w_1_360_s_0_540=4.08e-11
+  mcm2l1p1_ca_w_1_360_s_0_720=2.27e-04 mcm2l1p1_cc_w_1_360_s_0_720=1.05e-11 mcm2l1p1_cf_w_1_360_s_0_720=4.74e-11
+  mcm2l1p1_ca_w_1_360_s_1_080=2.27e-04 mcm2l1p1_cc_w_1_360_s_1_080=3.40e-12 mcm2l1p1_cf_w_1_360_s_1_080=5.37e-11
+  mcm2l1p1_ca_w_1_360_s_1_980=2.27e-04 mcm2l1p1_cc_w_1_360_s_1_980=3.00e-13 mcm2l1p1_cf_w_1_360_s_1_980=5.67e-11
+  mcm2l1p1_ca_w_1_360_s_4_500=2.27e-04 mcm2l1p1_cc_w_1_360_s_4_500=0.00e+00 mcm2l1p1_cf_w_1_360_s_4_500=5.70e-11
+  mcm3l1f_ca_w_0_170_s_0_180=7.60e-05 mcm3l1f_cc_w_0_170_s_0_180=9.72e-11 mcm3l1f_cf_w_0_170_s_0_180=5.46e-12
+  mcm3l1f_ca_w_0_170_s_0_225=7.60e-05 mcm3l1f_cc_w_0_170_s_0_225=7.80e-11 mcm3l1f_cf_w_0_170_s_0_225=7.06e-12
+  mcm3l1f_ca_w_0_170_s_0_270=7.60e-05 mcm3l1f_cc_w_0_170_s_0_270=6.57e-11 mcm3l1f_cf_w_0_170_s_0_270=8.62e-12
+  mcm3l1f_ca_w_0_170_s_0_360=7.60e-05 mcm3l1f_cc_w_0_170_s_0_360=5.01e-11 mcm3l1f_cf_w_0_170_s_0_360=1.17e-11
+  mcm3l1f_ca_w_0_170_s_0_450=7.60e-05 mcm3l1f_cc_w_0_170_s_0_450=4.03e-11 mcm3l1f_cf_w_0_170_s_0_450=1.45e-11
+  mcm3l1f_ca_w_0_170_s_0_540=7.60e-05 mcm3l1f_cc_w_0_170_s_0_540=3.32e-11 mcm3l1f_cf_w_0_170_s_0_540=1.72e-11
+  mcm3l1f_ca_w_0_170_s_0_720=7.60e-05 mcm3l1f_cc_w_0_170_s_0_720=2.37e-11 mcm3l1f_cf_w_0_170_s_0_720=2.17e-11
+  mcm3l1f_ca_w_0_170_s_1_080=7.60e-05 mcm3l1f_cc_w_0_170_s_1_080=1.31e-11 mcm3l1f_cf_w_0_170_s_1_080=2.85e-11
+  mcm3l1f_ca_w_0_170_s_1_980=7.60e-05 mcm3l1f_cc_w_0_170_s_1_980=3.39e-12 mcm3l1f_cf_w_0_170_s_1_980=3.66e-11
+  mcm3l1f_ca_w_0_170_s_4_500=7.60e-05 mcm3l1f_cc_w_0_170_s_4_500=1.25e-13 mcm3l1f_cf_w_0_170_s_4_500=3.97e-11
+  mcm3l1f_ca_w_1_360_s_0_180=7.60e-05 mcm3l1f_cc_w_1_360_s_0_180=1.07e-10 mcm3l1f_cf_w_1_360_s_0_180=5.44e-12
+  mcm3l1f_ca_w_1_360_s_0_225=7.60e-05 mcm3l1f_cc_w_1_360_s_0_225=8.64e-11 mcm3l1f_cf_w_1_360_s_0_225=7.05e-12
+  mcm3l1f_ca_w_1_360_s_0_270=7.60e-05 mcm3l1f_cc_w_1_360_s_0_270=7.30e-11 mcm3l1f_cf_w_1_360_s_0_270=8.63e-12
+  mcm3l1f_ca_w_1_360_s_0_360=7.60e-05 mcm3l1f_cc_w_1_360_s_0_360=5.60e-11 mcm3l1f_cf_w_1_360_s_0_360=1.17e-11
+  mcm3l1f_ca_w_1_360_s_0_450=7.60e-05 mcm3l1f_cc_w_1_360_s_0_450=4.52e-11 mcm3l1f_cf_w_1_360_s_0_450=1.45e-11
+  mcm3l1f_ca_w_1_360_s_0_540=7.60e-05 mcm3l1f_cc_w_1_360_s_0_540=3.74e-11 mcm3l1f_cf_w_1_360_s_0_540=1.72e-11
+  mcm3l1f_ca_w_1_360_s_0_720=7.60e-05 mcm3l1f_cc_w_1_360_s_0_720=2.69e-11 mcm3l1f_cf_w_1_360_s_0_720=2.20e-11
+  mcm3l1f_ca_w_1_360_s_1_080=7.60e-05 mcm3l1f_cc_w_1_360_s_1_080=1.51e-11 mcm3l1f_cf_w_1_360_s_1_080=2.93e-11
+  mcm3l1f_ca_w_1_360_s_1_980=7.60e-05 mcm3l1f_cc_w_1_360_s_1_980=4.05e-12 mcm3l1f_cf_w_1_360_s_1_980=3.83e-11
+  mcm3l1f_ca_w_1_360_s_4_500=7.60e-05 mcm3l1f_cc_w_1_360_s_4_500=1.65e-13 mcm3l1f_cf_w_1_360_s_4_500=4.21e-11
+  mcm3l1d_ca_w_0_170_s_0_180=9.72e-05 mcm3l1d_cc_w_0_170_s_0_180=9.46e-11 mcm3l1d_cf_w_0_170_s_0_180=6.93e-12
+  mcm3l1d_ca_w_0_170_s_0_225=9.72e-05 mcm3l1d_cc_w_0_170_s_0_225=7.53e-11 mcm3l1d_cf_w_0_170_s_0_225=8.95e-12
+  mcm3l1d_ca_w_0_170_s_0_270=9.72e-05 mcm3l1d_cc_w_0_170_s_0_270=6.28e-11 mcm3l1d_cf_w_0_170_s_0_270=1.09e-11
+  mcm3l1d_ca_w_0_170_s_0_360=9.72e-05 mcm3l1d_cc_w_0_170_s_0_360=4.70e-11 mcm3l1d_cf_w_0_170_s_0_360=1.47e-11
+  mcm3l1d_ca_w_0_170_s_0_450=9.72e-05 mcm3l1d_cc_w_0_170_s_0_450=3.71e-11 mcm3l1d_cf_w_0_170_s_0_450=1.80e-11
+  mcm3l1d_ca_w_0_170_s_0_540=9.72e-05 mcm3l1d_cc_w_0_170_s_0_540=3.00e-11 mcm3l1d_cf_w_0_170_s_0_540=2.12e-11
+  mcm3l1d_ca_w_0_170_s_0_720=9.72e-05 mcm3l1d_cc_w_0_170_s_0_720=2.06e-11 mcm3l1d_cf_w_0_170_s_0_720=2.64e-11
+  mcm3l1d_ca_w_0_170_s_1_080=9.72e-05 mcm3l1d_cc_w_0_170_s_1_080=1.05e-11 mcm3l1d_cf_w_0_170_s_1_080=3.36e-11
+  mcm3l1d_ca_w_0_170_s_1_980=9.72e-05 mcm3l1d_cc_w_0_170_s_1_980=2.28e-12 mcm3l1d_cf_w_0_170_s_1_980=4.08e-11
+  mcm3l1d_ca_w_0_170_s_4_500=9.72e-05 mcm3l1d_cc_w_0_170_s_4_500=6.00e-14 mcm3l1d_cf_w_0_170_s_4_500=4.29e-11
+  mcm3l1d_ca_w_1_360_s_0_180=9.72e-05 mcm3l1d_cc_w_1_360_s_0_180=1.03e-10 mcm3l1d_cf_w_1_360_s_0_180=6.91e-12
+  mcm3l1d_ca_w_1_360_s_0_225=9.72e-05 mcm3l1d_cc_w_1_360_s_0_225=8.24e-11 mcm3l1d_cf_w_1_360_s_0_225=8.93e-12
+  mcm3l1d_ca_w_1_360_s_0_270=9.72e-05 mcm3l1d_cc_w_1_360_s_0_270=6.92e-11 mcm3l1d_cf_w_1_360_s_0_270=1.09e-11
+  mcm3l1d_ca_w_1_360_s_0_360=9.72e-05 mcm3l1d_cc_w_1_360_s_0_360=5.23e-11 mcm3l1d_cf_w_1_360_s_0_360=1.46e-11
+  mcm3l1d_ca_w_1_360_s_0_450=9.72e-05 mcm3l1d_cc_w_1_360_s_0_450=4.14e-11 mcm3l1d_cf_w_1_360_s_0_450=1.81e-11
+  mcm3l1d_ca_w_1_360_s_0_540=9.72e-05 mcm3l1d_cc_w_1_360_s_0_540=3.37e-11 mcm3l1d_cf_w_1_360_s_0_540=2.13e-11
+  mcm3l1d_ca_w_1_360_s_0_720=9.72e-05 mcm3l1d_cc_w_1_360_s_0_720=2.35e-11 mcm3l1d_cf_w_1_360_s_0_720=2.67e-11
+  mcm3l1d_ca_w_1_360_s_1_080=9.72e-05 mcm3l1d_cc_w_1_360_s_1_080=1.23e-11 mcm3l1d_cf_w_1_360_s_1_080=3.44e-11
+  mcm3l1d_ca_w_1_360_s_1_980=9.72e-05 mcm3l1d_cc_w_1_360_s_1_980=2.82e-12 mcm3l1d_cf_w_1_360_s_1_980=4.27e-11
+  mcm3l1d_ca_w_1_360_s_4_500=9.72e-05 mcm3l1d_cc_w_1_360_s_4_500=1.05e-13 mcm3l1d_cf_w_1_360_s_4_500=4.53e-11
+  mcm3l1p1_ca_w_0_170_s_0_180=2.01e-04 mcm3l1p1_cc_w_0_170_s_0_180=8.68e-11 mcm3l1p1_cf_w_0_170_s_0_180=1.38e-11
+  mcm3l1p1_ca_w_0_170_s_0_225=2.01e-04 mcm3l1p1_cc_w_0_170_s_0_225=6.71e-11 mcm3l1p1_cf_w_0_170_s_0_225=1.75e-11
+  mcm3l1p1_ca_w_0_170_s_0_270=2.01e-04 mcm3l1p1_cc_w_0_170_s_0_270=5.45e-11 mcm3l1p1_cf_w_0_170_s_0_270=2.10e-11
+  mcm3l1p1_ca_w_0_170_s_0_360=2.01e-04 mcm3l1p1_cc_w_0_170_s_0_360=3.85e-11 mcm3l1p1_cf_w_0_170_s_0_360=2.73e-11
+  mcm3l1p1_ca_w_0_170_s_0_450=2.01e-04 mcm3l1p1_cc_w_0_170_s_0_450=2.87e-11 mcm3l1p1_cf_w_0_170_s_0_450=3.25e-11
+  mcm3l1p1_ca_w_0_170_s_0_540=2.01e-04 mcm3l1p1_cc_w_0_170_s_0_540=2.19e-11 mcm3l1p1_cf_w_0_170_s_0_540=3.69e-11
+  mcm3l1p1_ca_w_0_170_s_0_720=2.01e-04 mcm3l1p1_cc_w_0_170_s_0_720=1.34e-11 mcm3l1p1_cf_w_0_170_s_0_720=4.32e-11
+  mcm3l1p1_ca_w_0_170_s_1_080=2.01e-04 mcm3l1p1_cc_w_0_170_s_1_080=5.63e-12 mcm3l1p1_cf_w_0_170_s_1_080=4.99e-11
+  mcm3l1p1_ca_w_0_170_s_1_980=2.01e-04 mcm3l1p1_cc_w_0_170_s_1_980=8.85e-13 mcm3l1p1_cf_w_0_170_s_1_980=5.44e-11
+  mcm3l1p1_ca_w_0_170_s_4_500=2.01e-04 mcm3l1p1_cc_w_0_170_s_4_500=4.50e-14 mcm3l1p1_cf_w_0_170_s_4_500=5.53e-11
+  mcm3l1p1_ca_w_1_360_s_0_180=2.01e-04 mcm3l1p1_cc_w_1_360_s_0_180=9.37e-11 mcm3l1p1_cf_w_1_360_s_0_180=1.38e-11
+  mcm3l1p1_ca_w_1_360_s_0_225=2.01e-04 mcm3l1p1_cc_w_1_360_s_0_225=7.34e-11 mcm3l1p1_cf_w_1_360_s_0_225=1.75e-11
+  mcm3l1p1_ca_w_1_360_s_0_270=2.01e-04 mcm3l1p1_cc_w_1_360_s_0_270=6.01e-11 mcm3l1p1_cf_w_1_360_s_0_270=2.10e-11
+  mcm3l1p1_ca_w_1_360_s_0_360=2.01e-04 mcm3l1p1_cc_w_1_360_s_0_360=4.33e-11 mcm3l1p1_cf_w_1_360_s_0_360=2.73e-11
+  mcm3l1p1_ca_w_1_360_s_0_450=2.01e-04 mcm3l1p1_cc_w_1_360_s_0_450=3.27e-11 mcm3l1p1_cf_w_1_360_s_0_450=3.26e-11
+  mcm3l1p1_ca_w_1_360_s_0_540=2.01e-04 mcm3l1p1_cc_w_1_360_s_0_540=2.54e-11 mcm3l1p1_cf_w_1_360_s_0_540=3.71e-11
+  mcm3l1p1_ca_w_1_360_s_0_720=2.01e-04 mcm3l1p1_cc_w_1_360_s_0_720=1.61e-11 mcm3l1p1_cf_w_1_360_s_0_720=4.37e-11
+  mcm3l1p1_ca_w_1_360_s_1_080=2.01e-04 mcm3l1p1_cc_w_1_360_s_1_080=7.15e-12 mcm3l1p1_cf_w_1_360_s_1_080=5.13e-11
+  mcm3l1p1_ca_w_1_360_s_1_980=2.01e-04 mcm3l1p1_cc_w_1_360_s_1_980=1.19e-12 mcm3l1p1_cf_w_1_360_s_1_980=5.70e-11
+  mcm3l1p1_ca_w_1_360_s_4_500=2.01e-04 mcm3l1p1_cc_w_1_360_s_4_500=4.00e-14 mcm3l1p1_cf_w_1_360_s_4_500=5.81e-11
+  mcm4l1f_ca_w_0_170_s_0_180=6.40e-05 mcm4l1f_cc_w_0_170_s_0_180=9.89e-11 mcm4l1f_cf_w_0_170_s_0_180=4.60e-12
+  mcm4l1f_ca_w_0_170_s_0_225=6.40e-05 mcm4l1f_cc_w_0_170_s_0_225=7.99e-11 mcm4l1f_cf_w_0_170_s_0_225=5.96e-12
+  mcm4l1f_ca_w_0_170_s_0_270=6.40e-05 mcm4l1f_cc_w_0_170_s_0_270=6.78e-11 mcm4l1f_cf_w_0_170_s_0_270=7.29e-12
+  mcm4l1f_ca_w_0_170_s_0_360=6.40e-05 mcm4l1f_cc_w_0_170_s_0_360=5.25e-11 mcm4l1f_cf_w_0_170_s_0_360=9.95e-12
+  mcm4l1f_ca_w_0_170_s_0_450=6.40e-05 mcm4l1f_cc_w_0_170_s_0_450=4.30e-11 mcm4l1f_cf_w_0_170_s_0_450=1.23e-11
+  mcm4l1f_ca_w_0_170_s_0_540=6.40e-05 mcm4l1f_cc_w_0_170_s_0_540=3.60e-11 mcm4l1f_cf_w_0_170_s_0_540=1.48e-11
+  mcm4l1f_ca_w_0_170_s_0_720=6.40e-05 mcm4l1f_cc_w_0_170_s_0_720=2.67e-11 mcm4l1f_cf_w_0_170_s_0_720=1.88e-11
+  mcm4l1f_ca_w_0_170_s_1_080=6.40e-05 mcm4l1f_cc_w_0_170_s_1_080=1.61e-11 mcm4l1f_cf_w_0_170_s_1_080=2.52e-11
+  mcm4l1f_ca_w_0_170_s_1_980=6.40e-05 mcm4l1f_cc_w_0_170_s_1_980=5.52e-12 mcm4l1f_cf_w_0_170_s_1_980=3.35e-11
+  mcm4l1f_ca_w_0_170_s_4_500=6.40e-05 mcm4l1f_cc_w_0_170_s_4_500=4.45e-13 mcm4l1f_cf_w_0_170_s_4_500=3.83e-11
+  mcm4l1f_ca_w_1_360_s_0_180=6.40e-05 mcm4l1f_cc_w_1_360_s_0_180=1.12e-10 mcm4l1f_cf_w_1_360_s_0_180=4.59e-12
+  mcm4l1f_ca_w_1_360_s_0_225=6.40e-05 mcm4l1f_cc_w_1_360_s_0_225=9.19e-11 mcm4l1f_cf_w_1_360_s_0_225=5.96e-12
+  mcm4l1f_ca_w_1_360_s_0_270=6.40e-05 mcm4l1f_cc_w_1_360_s_0_270=7.85e-11 mcm4l1f_cf_w_1_360_s_0_270=7.30e-12
+  mcm4l1f_ca_w_1_360_s_0_360=6.40e-05 mcm4l1f_cc_w_1_360_s_0_360=6.17e-11 mcm4l1f_cf_w_1_360_s_0_360=9.90e-12
+  mcm4l1f_ca_w_1_360_s_0_450=6.40e-05 mcm4l1f_cc_w_1_360_s_0_450=5.09e-11 mcm4l1f_cf_w_1_360_s_0_450=1.24e-11
+  mcm4l1f_ca_w_1_360_s_0_540=6.40e-05 mcm4l1f_cc_w_1_360_s_0_540=4.31e-11 mcm4l1f_cf_w_1_360_s_0_540=1.47e-11
+  mcm4l1f_ca_w_1_360_s_0_720=6.40e-05 mcm4l1f_cc_w_1_360_s_0_720=3.25e-11 mcm4l1f_cf_w_1_360_s_0_720=1.89e-11
+  mcm4l1f_ca_w_1_360_s_1_080=6.40e-05 mcm4l1f_cc_w_1_360_s_1_080=2.02e-11 mcm4l1f_cf_w_1_360_s_1_080=2.58e-11
+  mcm4l1f_ca_w_1_360_s_1_980=6.40e-05 mcm4l1f_cc_w_1_360_s_1_980=7.37e-12 mcm4l1f_cf_w_1_360_s_1_980=3.55e-11
+  mcm4l1f_ca_w_1_360_s_4_500=6.40e-05 mcm4l1f_cc_w_1_360_s_4_500=6.20e-13 mcm4l1f_cf_w_1_360_s_4_500=4.18e-11
+  mcm4l1d_ca_w_0_170_s_0_180=8.52e-05 mcm4l1d_cc_w_0_170_s_0_180=9.64e-11 mcm4l1d_cf_w_0_170_s_0_180=6.07e-12
+  mcm4l1d_ca_w_0_170_s_0_225=8.52e-05 mcm4l1d_cc_w_0_170_s_0_225=7.71e-11 mcm4l1d_cf_w_0_170_s_0_225=7.85e-12
+  mcm4l1d_ca_w_0_170_s_0_270=8.52e-05 mcm4l1d_cc_w_0_170_s_0_270=6.50e-11 mcm4l1d_cf_w_0_170_s_0_270=9.58e-12
+  mcm4l1d_ca_w_0_170_s_0_360=8.52e-05 mcm4l1d_cc_w_0_170_s_0_360=4.94e-11 mcm4l1d_cf_w_0_170_s_0_360=1.30e-11
+  mcm4l1d_ca_w_0_170_s_0_450=8.52e-05 mcm4l1d_cc_w_0_170_s_0_450=3.98e-11 mcm4l1d_cf_w_0_170_s_0_450=1.59e-11
+  mcm4l1d_ca_w_0_170_s_0_540=8.52e-05 mcm4l1d_cc_w_0_170_s_0_540=3.27e-11 mcm4l1d_cf_w_0_170_s_0_540=1.89e-11
+  mcm4l1d_ca_w_0_170_s_0_720=8.52e-05 mcm4l1d_cc_w_0_170_s_0_720=2.35e-11 mcm4l1d_cf_w_0_170_s_0_720=2.37e-11
+  mcm4l1d_ca_w_0_170_s_1_080=8.52e-05 mcm4l1d_cc_w_0_170_s_1_080=1.33e-11 mcm4l1d_cf_w_0_170_s_1_080=3.07e-11
+  mcm4l1d_ca_w_0_170_s_1_980=8.52e-05 mcm4l1d_cc_w_0_170_s_1_980=4.01e-12 mcm4l1d_cf_w_0_170_s_1_980=3.85e-11
+  mcm4l1d_ca_w_0_170_s_4_500=8.52e-05 mcm4l1d_cc_w_0_170_s_4_500=2.95e-13 mcm4l1d_cf_w_0_170_s_4_500=4.21e-11
+  mcm4l1d_ca_w_1_360_s_0_180=8.52e-05 mcm4l1d_cc_w_1_360_s_0_180=1.08e-10 mcm4l1d_cf_w_1_360_s_0_180=6.06e-12
+  mcm4l1d_ca_w_1_360_s_0_225=8.52e-05 mcm4l1d_cc_w_1_360_s_0_225=8.80e-11 mcm4l1d_cf_w_1_360_s_0_225=7.85e-12
+  mcm4l1d_ca_w_1_360_s_0_270=8.52e-05 mcm4l1d_cc_w_1_360_s_0_270=7.47e-11 mcm4l1d_cf_w_1_360_s_0_270=9.58e-12
+  mcm4l1d_ca_w_1_360_s_0_360=8.52e-05 mcm4l1d_cc_w_1_360_s_0_360=5.78e-11 mcm4l1d_cf_w_1_360_s_0_360=1.29e-11
+  mcm4l1d_ca_w_1_360_s_0_450=8.52e-05 mcm4l1d_cc_w_1_360_s_0_450=4.70e-11 mcm4l1d_cf_w_1_360_s_0_450=1.60e-11
+  mcm4l1d_ca_w_1_360_s_0_540=8.52e-05 mcm4l1d_cc_w_1_360_s_0_540=3.94e-11 mcm4l1d_cf_w_1_360_s_0_540=1.89e-11
+  mcm4l1d_ca_w_1_360_s_0_720=8.52e-05 mcm4l1d_cc_w_1_360_s_0_720=2.89e-11 mcm4l1d_cf_w_1_360_s_0_720=2.39e-11
+  mcm4l1d_ca_w_1_360_s_1_080=8.52e-05 mcm4l1d_cc_w_1_360_s_1_080=1.71e-11 mcm4l1d_cf_w_1_360_s_1_080=3.14e-11
+  mcm4l1d_ca_w_1_360_s_1_980=8.52e-05 mcm4l1d_cc_w_1_360_s_1_980=5.64e-12 mcm4l1d_cf_w_1_360_s_1_980=4.09e-11
+  mcm4l1d_ca_w_1_360_s_4_500=8.52e-05 mcm4l1d_cc_w_1_360_s_4_500=3.95e-13 mcm4l1d_cf_w_1_360_s_4_500=4.59e-11
+  mcm4l1p1_ca_w_0_170_s_0_180=1.88e-04 mcm4l1p1_cc_w_0_170_s_0_180=8.85e-11 mcm4l1p1_cf_w_0_170_s_0_180=1.29e-11
+  mcm4l1p1_ca_w_0_170_s_0_225=1.88e-04 mcm4l1p1_cc_w_0_170_s_0_225=6.90e-11 mcm4l1p1_cf_w_0_170_s_0_225=1.65e-11
+  mcm4l1p1_ca_w_0_170_s_0_270=1.88e-04 mcm4l1p1_cc_w_0_170_s_0_270=5.67e-11 mcm4l1p1_cf_w_0_170_s_0_270=1.97e-11
+  mcm4l1p1_ca_w_0_170_s_0_360=1.88e-04 mcm4l1p1_cc_w_0_170_s_0_360=4.07e-11 mcm4l1p1_cf_w_0_170_s_0_360=2.58e-11
+  mcm4l1p1_ca_w_0_170_s_0_450=1.88e-04 mcm4l1p1_cc_w_0_170_s_0_450=3.12e-11 mcm4l1p1_cf_w_0_170_s_0_450=3.07e-11
+  mcm4l1p1_ca_w_0_170_s_0_540=1.88e-04 mcm4l1p1_cc_w_0_170_s_0_540=2.42e-11 mcm4l1p1_cf_w_0_170_s_0_540=3.51e-11
+  mcm4l1p1_ca_w_0_170_s_0_720=1.88e-04 mcm4l1p1_cc_w_0_170_s_0_720=1.57e-11 mcm4l1p1_cf_w_0_170_s_0_720=4.13e-11
+  mcm4l1p1_ca_w_0_170_s_1_080=1.88e-04 mcm4l1p1_cc_w_0_170_s_1_080=7.48e-12 mcm4l1p1_cf_w_0_170_s_1_080=4.83e-11
+  mcm4l1p1_ca_w_0_170_s_1_980=1.88e-04 mcm4l1p1_cc_w_0_170_s_1_980=1.80e-12 mcm4l1p1_cf_w_0_170_s_1_980=5.36e-11
+  mcm4l1p1_ca_w_0_170_s_4_500=1.88e-04 mcm4l1p1_cc_w_0_170_s_4_500=1.30e-13 mcm4l1p1_cf_w_0_170_s_4_500=5.53e-11
+  mcm4l1p1_ca_w_1_360_s_0_180=1.88e-04 mcm4l1p1_cc_w_1_360_s_0_180=9.91e-11 mcm4l1p1_cf_w_1_360_s_0_180=1.31e-11
+  mcm4l1p1_ca_w_1_360_s_0_225=1.88e-04 mcm4l1p1_cc_w_1_360_s_0_225=7.89e-11 mcm4l1p1_cf_w_1_360_s_0_225=1.66e-11
+  mcm4l1p1_ca_w_1_360_s_0_270=1.88e-04 mcm4l1p1_cc_w_1_360_s_0_270=6.56e-11 mcm4l1p1_cf_w_1_360_s_0_270=1.99e-11
+  mcm4l1p1_ca_w_1_360_s_0_360=1.88e-04 mcm4l1p1_cc_w_1_360_s_0_360=4.88e-11 mcm4l1p1_cf_w_1_360_s_0_360=2.58e-11
+  mcm4l1p1_ca_w_1_360_s_0_450=1.88e-04 mcm4l1p1_cc_w_1_360_s_0_450=3.81e-11 mcm4l1p1_cf_w_1_360_s_0_450=3.09e-11
+  mcm4l1p1_ca_w_1_360_s_0_540=1.88e-04 mcm4l1p1_cc_w_1_360_s_0_540=3.08e-11 mcm4l1p1_cf_w_1_360_s_0_540=3.52e-11
+  mcm4l1p1_ca_w_1_360_s_0_720=1.88e-04 mcm4l1p1_cc_w_1_360_s_0_720=2.11e-11 mcm4l1p1_cf_w_1_360_s_0_720=4.19e-11
+  mcm4l1p1_ca_w_1_360_s_1_080=1.88e-04 mcm4l1p1_cc_w_1_360_s_1_080=1.12e-11 mcm4l1p1_cf_w_1_360_s_1_080=5.00e-11
+  mcm4l1p1_ca_w_1_360_s_1_980=1.88e-04 mcm4l1p1_cc_w_1_360_s_1_980=3.18e-12 mcm4l1p1_cf_w_1_360_s_1_980=5.74e-11
+  mcm4l1p1_ca_w_1_360_s_4_500=1.88e-04 mcm4l1p1_cc_w_1_360_s_4_500=2.25e-13 mcm4l1p1_cf_w_1_360_s_4_500=6.03e-11
+  mcm5l1f_ca_w_0_170_s_0_180=5.92e-05 mcm5l1f_cc_w_0_170_s_0_180=9.96e-11 mcm5l1f_cf_w_0_170_s_0_180=4.25e-12
+  mcm5l1f_ca_w_0_170_s_0_225=5.92e-05 mcm5l1f_cc_w_0_170_s_0_225=8.06e-11 mcm5l1f_cf_w_0_170_s_0_225=5.52e-12
+  mcm5l1f_ca_w_0_170_s_0_270=5.92e-05 mcm5l1f_cc_w_0_170_s_0_270=6.87e-11 mcm5l1f_cf_w_0_170_s_0_270=6.75e-12
+  mcm5l1f_ca_w_0_170_s_0_360=5.92e-05 mcm5l1f_cc_w_0_170_s_0_360=5.34e-11 mcm5l1f_cf_w_0_170_s_0_360=9.21e-12
+  mcm5l1f_ca_w_0_170_s_0_450=5.92e-05 mcm5l1f_cc_w_0_170_s_0_450=4.42e-11 mcm5l1f_cf_w_0_170_s_0_450=1.14e-11
+  mcm5l1f_ca_w_0_170_s_0_540=5.92e-05 mcm5l1f_cc_w_0_170_s_0_540=3.72e-11 mcm5l1f_cf_w_0_170_s_0_540=1.38e-11
+  mcm5l1f_ca_w_0_170_s_0_720=5.92e-05 mcm5l1f_cc_w_0_170_s_0_720=2.81e-11 mcm5l1f_cf_w_0_170_s_0_720=1.76e-11
+  mcm5l1f_ca_w_0_170_s_1_080=5.92e-05 mcm5l1f_cc_w_0_170_s_1_080=1.76e-11 mcm5l1f_cf_w_0_170_s_1_080=2.38e-11
+  mcm5l1f_ca_w_0_170_s_1_980=5.92e-05 mcm5l1f_cc_w_0_170_s_1_980=6.80e-12 mcm5l1f_cf_w_0_170_s_1_980=3.21e-11
+  mcm5l1f_ca_w_0_170_s_4_500=5.92e-05 mcm5l1f_cc_w_0_170_s_4_500=8.45e-13 mcm5l1f_cf_w_0_170_s_4_500=3.76e-11
+  mcm5l1f_ca_w_1_360_s_0_180=5.92e-05 mcm5l1f_cc_w_1_360_s_0_180=1.15e-10 mcm5l1f_cf_w_1_360_s_0_180=4.25e-12
+  mcm5l1f_ca_w_1_360_s_0_225=5.92e-05 mcm5l1f_cc_w_1_360_s_0_225=9.46e-11 mcm5l1f_cf_w_1_360_s_0_225=5.51e-12
+  mcm5l1f_ca_w_1_360_s_0_270=5.92e-05 mcm5l1f_cc_w_1_360_s_0_270=8.14e-11 mcm5l1f_cf_w_1_360_s_0_270=6.76e-12
+  mcm5l1f_ca_w_1_360_s_0_360=5.92e-05 mcm5l1f_cc_w_1_360_s_0_360=6.46e-11 mcm5l1f_cf_w_1_360_s_0_360=9.17e-12
+  mcm5l1f_ca_w_1_360_s_0_450=5.92e-05 mcm5l1f_cc_w_1_360_s_0_450=5.38e-11 mcm5l1f_cf_w_1_360_s_0_450=1.15e-11
+  mcm5l1f_ca_w_1_360_s_0_540=5.92e-05 mcm5l1f_cc_w_1_360_s_0_540=4.61e-11 mcm5l1f_cf_w_1_360_s_0_540=1.37e-11
+  mcm5l1f_ca_w_1_360_s_0_720=5.92e-05 mcm5l1f_cc_w_1_360_s_0_720=3.56e-11 mcm5l1f_cf_w_1_360_s_0_720=1.76e-11
+  mcm5l1f_ca_w_1_360_s_1_080=5.92e-05 mcm5l1f_cc_w_1_360_s_1_080=2.32e-11 mcm5l1f_cf_w_1_360_s_1_080=2.42e-11
+  mcm5l1f_ca_w_1_360_s_1_980=5.92e-05 mcm5l1f_cc_w_1_360_s_1_980=9.77e-12 mcm5l1f_cf_w_1_360_s_1_980=3.41e-11
+  mcm5l1f_ca_w_1_360_s_4_500=5.92e-05 mcm5l1f_cc_w_1_360_s_4_500=1.39e-12 mcm5l1f_cf_w_1_360_s_4_500=4.18e-11
+  mcm5l1d_ca_w_0_170_s_0_180=8.04e-05 mcm5l1d_cc_w_0_170_s_0_180=9.71e-11 mcm5l1d_cf_w_0_170_s_0_180=5.73e-12
+  mcm5l1d_ca_w_0_170_s_0_225=8.04e-05 mcm5l1d_cc_w_0_170_s_0_225=7.79e-11 mcm5l1d_cf_w_0_170_s_0_225=7.41e-12
+  mcm5l1d_ca_w_0_170_s_0_270=8.04e-05 mcm5l1d_cc_w_0_170_s_0_270=6.59e-11 mcm5l1d_cf_w_0_170_s_0_270=9.04e-12
+  mcm5l1d_ca_w_0_170_s_0_360=8.04e-05 mcm5l1d_cc_w_0_170_s_0_360=5.03e-11 mcm5l1d_cf_w_0_170_s_0_360=1.23e-11
+  mcm5l1d_ca_w_0_170_s_0_450=8.04e-05 mcm5l1d_cc_w_0_170_s_0_450=4.10e-11 mcm5l1d_cf_w_0_170_s_0_450=1.51e-11
+  mcm5l1d_ca_w_0_170_s_0_540=8.04e-05 mcm5l1d_cc_w_0_170_s_0_540=3.39e-11 mcm5l1d_cf_w_0_170_s_0_540=1.79e-11
+  mcm5l1d_ca_w_0_170_s_0_720=8.04e-05 mcm5l1d_cc_w_0_170_s_0_720=2.47e-11 mcm5l1d_cf_w_0_170_s_0_720=2.26e-11
+  mcm5l1d_ca_w_0_170_s_1_080=8.04e-05 mcm5l1d_cc_w_0_170_s_1_080=1.46e-11 mcm5l1d_cf_w_0_170_s_1_080=2.95e-11
+  mcm5l1d_ca_w_0_170_s_1_980=8.04e-05 mcm5l1d_cc_w_0_170_s_1_980=5.03e-12 mcm5l1d_cf_w_0_170_s_1_980=3.74e-11
+  mcm5l1d_ca_w_0_170_s_4_500=8.04e-05 mcm5l1d_cc_w_0_170_s_4_500=5.70e-13 mcm5l1d_cf_w_0_170_s_4_500=4.17e-11
+  mcm5l1d_ca_w_1_360_s_0_180=8.04e-05 mcm5l1d_cc_w_1_360_s_0_180=1.11e-10 mcm5l1d_cf_w_1_360_s_0_180=5.72e-12
+  mcm5l1d_ca_w_1_360_s_0_225=8.04e-05 mcm5l1d_cc_w_1_360_s_0_225=9.07e-11 mcm5l1d_cf_w_1_360_s_0_225=7.40e-12
+  mcm5l1d_ca_w_1_360_s_0_270=8.04e-05 mcm5l1d_cc_w_1_360_s_0_270=7.75e-11 mcm5l1d_cf_w_1_360_s_0_270=9.04e-12
+  mcm5l1d_ca_w_1_360_s_0_360=8.04e-05 mcm5l1d_cc_w_1_360_s_0_360=6.07e-11 mcm5l1d_cf_w_1_360_s_0_360=1.22e-11
+  mcm5l1d_ca_w_1_360_s_0_450=8.04e-05 mcm5l1d_cc_w_1_360_s_0_450=4.99e-11 mcm5l1d_cf_w_1_360_s_0_450=1.51e-11
+  mcm5l1d_ca_w_1_360_s_0_540=8.04e-05 mcm5l1d_cc_w_1_360_s_0_540=4.23e-11 mcm5l1d_cf_w_1_360_s_0_540=1.79e-11
+  mcm5l1d_ca_w_1_360_s_0_720=8.04e-05 mcm5l1d_cc_w_1_360_s_0_720=3.19e-11 mcm5l1d_cf_w_1_360_s_0_720=2.27e-11
+  mcm5l1d_ca_w_1_360_s_1_080=8.04e-05 mcm5l1d_cc_w_1_360_s_1_080=2.00e-11 mcm5l1d_cf_w_1_360_s_1_080=3.01e-11
+  mcm5l1d_ca_w_1_360_s_1_980=8.04e-05 mcm5l1d_cc_w_1_360_s_1_980=7.81e-12 mcm5l1d_cf_w_1_360_s_1_980=4.00e-11
+  mcm5l1d_ca_w_1_360_s_4_500=8.04e-05 mcm5l1d_cc_w_1_360_s_4_500=9.95e-13 mcm5l1d_cf_w_1_360_s_4_500=4.64e-11
+  mcm5l1p1_ca_w_0_170_s_0_180=1.84e-04 mcm5l1p1_cc_w_0_170_s_0_180=8.92e-11 mcm5l1p1_cf_w_0_170_s_0_180=1.26e-11
+  mcm5l1p1_ca_w_0_170_s_0_225=1.84e-04 mcm5l1p1_cc_w_0_170_s_0_225=6.98e-11 mcm5l1p1_cf_w_0_170_s_0_225=1.60e-11
+  mcm5l1p1_ca_w_0_170_s_0_270=1.84e-04 mcm5l1p1_cc_w_0_170_s_0_270=5.75e-11 mcm5l1p1_cf_w_0_170_s_0_270=1.92e-11
+  mcm5l1p1_ca_w_0_170_s_0_360=1.84e-04 mcm5l1p1_cc_w_0_170_s_0_360=4.17e-11 mcm5l1p1_cf_w_0_170_s_0_360=2.52e-11
+  mcm5l1p1_ca_w_0_170_s_0_450=1.84e-04 mcm5l1p1_cc_w_0_170_s_0_450=3.23e-11 mcm5l1p1_cf_w_0_170_s_0_450=2.99e-11
+  mcm5l1p1_ca_w_0_170_s_0_540=1.84e-04 mcm5l1p1_cc_w_0_170_s_0_540=2.53e-11 mcm5l1p1_cf_w_0_170_s_0_540=3.44e-11
+  mcm5l1p1_ca_w_0_170_s_0_720=1.84e-04 mcm5l1p1_cc_w_0_170_s_0_720=1.67e-11 mcm5l1p1_cf_w_0_170_s_0_720=4.06e-11
+  mcm5l1p1_ca_w_0_170_s_1_080=1.84e-04 mcm5l1p1_cc_w_0_170_s_1_080=8.43e-12 mcm5l1p1_cf_w_0_170_s_1_080=4.76e-11
+  mcm5l1p1_ca_w_0_170_s_1_980=1.84e-04 mcm5l1p1_cc_w_0_170_s_1_980=2.40e-12 mcm5l1p1_cf_w_0_170_s_1_980=5.32e-11
+  mcm5l1p1_ca_w_0_170_s_4_500=1.84e-04 mcm5l1p1_cc_w_0_170_s_4_500=2.50e-13 mcm5l1p1_cf_w_0_170_s_4_500=5.53e-11
+  mcm5l1p1_ca_w_1_360_s_0_180=1.84e-04 mcm5l1p1_cc_w_1_360_s_0_180=1.02e-10 mcm5l1p1_cf_w_1_360_s_0_180=1.28e-11
+  mcm5l1p1_ca_w_1_360_s_0_225=1.84e-04 mcm5l1p1_cc_w_1_360_s_0_225=8.16e-11 mcm5l1p1_cf_w_1_360_s_0_225=1.62e-11
+  mcm5l1p1_ca_w_1_360_s_0_270=1.84e-04 mcm5l1p1_cc_w_1_360_s_0_270=6.84e-11 mcm5l1p1_cf_w_1_360_s_0_270=1.94e-11
+  mcm5l1p1_ca_w_1_360_s_0_360=1.84e-04 mcm5l1p1_cc_w_1_360_s_0_360=5.16e-11 mcm5l1p1_cf_w_1_360_s_0_360=2.52e-11
+  mcm5l1p1_ca_w_1_360_s_0_450=1.84e-04 mcm5l1p1_cc_w_1_360_s_0_450=4.09e-11 mcm5l1p1_cf_w_1_360_s_0_450=3.02e-11
+  mcm5l1p1_ca_w_1_360_s_0_540=1.84e-04 mcm5l1p1_cc_w_1_360_s_0_540=3.37e-11 mcm5l1p1_cf_w_1_360_s_0_540=3.45e-11
+  mcm5l1p1_ca_w_1_360_s_0_720=1.84e-04 mcm5l1p1_cc_w_1_360_s_0_720=2.39e-11 mcm5l1p1_cf_w_1_360_s_0_720=4.11e-11
+  mcm5l1p1_ca_w_1_360_s_1_080=1.84e-04 mcm5l1p1_cc_w_1_360_s_1_080=1.37e-11 mcm5l1p1_cf_w_1_360_s_1_080=4.93e-11
+  mcm5l1p1_ca_w_1_360_s_1_980=1.84e-04 mcm5l1p1_cc_w_1_360_s_1_980=4.75e-12 mcm5l1p1_cf_w_1_360_s_1_980=5.75e-11
+  mcm5l1p1_ca_w_1_360_s_4_500=1.84e-04 mcm5l1p1_cc_w_1_360_s_4_500=5.50e-13 mcm5l1p1_cf_w_1_360_s_4_500=6.15e-11
+  mcrdll1f_ca_w_0_170_s_0_180=5.35e-05 mcrdll1f_cc_w_0_170_s_0_180=1.00e-10 mcrdll1f_cf_w_0_170_s_0_180=3.84e-12
+  mcrdll1f_ca_w_0_170_s_0_225=5.35e-05 mcrdll1f_cc_w_0_170_s_0_225=8.15e-11 mcrdll1f_cf_w_0_170_s_0_225=4.98e-12
+  mcrdll1f_ca_w_0_170_s_0_270=5.35e-05 mcrdll1f_cc_w_0_170_s_0_270=6.98e-11 mcrdll1f_cf_w_0_170_s_0_270=6.10e-12
+  mcrdll1f_ca_w_0_170_s_0_360=5.35e-05 mcrdll1f_cc_w_0_170_s_0_360=5.46e-11 mcrdll1f_cf_w_0_170_s_0_360=8.33e-12
+  mcrdll1f_ca_w_0_170_s_0_450=5.35e-05 mcrdll1f_cc_w_0_170_s_0_450=4.56e-11 mcrdll1f_cf_w_0_170_s_0_450=1.03e-11
+  mcrdll1f_ca_w_0_170_s_0_540=5.35e-05 mcrdll1f_cc_w_0_170_s_0_540=3.87e-11 mcrdll1f_cf_w_0_170_s_0_540=1.25e-11
+  mcrdll1f_ca_w_0_170_s_0_720=5.35e-05 mcrdll1f_cc_w_0_170_s_0_720=2.98e-11 mcrdll1f_cf_w_0_170_s_0_720=1.61e-11
+  mcrdll1f_ca_w_0_170_s_1_080=5.35e-05 mcrdll1f_cc_w_0_170_s_1_080=1.95e-11 mcrdll1f_cf_w_0_170_s_1_080=2.20e-11
+  mcrdll1f_ca_w_0_170_s_1_980=5.35e-05 mcrdll1f_cc_w_0_170_s_1_980=8.80e-12 mcrdll1f_cf_w_0_170_s_1_980=3.02e-11
+  mcrdll1f_ca_w_0_170_s_4_500=5.35e-05 mcrdll1f_cc_w_0_170_s_4_500=1.81e-12 mcrdll1f_cf_w_0_170_s_4_500=3.66e-11
+  mcrdll1f_ca_w_1_360_s_0_180=5.35e-05 mcrdll1f_cc_w_1_360_s_0_180=1.18e-10 mcrdll1f_cf_w_1_360_s_0_180=3.84e-12
+  mcrdll1f_ca_w_1_360_s_0_225=5.35e-05 mcrdll1f_cc_w_1_360_s_0_225=9.83e-11 mcrdll1f_cf_w_1_360_s_0_225=4.98e-12
+  mcrdll1f_ca_w_1_360_s_0_270=5.35e-05 mcrdll1f_cc_w_1_360_s_0_270=8.51e-11 mcrdll1f_cf_w_1_360_s_0_270=6.11e-12
+  mcrdll1f_ca_w_1_360_s_0_360=5.35e-05 mcrdll1f_cc_w_1_360_s_0_360=6.84e-11 mcrdll1f_cf_w_1_360_s_0_360=8.29e-12
+  mcrdll1f_ca_w_1_360_s_0_450=5.35e-05 mcrdll1f_cc_w_1_360_s_0_450=5.78e-11 mcrdll1f_cf_w_1_360_s_0_450=1.04e-11
+  mcrdll1f_ca_w_1_360_s_0_540=5.35e-05 mcrdll1f_cc_w_1_360_s_0_540=5.03e-11 mcrdll1f_cf_w_1_360_s_0_540=1.24e-11
+  mcrdll1f_ca_w_1_360_s_0_720=5.35e-05 mcrdll1f_cc_w_1_360_s_0_720=3.99e-11 mcrdll1f_cf_w_1_360_s_0_720=1.60e-11
+  mcrdll1f_ca_w_1_360_s_1_080=5.35e-05 mcrdll1f_cc_w_1_360_s_1_080=2.78e-11 mcrdll1f_cf_w_1_360_s_1_080=2.22e-11
+  mcrdll1f_ca_w_1_360_s_1_980=5.35e-05 mcrdll1f_cc_w_1_360_s_1_980=1.39e-11 mcrdll1f_cf_w_1_360_s_1_980=3.21e-11
+  mcrdll1f_ca_w_1_360_s_4_500=5.35e-05 mcrdll1f_cc_w_1_360_s_4_500=3.60e-12 mcrdll1f_cf_w_1_360_s_4_500=4.15e-11
+  mcrdll1d_ca_w_0_170_s_0_180=7.47e-05 mcrdll1d_cc_w_0_170_s_0_180=9.78e-11 mcrdll1d_cf_w_0_170_s_0_180=5.32e-12
+  mcrdll1d_ca_w_0_170_s_0_225=7.47e-05 mcrdll1d_cc_w_0_170_s_0_225=7.88e-11 mcrdll1d_cf_w_0_170_s_0_225=6.88e-12
+  mcrdll1d_ca_w_0_170_s_0_270=7.47e-05 mcrdll1d_cc_w_0_170_s_0_270=6.68e-11 mcrdll1d_cf_w_0_170_s_0_270=8.38e-12
+  mcrdll1d_ca_w_0_170_s_0_360=7.47e-05 mcrdll1d_cc_w_0_170_s_0_360=5.15e-11 mcrdll1d_cf_w_0_170_s_0_360=1.14e-11
+  mcrdll1d_ca_w_0_170_s_0_450=7.47e-05 mcrdll1d_cc_w_0_170_s_0_450=4.23e-11 mcrdll1d_cf_w_0_170_s_0_450=1.40e-11
+  mcrdll1d_ca_w_0_170_s_0_540=7.47e-05 mcrdll1d_cc_w_0_170_s_0_540=3.53e-11 mcrdll1d_cf_w_0_170_s_0_540=1.68e-11
+  mcrdll1d_ca_w_0_170_s_0_720=7.47e-05 mcrdll1d_cc_w_0_170_s_0_720=2.63e-11 mcrdll1d_cf_w_0_170_s_0_720=2.13e-11
+  mcrdll1d_ca_w_0_170_s_1_080=7.47e-05 mcrdll1d_cc_w_0_170_s_1_080=1.63e-11 mcrdll1d_cf_w_0_170_s_1_080=2.79e-11
+  mcrdll1d_ca_w_0_170_s_1_980=7.47e-05 mcrdll1d_cc_w_0_170_s_1_980=6.66e-12 mcrdll1d_cf_w_0_170_s_1_980=3.60e-11
+  mcrdll1d_ca_w_0_170_s_4_500=7.47e-05 mcrdll1d_cc_w_0_170_s_4_500=1.26e-12 mcrdll1d_cf_w_0_170_s_4_500=4.11e-11
+  mcrdll1d_ca_w_1_360_s_0_180=7.47e-05 mcrdll1d_cc_w_1_360_s_0_180=1.14e-10 mcrdll1d_cf_w_1_360_s_0_180=5.32e-12
+  mcrdll1d_ca_w_1_360_s_0_225=7.47e-05 mcrdll1d_cc_w_1_360_s_0_225=9.43e-11 mcrdll1d_cf_w_1_360_s_0_225=6.88e-12
+  mcrdll1d_ca_w_1_360_s_0_270=7.47e-05 mcrdll1d_cc_w_1_360_s_0_270=8.12e-11 mcrdll1d_cf_w_1_360_s_0_270=8.40e-12
+  mcrdll1d_ca_w_1_360_s_0_360=7.47e-05 mcrdll1d_cc_w_1_360_s_0_360=6.46e-11 mcrdll1d_cf_w_1_360_s_0_360=1.13e-11
+  mcrdll1d_ca_w_1_360_s_0_450=7.47e-05 mcrdll1d_cc_w_1_360_s_0_450=5.39e-11 mcrdll1d_cf_w_1_360_s_0_450=1.41e-11
+  mcrdll1d_ca_w_1_360_s_0_540=7.47e-05 mcrdll1d_cc_w_1_360_s_0_540=4.65e-11 mcrdll1d_cf_w_1_360_s_0_540=1.66e-11
+  mcrdll1d_ca_w_1_360_s_0_720=7.47e-05 mcrdll1d_cc_w_1_360_s_0_720=3.61e-11 mcrdll1d_cf_w_1_360_s_0_720=2.12e-11
+  mcrdll1d_ca_w_1_360_s_1_080=7.47e-05 mcrdll1d_cc_w_1_360_s_1_080=2.43e-11 mcrdll1d_cf_w_1_360_s_1_080=2.83e-11
+  mcrdll1d_ca_w_1_360_s_1_980=7.47e-05 mcrdll1d_cc_w_1_360_s_1_980=1.15e-11 mcrdll1d_cf_w_1_360_s_1_980=3.86e-11
+  mcrdll1d_ca_w_1_360_s_4_500=7.47e-05 mcrdll1d_cc_w_1_360_s_4_500=2.77e-12 mcrdll1d_cf_w_1_360_s_4_500=4.67e-11
+  mcrdll1p1_ca_w_0_170_s_0_180=1.78e-04 mcrdll1p1_cc_w_0_170_s_0_180=8.99e-11 mcrdll1p1_cf_w_0_170_s_0_180=1.22e-11
+  mcrdll1p1_ca_w_0_170_s_0_225=1.78e-04 mcrdll1p1_cc_w_0_170_s_0_225=7.06e-11 mcrdll1p1_cf_w_0_170_s_0_225=1.55e-11
+  mcrdll1p1_ca_w_0_170_s_0_270=1.78e-04 mcrdll1p1_cc_w_0_170_s_0_270=5.86e-11 mcrdll1p1_cf_w_0_170_s_0_270=1.85e-11
+  mcrdll1p1_ca_w_0_170_s_0_360=1.78e-04 mcrdll1p1_cc_w_0_170_s_0_360=4.28e-11 mcrdll1p1_cf_w_0_170_s_0_360=2.43e-11
+  mcrdll1p1_ca_w_0_170_s_0_450=1.78e-04 mcrdll1p1_cc_w_0_170_s_0_450=3.36e-11 mcrdll1p1_cf_w_0_170_s_0_450=2.89e-11
+  mcrdll1p1_ca_w_0_170_s_0_540=1.78e-04 mcrdll1p1_cc_w_0_170_s_0_540=2.65e-11 mcrdll1p1_cf_w_0_170_s_0_540=3.34e-11
+  mcrdll1p1_ca_w_0_170_s_0_720=1.78e-04 mcrdll1p1_cc_w_0_170_s_0_720=1.80e-11 mcrdll1p1_cf_w_0_170_s_0_720=3.95e-11
+  mcrdll1p1_ca_w_0_170_s_1_080=1.78e-04 mcrdll1p1_cc_w_0_170_s_1_080=9.57e-12 mcrdll1p1_cf_w_0_170_s_1_080=4.67e-11
+  mcrdll1p1_ca_w_0_170_s_1_980=1.78e-04 mcrdll1p1_cc_w_0_170_s_1_980=3.29e-12 mcrdll1p1_cf_w_0_170_s_1_980=5.26e-11
+  mcrdll1p1_ca_w_0_170_s_4_500=1.78e-04 mcrdll1p1_cc_w_0_170_s_4_500=6.15e-13 mcrdll1p1_cf_w_0_170_s_4_500=5.52e-11
+  mcrdll1p1_ca_w_1_360_s_0_180=1.78e-04 mcrdll1p1_cc_w_1_360_s_0_180=1.05e-10 mcrdll1p1_cf_w_1_360_s_0_180=1.24e-11
+  mcrdll1p1_ca_w_1_360_s_0_225=1.78e-04 mcrdll1p1_cc_w_1_360_s_0_225=8.53e-11 mcrdll1p1_cf_w_1_360_s_0_225=1.57e-11
+  mcrdll1p1_ca_w_1_360_s_0_270=1.78e-04 mcrdll1p1_cc_w_1_360_s_0_270=7.22e-11 mcrdll1p1_cf_w_1_360_s_0_270=1.88e-11
+  mcrdll1p1_ca_w_1_360_s_0_360=1.78e-04 mcrdll1p1_cc_w_1_360_s_0_360=5.54e-11 mcrdll1p1_cf_w_1_360_s_0_360=2.44e-11
+  mcrdll1p1_ca_w_1_360_s_0_450=1.78e-04 mcrdll1p1_cc_w_1_360_s_0_450=4.50e-11 mcrdll1p1_cf_w_1_360_s_0_450=2.92e-11
+  mcrdll1p1_ca_w_1_360_s_0_540=1.78e-04 mcrdll1p1_cc_w_1_360_s_0_540=3.76e-11 mcrdll1p1_cf_w_1_360_s_0_540=3.34e-11
+  mcrdll1p1_ca_w_1_360_s_0_720=1.78e-04 mcrdll1p1_cc_w_1_360_s_0_720=2.78e-11 mcrdll1p1_cf_w_1_360_s_0_720=4.00e-11
+  mcrdll1p1_ca_w_1_360_s_1_080=1.78e-04 mcrdll1p1_cc_w_1_360_s_1_080=1.74e-11 mcrdll1p1_cf_w_1_360_s_1_080=4.83e-11
+  mcrdll1p1_ca_w_1_360_s_1_980=1.78e-04 mcrdll1p1_cc_w_1_360_s_1_980=7.57e-12 mcrdll1p1_cf_w_1_360_s_1_980=5.74e-11
+  mcrdll1p1_ca_w_1_360_s_4_500=1.78e-04 mcrdll1p1_cc_w_1_360_s_4_500=1.74e-12 mcrdll1p1_cf_w_1_360_s_4_500=6.29e-11
+  mcm2m1f_ca_w_0_140_s_0_140=3.49e-04 mcm2m1f_cc_w_0_140_s_0_140=1.08e-10 mcm2m1f_cf_w_0_140_s_0_140=1.58e-11
+  mcm2m1f_ca_w_0_140_s_0_175=3.49e-04 mcm2m1f_cc_w_0_140_s_0_175=1.02e-10 mcm2m1f_cf_w_0_140_s_0_175=2.01e-11
+  mcm2m1f_ca_w_0_140_s_0_210=3.49e-04 mcm2m1f_cc_w_0_140_s_0_210=9.42e-11 mcm2m1f_cf_w_0_140_s_0_210=2.39e-11
+  mcm2m1f_ca_w_0_140_s_0_280=3.49e-04 mcm2m1f_cc_w_0_140_s_0_280=7.66e-11 mcm2m1f_cf_w_0_140_s_0_280=3.08e-11
+  mcm2m1f_ca_w_0_140_s_0_350=3.49e-04 mcm2m1f_cc_w_0_140_s_0_350=6.16e-11 mcm2m1f_cf_w_0_140_s_0_350=3.69e-11
+  mcm2m1f_ca_w_0_140_s_0_420=3.49e-04 mcm2m1f_cc_w_0_140_s_0_420=4.89e-11 mcm2m1f_cf_w_0_140_s_0_420=4.25e-11
+  mcm2m1f_ca_w_0_140_s_0_560=3.49e-04 mcm2m1f_cc_w_0_140_s_0_560=3.25e-11 mcm2m1f_cf_w_0_140_s_0_560=5.10e-11
+  mcm2m1f_ca_w_0_140_s_0_840=3.49e-04 mcm2m1f_cc_w_0_140_s_0_840=1.62e-11 mcm2m1f_cf_w_0_140_s_0_840=6.25e-11
+  mcm2m1f_ca_w_0_140_s_1_540=3.49e-04 mcm2m1f_cc_w_0_140_s_1_540=3.68e-12 mcm2m1f_cf_w_0_140_s_1_540=7.39e-11
+  mcm2m1f_ca_w_0_140_s_3_500=3.49e-04 mcm2m1f_cc_w_0_140_s_3_500=1.60e-13 mcm2m1f_cf_w_0_140_s_3_500=7.78e-11
+  mcm2m1f_ca_w_1_120_s_0_140=3.49e-04 mcm2m1f_cc_w_1_120_s_0_140=1.15e-10 mcm2m1f_cf_w_1_120_s_0_140=1.58e-11
+  mcm2m1f_ca_w_1_120_s_0_175=3.49e-04 mcm2m1f_cc_w_1_120_s_0_175=1.09e-10 mcm2m1f_cf_w_1_120_s_0_175=2.01e-11
+  mcm2m1f_ca_w_1_120_s_0_210=3.49e-04 mcm2m1f_cc_w_1_120_s_0_210=9.97e-11 mcm2m1f_cf_w_1_120_s_0_210=2.39e-11
+  mcm2m1f_ca_w_1_120_s_0_280=3.49e-04 mcm2m1f_cc_w_1_120_s_0_280=8.09e-11 mcm2m1f_cf_w_1_120_s_0_280=3.08e-11
+  mcm2m1f_ca_w_1_120_s_0_350=3.49e-04 mcm2m1f_cc_w_1_120_s_0_350=6.56e-11 mcm2m1f_cf_w_1_120_s_0_350=3.69e-11
+  mcm2m1f_ca_w_1_120_s_0_420=3.49e-04 mcm2m1f_cc_w_1_120_s_0_420=5.23e-11 mcm2m1f_cf_w_1_120_s_0_420=4.25e-11
+  mcm2m1f_ca_w_1_120_s_0_560=3.49e-04 mcm2m1f_cc_w_1_120_s_0_560=3.49e-11 mcm2m1f_cf_w_1_120_s_0_560=5.12e-11
+  mcm2m1f_ca_w_1_120_s_0_840=3.49e-04 mcm2m1f_cc_w_1_120_s_0_840=1.77e-11 mcm2m1f_cf_w_1_120_s_0_840=6.28e-11
+  mcm2m1f_ca_w_1_120_s_1_540=3.49e-04 mcm2m1f_cc_w_1_120_s_1_540=4.12e-12 mcm2m1f_cf_w_1_120_s_1_540=7.48e-11
+  mcm2m1f_ca_w_1_120_s_3_500=3.49e-04 mcm2m1f_cc_w_1_120_s_3_500=1.35e-13 mcm2m1f_cf_w_1_120_s_3_500=7.91e-11
+  mcm2m1d_ca_w_0_140_s_0_140=3.58e-04 mcm2m1d_cc_w_0_140_s_0_140=1.06e-10 mcm2m1d_cf_w_0_140_s_0_140=1.63e-11
+  mcm2m1d_ca_w_0_140_s_0_175=3.58e-04 mcm2m1d_cc_w_0_140_s_0_175=1.01e-10 mcm2m1d_cf_w_0_140_s_0_175=2.08e-11
+  mcm2m1d_ca_w_0_140_s_0_210=3.58e-04 mcm2m1d_cc_w_0_140_s_0_210=9.28e-11 mcm2m1d_cf_w_0_140_s_0_210=2.48e-11
+  mcm2m1d_ca_w_0_140_s_0_280=3.58e-04 mcm2m1d_cc_w_0_140_s_0_280=7.50e-11 mcm2m1d_cf_w_0_140_s_0_280=3.19e-11
+  mcm2m1d_ca_w_0_140_s_0_350=3.58e-04 mcm2m1d_cc_w_0_140_s_0_350=5.99e-11 mcm2m1d_cf_w_0_140_s_0_350=3.83e-11
+  mcm2m1d_ca_w_0_140_s_0_420=3.58e-04 mcm2m1d_cc_w_0_140_s_0_420=4.70e-11 mcm2m1d_cf_w_0_140_s_0_420=4.43e-11
+  mcm2m1d_ca_w_0_140_s_0_560=3.58e-04 mcm2m1d_cc_w_0_140_s_0_560=3.04e-11 mcm2m1d_cf_w_0_140_s_0_560=5.32e-11
+  mcm2m1d_ca_w_0_140_s_0_840=3.58e-04 mcm2m1d_cc_w_0_140_s_0_840=1.44e-11 mcm2m1d_cf_w_0_140_s_0_840=6.50e-11
+  mcm2m1d_ca_w_0_140_s_1_540=3.58e-04 mcm2m1d_cc_w_0_140_s_1_540=2.75e-12 mcm2m1d_cf_w_0_140_s_1_540=7.59e-11
+  mcm2m1d_ca_w_0_140_s_3_500=3.58e-04 mcm2m1d_cc_w_0_140_s_3_500=1.05e-13 mcm2m1d_cf_w_0_140_s_3_500=7.90e-11
+  mcm2m1d_ca_w_1_120_s_0_140=3.58e-04 mcm2m1d_cc_w_1_120_s_0_140=1.13e-10 mcm2m1d_cf_w_1_120_s_0_140=1.64e-11
+  mcm2m1d_ca_w_1_120_s_0_175=3.58e-04 mcm2m1d_cc_w_1_120_s_0_175=1.06e-10 mcm2m1d_cf_w_1_120_s_0_175=2.08e-11
+  mcm2m1d_ca_w_1_120_s_0_210=3.58e-04 mcm2m1d_cc_w_1_120_s_0_210=9.70e-11 mcm2m1d_cf_w_1_120_s_0_210=2.48e-11
+  mcm2m1d_ca_w_1_120_s_0_280=3.58e-04 mcm2m1d_cc_w_1_120_s_0_280=7.81e-11 mcm2m1d_cf_w_1_120_s_0_280=3.20e-11
+  mcm2m1d_ca_w_1_120_s_0_350=3.58e-04 mcm2m1d_cc_w_1_120_s_0_350=6.27e-11 mcm2m1d_cf_w_1_120_s_0_350=3.84e-11
+  mcm2m1d_ca_w_1_120_s_0_420=3.58e-04 mcm2m1d_cc_w_1_120_s_0_420=4.96e-11 mcm2m1d_cf_w_1_120_s_0_420=4.43e-11
+  mcm2m1d_ca_w_1_120_s_0_560=3.58e-04 mcm2m1d_cc_w_1_120_s_0_560=3.23e-11 mcm2m1d_cf_w_1_120_s_0_560=5.33e-11
+  mcm2m1d_ca_w_1_120_s_0_840=3.58e-04 mcm2m1d_cc_w_1_120_s_0_840=1.53e-11 mcm2m1d_cf_w_1_120_s_0_840=6.52e-11
+  mcm2m1d_ca_w_1_120_s_1_540=3.58e-04 mcm2m1d_cc_w_1_120_s_1_540=2.98e-12 mcm2m1d_cf_w_1_120_s_1_540=7.66e-11
+  mcm2m1d_ca_w_1_120_s_3_500=3.58e-04 mcm2m1d_cc_w_1_120_s_3_500=9.50e-14 mcm2m1d_cf_w_1_120_s_3_500=8.02e-11
+  mcm2m1p1_ca_w_0_140_s_0_140=3.86e-04 mcm2m1p1_cc_w_0_140_s_0_140=1.03e-10 mcm2m1p1_cf_w_0_140_s_0_140=1.78e-11
+  mcm2m1p1_ca_w_0_140_s_0_175=3.86e-04 mcm2m1p1_cc_w_0_140_s_0_175=9.73e-11 mcm2m1p1_cf_w_0_140_s_0_175=2.27e-11
+  mcm2m1p1_ca_w_0_140_s_0_210=3.86e-04 mcm2m1p1_cc_w_0_140_s_0_210=8.94e-11 mcm2m1p1_cf_w_0_140_s_0_210=2.72e-11
+  mcm2m1p1_ca_w_0_140_s_0_280=3.86e-04 mcm2m1p1_cc_w_0_140_s_0_280=7.10e-11 mcm2m1p1_cf_w_0_140_s_0_280=3.53e-11
+  mcm2m1p1_ca_w_0_140_s_0_350=3.86e-04 mcm2m1p1_cc_w_0_140_s_0_350=5.56e-11 mcm2m1p1_cf_w_0_140_s_0_350=4.25e-11
+  mcm2m1p1_ca_w_0_140_s_0_420=3.86e-04 mcm2m1p1_cc_w_0_140_s_0_420=4.25e-11 mcm2m1p1_cf_w_0_140_s_0_420=4.90e-11
+  mcm2m1p1_ca_w_0_140_s_0_560=3.86e-04 mcm2m1p1_cc_w_0_140_s_0_560=2.62e-11 mcm2m1p1_cf_w_0_140_s_0_560=5.90e-11
+  mcm2m1p1_ca_w_0_140_s_0_840=3.86e-04 mcm2m1p1_cc_w_0_140_s_0_840=1.06e-11 mcm2m1p1_cf_w_0_140_s_0_840=7.15e-11
+  mcm2m1p1_ca_w_0_140_s_1_540=3.86e-04 mcm2m1p1_cc_w_0_140_s_1_540=1.32e-12 mcm2m1p1_cf_w_0_140_s_1_540=8.08e-11
+  mcm2m1p1_ca_w_0_140_s_3_500=3.86e-04 mcm2m1p1_cc_w_0_140_s_3_500=3.50e-14 mcm2m1p1_cf_w_0_140_s_3_500=8.27e-11
+  mcm2m1p1_ca_w_1_120_s_0_140=3.86e-04 mcm2m1p1_cc_w_1_120_s_0_140=1.07e-10 mcm2m1p1_cf_w_1_120_s_0_140=1.79e-11
+  mcm2m1p1_ca_w_1_120_s_0_175=3.86e-04 mcm2m1p1_cc_w_1_120_s_0_175=1.00e-10 mcm2m1p1_cf_w_1_120_s_0_175=2.28e-11
+  mcm2m1p1_ca_w_1_120_s_0_210=3.86e-04 mcm2m1p1_cc_w_1_120_s_0_210=9.11e-11 mcm2m1p1_cf_w_1_120_s_0_210=2.73e-11
+  mcm2m1p1_ca_w_1_120_s_0_280=3.86e-04 mcm2m1p1_cc_w_1_120_s_0_280=7.25e-11 mcm2m1p1_cf_w_1_120_s_0_280=3.54e-11
+  mcm2m1p1_ca_w_1_120_s_0_350=3.86e-04 mcm2m1p1_cc_w_1_120_s_0_350=5.68e-11 mcm2m1p1_cf_w_1_120_s_0_350=4.26e-11
+  mcm2m1p1_ca_w_1_120_s_0_420=3.86e-04 mcm2m1p1_cc_w_1_120_s_0_420=4.38e-11 mcm2m1p1_cf_w_1_120_s_0_420=4.91e-11
+  mcm2m1p1_ca_w_1_120_s_0_560=3.86e-04 mcm2m1p1_cc_w_1_120_s_0_560=2.67e-11 mcm2m1p1_cf_w_1_120_s_0_560=5.91e-11
+  mcm2m1p1_ca_w_1_120_s_0_840=3.86e-04 mcm2m1p1_cc_w_1_120_s_0_840=1.09e-11 mcm2m1p1_cf_w_1_120_s_0_840=7.17e-11
+  mcm2m1p1_ca_w_1_120_s_1_540=3.86e-04 mcm2m1p1_cc_w_1_120_s_1_540=1.35e-12 mcm2m1p1_cf_w_1_120_s_1_540=8.12e-11
+  mcm2m1p1_ca_w_1_120_s_3_500=3.86e-04 mcm2m1p1_cc_w_1_120_s_3_500=0.00e+00 mcm2m1p1_cf_w_1_120_s_3_500=8.32e-11
+  mcm2m1l1_ca_w_0_140_s_0_140=5.28e-04 mcm2m1l1_cc_w_0_140_s_0_140=9.37e-11 mcm2m1l1_cf_w_0_140_s_0_140=2.44e-11
+  mcm2m1l1_ca_w_0_140_s_0_175=5.28e-04 mcm2m1l1_cc_w_0_140_s_0_175=8.65e-11 mcm2m1l1_cf_w_0_140_s_0_175=3.18e-11
+  mcm2m1l1_ca_w_0_140_s_0_210=5.28e-04 mcm2m1l1_cc_w_0_140_s_0_210=7.83e-11 mcm2m1l1_cf_w_0_140_s_0_210=3.85e-11
+  mcm2m1l1_ca_w_0_140_s_0_280=5.28e-04 mcm2m1l1_cc_w_0_140_s_0_280=5.99e-11 mcm2m1l1_cf_w_0_140_s_0_280=5.05e-11
+  mcm2m1l1_ca_w_0_140_s_0_350=5.28e-04 mcm2m1l1_cc_w_0_140_s_0_350=4.44e-11 mcm2m1l1_cf_w_0_140_s_0_350=6.08e-11
+  mcm2m1l1_ca_w_0_140_s_0_420=5.28e-04 mcm2m1l1_cc_w_0_140_s_0_420=3.20e-11 mcm2m1l1_cf_w_0_140_s_0_420=6.97e-11
+  mcm2m1l1_ca_w_0_140_s_0_560=5.28e-04 mcm2m1l1_cc_w_0_140_s_0_560=1.65e-11 mcm2m1l1_cf_w_0_140_s_0_560=8.23e-11
+  mcm2m1l1_ca_w_0_140_s_0_840=5.28e-04 mcm2m1l1_cc_w_0_140_s_0_840=4.55e-12 mcm2m1l1_cf_w_0_140_s_0_840=9.45e-11
+  mcm2m1l1_ca_w_0_140_s_1_540=5.28e-04 mcm2m1l1_cc_w_0_140_s_1_540=3.50e-13 mcm2m1l1_cf_w_0_140_s_1_540=1.01e-10
+  mcm2m1l1_ca_w_0_140_s_3_500=5.28e-04 mcm2m1l1_cc_w_0_140_s_3_500=0.00e+00 mcm2m1l1_cf_w_0_140_s_3_500=1.02e-10
+  mcm2m1l1_ca_w_1_120_s_0_140=5.28e-04 mcm2m1l1_cc_w_1_120_s_0_140=9.36e-11 mcm2m1l1_cf_w_1_120_s_0_140=2.45e-11
+  mcm2m1l1_ca_w_1_120_s_0_175=5.28e-04 mcm2m1l1_cc_w_1_120_s_0_175=8.75e-11 mcm2m1l1_cf_w_1_120_s_0_175=3.19e-11
+  mcm2m1l1_ca_w_1_120_s_0_210=5.28e-04 mcm2m1l1_cc_w_1_120_s_0_210=7.85e-11 mcm2m1l1_cf_w_1_120_s_0_210=3.86e-11
+  mcm2m1l1_ca_w_1_120_s_0_280=5.28e-04 mcm2m1l1_cc_w_1_120_s_0_280=5.99e-11 mcm2m1l1_cf_w_1_120_s_0_280=5.07e-11
+  mcm2m1l1_ca_w_1_120_s_0_350=5.28e-04 mcm2m1l1_cc_w_1_120_s_0_350=4.44e-11 mcm2m1l1_cf_w_1_120_s_0_350=6.11e-11
+  mcm2m1l1_ca_w_1_120_s_0_420=5.28e-04 mcm2m1l1_cc_w_1_120_s_0_420=3.20e-11 mcm2m1l1_cf_w_1_120_s_0_420=6.99e-11
+  mcm2m1l1_ca_w_1_120_s_0_560=5.28e-04 mcm2m1l1_cc_w_1_120_s_0_560=1.64e-11 mcm2m1l1_cf_w_1_120_s_0_560=8.26e-11
+  mcm2m1l1_ca_w_1_120_s_0_840=5.28e-04 mcm2m1l1_cc_w_1_120_s_0_840=4.55e-12 mcm2m1l1_cf_w_1_120_s_0_840=9.48e-11
+  mcm2m1l1_ca_w_1_120_s_1_540=5.28e-04 mcm2m1l1_cc_w_1_120_s_1_540=3.00e-13 mcm2m1l1_cf_w_1_120_s_1_540=1.01e-10
+  mcm2m1l1_ca_w_1_120_s_3_500=5.28e-04 mcm2m1l1_cc_w_1_120_s_3_500=5.00e-14 mcm2m1l1_cf_w_1_120_s_3_500=1.02e-10
+  mcm3m1f_ca_w_0_140_s_0_140=8.09e-05 mcm3m1f_cc_w_0_140_s_0_140=1.25e-10 mcm3m1f_cf_w_0_140_s_0_140=4.32e-12
+  mcm3m1f_ca_w_0_140_s_0_175=8.09e-05 mcm3m1f_cc_w_0_140_s_0_175=1.19e-10 mcm3m1f_cf_w_0_140_s_0_175=5.69e-12
+  mcm3m1f_ca_w_0_140_s_0_210=8.09e-05 mcm3m1f_cc_w_0_140_s_0_210=1.11e-10 mcm3m1f_cf_w_0_140_s_0_210=7.05e-12
+  mcm3m1f_ca_w_0_140_s_0_280=8.09e-05 mcm3m1f_cc_w_0_140_s_0_280=9.30e-11 mcm3m1f_cf_w_0_140_s_0_280=9.70e-12
+  mcm3m1f_ca_w_0_140_s_0_350=8.09e-05 mcm3m1f_cc_w_0_140_s_0_350=7.76e-11 mcm3m1f_cf_w_0_140_s_0_350=1.23e-11
+  mcm3m1f_ca_w_0_140_s_0_420=8.09e-05 mcm3m1f_cc_w_0_140_s_0_420=6.48e-11 mcm3m1f_cf_w_0_140_s_0_420=1.48e-11
+  mcm3m1f_ca_w_0_140_s_0_560=8.09e-05 mcm3m1f_cc_w_0_140_s_0_560=4.77e-11 mcm3m1f_cf_w_0_140_s_0_560=1.95e-11
+  mcm3m1f_ca_w_0_140_s_0_840=8.09e-05 mcm3m1f_cc_w_0_140_s_0_840=2.88e-11 mcm3m1f_cf_w_0_140_s_0_840=2.75e-11
+  mcm3m1f_ca_w_0_140_s_1_540=8.09e-05 mcm3m1f_cc_w_0_140_s_1_540=9.94e-12 mcm3m1f_cf_w_0_140_s_1_540=4.04e-11
+  mcm3m1f_ca_w_0_140_s_3_500=8.09e-05 mcm3m1f_cc_w_0_140_s_3_500=6.75e-13 mcm3m1f_cf_w_0_140_s_3_500=4.88e-11
+  mcm3m1f_ca_w_1_120_s_0_140=8.09e-05 mcm3m1f_cc_w_1_120_s_0_140=1.35e-10 mcm3m1f_cf_w_1_120_s_0_140=4.39e-12
+  mcm3m1f_ca_w_1_120_s_0_175=8.09e-05 mcm3m1f_cc_w_1_120_s_0_175=1.29e-10 mcm3m1f_cf_w_1_120_s_0_175=5.75e-12
+  mcm3m1f_ca_w_1_120_s_0_210=8.09e-05 mcm3m1f_cc_w_1_120_s_0_210=1.20e-10 mcm3m1f_cf_w_1_120_s_0_210=7.10e-12
+  mcm3m1f_ca_w_1_120_s_0_280=8.09e-05 mcm3m1f_cc_w_1_120_s_0_280=1.00e-10 mcm3m1f_cf_w_1_120_s_0_280=9.76e-12
+  mcm3m1f_ca_w_1_120_s_0_350=8.09e-05 mcm3m1f_cc_w_1_120_s_0_350=8.38e-11 mcm3m1f_cf_w_1_120_s_0_350=1.24e-11
+  mcm3m1f_ca_w_1_120_s_0_420=8.09e-05 mcm3m1f_cc_w_1_120_s_0_420=7.03e-11 mcm3m1f_cf_w_1_120_s_0_420=1.49e-11
+  mcm3m1f_ca_w_1_120_s_0_560=8.09e-05 mcm3m1f_cc_w_1_120_s_0_560=5.15e-11 mcm3m1f_cf_w_1_120_s_0_560=1.97e-11
+  mcm3m1f_ca_w_1_120_s_0_840=8.09e-05 mcm3m1f_cc_w_1_120_s_0_840=3.10e-11 mcm3m1f_cf_w_1_120_s_0_840=2.79e-11
+  mcm3m1f_ca_w_1_120_s_1_540=8.09e-05 mcm3m1f_cc_w_1_120_s_1_540=1.08e-11 mcm3m1f_cf_w_1_120_s_1_540=4.13e-11
+  mcm3m1f_ca_w_1_120_s_3_500=8.09e-05 mcm3m1f_cc_w_1_120_s_3_500=7.25e-13 mcm3m1f_cf_w_1_120_s_3_500=5.05e-11
+  mcm3m1d_ca_w_0_140_s_0_140=9.07e-05 mcm3m1d_cc_w_0_140_s_0_140=1.24e-10 mcm3m1d_cf_w_0_140_s_0_140=4.85e-12
+  mcm3m1d_ca_w_0_140_s_0_175=9.07e-05 mcm3m1d_cc_w_0_140_s_0_175=1.18e-10 mcm3m1d_cf_w_0_140_s_0_175=6.38e-12
+  mcm3m1d_ca_w_0_140_s_0_210=9.07e-05 mcm3m1d_cc_w_0_140_s_0_210=1.09e-10 mcm3m1d_cf_w_0_140_s_0_210=7.91e-12
+  mcm3m1d_ca_w_0_140_s_0_280=9.07e-05 mcm3m1d_cc_w_0_140_s_0_280=9.14e-11 mcm3m1d_cf_w_0_140_s_0_280=1.09e-11
+  mcm3m1d_ca_w_0_140_s_0_350=9.07e-05 mcm3m1d_cc_w_0_140_s_0_350=7.59e-11 mcm3m1d_cf_w_0_140_s_0_350=1.38e-11
+  mcm3m1d_ca_w_0_140_s_0_420=9.07e-05 mcm3m1d_cc_w_0_140_s_0_420=6.28e-11 mcm3m1d_cf_w_0_140_s_0_420=1.66e-11
+  mcm3m1d_ca_w_0_140_s_0_560=9.07e-05 mcm3m1d_cc_w_0_140_s_0_560=4.56e-11 mcm3m1d_cf_w_0_140_s_0_560=2.18e-11
+  mcm3m1d_ca_w_0_140_s_0_840=9.07e-05 mcm3m1d_cc_w_0_140_s_0_840=2.67e-11 mcm3m1d_cf_w_0_140_s_0_840=3.05e-11
+  mcm3m1d_ca_w_0_140_s_1_540=9.07e-05 mcm3m1d_cc_w_0_140_s_1_540=8.30e-12 mcm3m1d_cf_w_0_140_s_1_540=4.38e-11
+  mcm3m1d_ca_w_0_140_s_3_500=9.07e-05 mcm3m1d_cc_w_0_140_s_3_500=4.40e-13 mcm3m1d_cf_w_0_140_s_3_500=5.12e-11
+  mcm3m1d_ca_w_1_120_s_0_140=9.07e-05 mcm3m1d_cc_w_1_120_s_0_140=1.32e-10 mcm3m1d_cf_w_1_120_s_0_140=4.93e-12
+  mcm3m1d_ca_w_1_120_s_0_175=9.07e-05 mcm3m1d_cc_w_1_120_s_0_175=1.26e-10 mcm3m1d_cf_w_1_120_s_0_175=6.47e-12
+  mcm3m1d_ca_w_1_120_s_0_210=9.07e-05 mcm3m1d_cc_w_1_120_s_0_210=1.17e-10 mcm3m1d_cf_w_1_120_s_0_210=8.00e-12
+  mcm3m1d_ca_w_1_120_s_0_280=9.07e-05 mcm3m1d_cc_w_1_120_s_0_280=9.75e-11 mcm3m1d_cf_w_1_120_s_0_280=1.10e-11
+  mcm3m1d_ca_w_1_120_s_0_350=9.07e-05 mcm3m1d_cc_w_1_120_s_0_350=8.10e-11 mcm3m1d_cf_w_1_120_s_0_350=1.39e-11
+  mcm3m1d_ca_w_1_120_s_0_420=9.07e-05 mcm3m1d_cc_w_1_120_s_0_420=6.74e-11 mcm3m1d_cf_w_1_120_s_0_420=1.67e-11
+  mcm3m1d_ca_w_1_120_s_0_560=9.07e-05 mcm3m1d_cc_w_1_120_s_0_560=4.87e-11 mcm3m1d_cf_w_1_120_s_0_560=2.20e-11
+  mcm3m1d_ca_w_1_120_s_0_840=9.07e-05 mcm3m1d_cc_w_1_120_s_0_840=2.84e-11 mcm3m1d_cf_w_1_120_s_0_840=3.09e-11
+  mcm3m1d_ca_w_1_120_s_1_540=9.07e-05 mcm3m1d_cc_w_1_120_s_1_540=8.97e-12 mcm3m1d_cf_w_1_120_s_1_540=4.46e-11
+  mcm3m1d_ca_w_1_120_s_3_500=9.07e-05 mcm3m1d_cc_w_1_120_s_3_500=4.50e-13 mcm3m1d_cf_w_1_120_s_3_500=5.26e-11
+  mcm3m1p1_ca_w_0_140_s_0_140=1.18e-04 mcm3m1p1_cc_w_0_140_s_0_140=1.19e-10 mcm3m1p1_cf_w_0_140_s_0_140=6.33e-12
+  mcm3m1p1_ca_w_0_140_s_0_175=1.18e-04 mcm3m1p1_cc_w_0_140_s_0_175=1.13e-10 mcm3m1p1_cf_w_0_140_s_0_175=8.35e-12
+  mcm3m1p1_ca_w_0_140_s_0_210=1.18e-04 mcm3m1p1_cc_w_0_140_s_0_210=1.05e-10 mcm3m1p1_cf_w_0_140_s_0_210=1.03e-11
+  mcm3m1p1_ca_w_0_140_s_0_280=1.18e-04 mcm3m1p1_cc_w_0_140_s_0_280=8.72e-11 mcm3m1p1_cf_w_0_140_s_0_280=1.42e-11
+  mcm3m1p1_ca_w_0_140_s_0_350=1.18e-04 mcm3m1p1_cc_w_0_140_s_0_350=7.16e-11 mcm3m1p1_cf_w_0_140_s_0_350=1.79e-11
+  mcm3m1p1_ca_w_0_140_s_0_420=1.18e-04 mcm3m1p1_cc_w_0_140_s_0_420=5.91e-11 mcm3m1p1_cf_w_0_140_s_0_420=2.14e-11
+  mcm3m1p1_ca_w_0_140_s_0_560=1.18e-04 mcm3m1p1_cc_w_0_140_s_0_560=4.11e-11 mcm3m1p1_cf_w_0_140_s_0_560=2.79e-11
+  mcm3m1p1_ca_w_0_140_s_0_840=1.18e-04 mcm3m1p1_cc_w_0_140_s_0_840=2.21e-11 mcm3m1p1_cf_w_0_140_s_0_840=3.82e-11
+  mcm3m1p1_ca_w_0_140_s_1_540=1.18e-04 mcm3m1p1_cc_w_0_140_s_1_540=5.59e-12 mcm3m1p1_cf_w_0_140_s_1_540=5.14e-11
+  mcm3m1p1_ca_w_0_140_s_3_500=1.18e-04 mcm3m1p1_cc_w_0_140_s_3_500=2.25e-13 mcm3m1p1_cf_w_0_140_s_3_500=5.69e-11
+  mcm3m1p1_ca_w_1_120_s_0_140=1.18e-04 mcm3m1p1_cc_w_1_120_s_0_140=1.27e-10 mcm3m1p1_cf_w_1_120_s_0_140=6.52e-12
+  mcm3m1p1_ca_w_1_120_s_0_175=1.18e-04 mcm3m1p1_cc_w_1_120_s_0_175=1.21e-10 mcm3m1p1_cf_w_1_120_s_0_175=8.55e-12
+  mcm3m1p1_ca_w_1_120_s_0_210=1.18e-04 mcm3m1p1_cc_w_1_120_s_0_210=1.12e-10 mcm3m1p1_cf_w_1_120_s_0_210=1.05e-11
+  mcm3m1p1_ca_w_1_120_s_0_280=1.18e-04 mcm3m1p1_cc_w_1_120_s_0_280=9.15e-11 mcm3m1p1_cf_w_1_120_s_0_280=1.44e-11
+  mcm3m1p1_ca_w_1_120_s_0_350=1.18e-04 mcm3m1p1_cc_w_1_120_s_0_350=7.48e-11 mcm3m1p1_cf_w_1_120_s_0_350=1.81e-11
+  mcm3m1p1_ca_w_1_120_s_0_420=1.18e-04 mcm3m1p1_cc_w_1_120_s_0_420=6.16e-11 mcm3m1p1_cf_w_1_120_s_0_420=2.16e-11
+  mcm3m1p1_ca_w_1_120_s_0_560=1.18e-04 mcm3m1p1_cc_w_1_120_s_0_560=4.31e-11 mcm3m1p1_cf_w_1_120_s_0_560=2.81e-11
+  mcm3m1p1_ca_w_1_120_s_0_840=1.18e-04 mcm3m1p1_cc_w_1_120_s_0_840=2.33e-11 mcm3m1p1_cf_w_1_120_s_0_840=3.86e-11
+  mcm3m1p1_ca_w_1_120_s_1_540=1.18e-04 mcm3m1p1_cc_w_1_120_s_1_540=5.95e-12 mcm3m1p1_cf_w_1_120_s_1_540=5.23e-11
+  mcm3m1p1_ca_w_1_120_s_3_500=1.18e-04 mcm3m1p1_cc_w_1_120_s_3_500=2.15e-13 mcm3m1p1_cf_w_1_120_s_3_500=5.82e-11
+  mcm3m1l1_ca_w_0_140_s_0_140=2.60e-04 mcm3m1l1_cc_w_0_140_s_0_140=1.09e-10 mcm3m1l1_cf_w_0_140_s_0_140=1.30e-11
+  mcm3m1l1_ca_w_0_140_s_0_175=2.60e-04 mcm3m1l1_cc_w_0_140_s_0_175=1.04e-10 mcm3m1l1_cf_w_0_140_s_0_175=1.75e-11
+  mcm3m1l1_ca_w_0_140_s_0_210=2.60e-04 mcm3m1l1_cc_w_0_140_s_0_210=9.52e-11 mcm3m1l1_cf_w_0_140_s_0_210=2.17e-11
+  mcm3m1l1_ca_w_0_140_s_0_280=2.60e-04 mcm3m1l1_cc_w_0_140_s_0_280=7.63e-11 mcm3m1l1_cf_w_0_140_s_0_280=2.94e-11
+  mcm3m1l1_ca_w_0_140_s_0_350=2.60e-04 mcm3m1l1_cc_w_0_140_s_0_350=6.03e-11 mcm3m1l1_cf_w_0_140_s_0_350=3.64e-11
+  mcm3m1l1_ca_w_0_140_s_0_420=2.60e-04 mcm3m1l1_cc_w_0_140_s_0_420=4.81e-11 mcm3m1l1_cf_w_0_140_s_0_420=4.25e-11
+  mcm3m1l1_ca_w_0_140_s_0_560=2.60e-04 mcm3m1l1_cc_w_0_140_s_0_560=3.07e-11 mcm3m1l1_cf_w_0_140_s_0_560=5.24e-11
+  mcm3m1l1_ca_w_0_140_s_0_840=2.60e-04 mcm3m1l1_cc_w_0_140_s_0_840=1.41e-11 mcm3m1l1_cf_w_0_140_s_0_840=6.51e-11
+  mcm3m1l1_ca_w_0_140_s_1_540=2.60e-04 mcm3m1l1_cc_w_0_140_s_1_540=2.47e-12 mcm3m1l1_cf_w_0_140_s_1_540=7.68e-11
+  mcm3m1l1_ca_w_0_140_s_3_500=2.60e-04 mcm3m1l1_cc_w_0_140_s_3_500=3.50e-14 mcm3m1l1_cf_w_0_140_s_3_500=8.01e-11
+  mcm3m1l1_ca_w_1_120_s_0_140=2.60e-04 mcm3m1l1_cc_w_1_120_s_0_140=1.15e-10 mcm3m1l1_cf_w_1_120_s_0_140=1.32e-11
+  mcm3m1l1_ca_w_1_120_s_0_175=2.60e-04 mcm3m1l1_cc_w_1_120_s_0_175=1.08e-10 mcm3m1l1_cf_w_1_120_s_0_175=1.77e-11
+  mcm3m1l1_ca_w_1_120_s_0_210=2.60e-04 mcm3m1l1_cc_w_1_120_s_0_210=9.86e-11 mcm3m1l1_cf_w_1_120_s_0_210=2.19e-11
+  mcm3m1l1_ca_w_1_120_s_0_280=2.60e-04 mcm3m1l1_cc_w_1_120_s_0_280=7.89e-11 mcm3m1l1_cf_w_1_120_s_0_280=2.95e-11
+  mcm3m1l1_ca_w_1_120_s_0_350=2.60e-04 mcm3m1l1_cc_w_1_120_s_0_350=6.28e-11 mcm3m1l1_cf_w_1_120_s_0_350=3.66e-11
+  mcm3m1l1_ca_w_1_120_s_0_420=2.60e-04 mcm3m1l1_cc_w_1_120_s_0_420=4.98e-11 mcm3m1l1_cf_w_1_120_s_0_420=4.27e-11
+  mcm3m1l1_ca_w_1_120_s_0_560=2.60e-04 mcm3m1l1_cc_w_1_120_s_0_560=3.23e-11 mcm3m1l1_cf_w_1_120_s_0_560=5.26e-11
+  mcm3m1l1_ca_w_1_120_s_0_840=2.60e-04 mcm3m1l1_cc_w_1_120_s_0_840=1.50e-11 mcm3m1l1_cf_w_1_120_s_0_840=6.55e-11
+  mcm3m1l1_ca_w_1_120_s_1_540=2.60e-04 mcm3m1l1_cc_w_1_120_s_1_540=2.74e-12 mcm3m1l1_cf_w_1_120_s_1_540=7.76e-11
+  mcm3m1l1_ca_w_1_120_s_3_500=2.60e-04 mcm3m1l1_cc_w_1_120_s_3_500=6.00e-14 mcm3m1l1_cf_w_1_120_s_3_500=8.12e-11
+  mcm4m1f_ca_w_0_140_s_0_140=5.42e-05 mcm4m1f_cc_w_0_140_s_0_140=1.28e-10 mcm4m1f_cf_w_0_140_s_0_140=2.93e-12
+  mcm4m1f_ca_w_0_140_s_0_175=5.42e-05 mcm4m1f_cc_w_0_140_s_0_175=1.21e-10 mcm4m1f_cf_w_0_140_s_0_175=3.86e-12
+  mcm4m1f_ca_w_0_140_s_0_210=5.42e-05 mcm4m1f_cc_w_0_140_s_0_210=1.14e-10 mcm4m1f_cf_w_0_140_s_0_210=4.80e-12
+  mcm4m1f_ca_w_0_140_s_0_280=5.42e-05 mcm4m1f_cc_w_0_140_s_0_280=9.73e-11 mcm4m1f_cf_w_0_140_s_0_280=6.64e-12
+  mcm4m1f_ca_w_0_140_s_0_350=5.42e-05 mcm4m1f_cc_w_0_140_s_0_350=8.23e-11 mcm4m1f_cf_w_0_140_s_0_350=8.43e-12
+  mcm4m1f_ca_w_0_140_s_0_420=5.42e-05 mcm4m1f_cc_w_0_140_s_0_420=7.00e-11 mcm4m1f_cf_w_0_140_s_0_420=1.02e-11
+  mcm4m1f_ca_w_0_140_s_0_560=5.42e-05 mcm4m1f_cc_w_0_140_s_0_560=5.34e-11 mcm4m1f_cf_w_0_140_s_0_560=1.36e-11
+  mcm4m1f_ca_w_0_140_s_0_840=5.42e-05 mcm4m1f_cc_w_0_140_s_0_840=3.51e-11 mcm4m1f_cf_w_0_140_s_0_840=1.97e-11
+  mcm4m1f_ca_w_0_140_s_1_540=5.42e-05 mcm4m1f_cc_w_0_140_s_1_540=1.55e-11 mcm4m1f_cf_w_0_140_s_1_540=3.07e-11
+  mcm4m1f_ca_w_0_140_s_3_500=5.42e-05 mcm4m1f_cc_w_0_140_s_3_500=2.17e-12 mcm4m1f_cf_w_0_140_s_3_500=4.19e-11
+  mcm4m1f_ca_w_1_120_s_0_140=5.42e-05 mcm4m1f_cc_w_1_120_s_0_140=1.44e-10 mcm4m1f_cf_w_1_120_s_0_140=3.01e-12
+  mcm4m1f_ca_w_1_120_s_0_175=5.42e-05 mcm4m1f_cc_w_1_120_s_0_175=1.37e-10 mcm4m1f_cf_w_1_120_s_0_175=3.95e-12
+  mcm4m1f_ca_w_1_120_s_0_210=5.42e-05 mcm4m1f_cc_w_1_120_s_0_210=1.29e-10 mcm4m1f_cf_w_1_120_s_0_210=4.88e-12
+  mcm4m1f_ca_w_1_120_s_0_280=5.42e-05 mcm4m1f_cc_w_1_120_s_0_280=1.09e-10 mcm4m1f_cf_w_1_120_s_0_280=6.70e-12
+  mcm4m1f_ca_w_1_120_s_0_350=5.42e-05 mcm4m1f_cc_w_1_120_s_0_350=9.24e-11 mcm4m1f_cf_w_1_120_s_0_350=8.50e-12
+  mcm4m1f_ca_w_1_120_s_0_420=5.42e-05 mcm4m1f_cc_w_1_120_s_0_420=7.93e-11 mcm4m1f_cf_w_1_120_s_0_420=1.03e-11
+  mcm4m1f_ca_w_1_120_s_0_560=5.42e-05 mcm4m1f_cc_w_1_120_s_0_560=6.06e-11 mcm4m1f_cf_w_1_120_s_0_560=1.37e-11
+  mcm4m1f_ca_w_1_120_s_0_840=5.42e-05 mcm4m1f_cc_w_1_120_s_0_840=3.99e-11 mcm4m1f_cf_w_1_120_s_0_840=1.99e-11
+  mcm4m1f_ca_w_1_120_s_1_540=5.42e-05 mcm4m1f_cc_w_1_120_s_1_540=1.78e-11 mcm4m1f_cf_w_1_120_s_1_540=3.15e-11
+  mcm4m1f_ca_w_1_120_s_3_500=5.42e-05 mcm4m1f_cc_w_1_120_s_3_500=2.58e-12 mcm4m1f_cf_w_1_120_s_3_500=4.41e-11
+  mcm4m1d_ca_w_0_140_s_0_140=6.39e-05 mcm4m1d_cc_w_0_140_s_0_140=1.27e-10 mcm4m1d_cf_w_0_140_s_0_140=3.45e-12
+  mcm4m1d_ca_w_0_140_s_0_175=6.39e-05 mcm4m1d_cc_w_0_140_s_0_175=1.20e-10 mcm4m1d_cf_w_0_140_s_0_175=4.56e-12
+  mcm4m1d_ca_w_0_140_s_0_210=6.39e-05 mcm4m1d_cc_w_0_140_s_0_210=1.13e-10 mcm4m1d_cf_w_0_140_s_0_210=5.66e-12
+  mcm4m1d_ca_w_0_140_s_0_280=6.39e-05 mcm4m1d_cc_w_0_140_s_0_280=9.58e-11 mcm4m1d_cf_w_0_140_s_0_280=7.82e-12
+  mcm4m1d_ca_w_0_140_s_0_350=6.39e-05 mcm4m1d_cc_w_0_140_s_0_350=8.07e-11 mcm4m1d_cf_w_0_140_s_0_350=9.92e-12
+  mcm4m1d_ca_w_0_140_s_0_420=6.39e-05 mcm4m1d_cc_w_0_140_s_0_420=6.81e-11 mcm4m1d_cf_w_0_140_s_0_420=1.20e-11
+  mcm4m1d_ca_w_0_140_s_0_560=6.39e-05 mcm4m1d_cc_w_0_140_s_0_560=5.13e-11 mcm4m1d_cf_w_0_140_s_0_560=1.59e-11
+  mcm4m1d_ca_w_0_140_s_0_840=6.39e-05 mcm4m1d_cc_w_0_140_s_0_840=3.30e-11 mcm4m1d_cf_w_0_140_s_0_840=2.27e-11
+  mcm4m1d_ca_w_0_140_s_1_540=6.39e-05 mcm4m1d_cc_w_0_140_s_1_540=1.36e-11 mcm4m1d_cf_w_0_140_s_1_540=3.45e-11
+  mcm4m1d_ca_w_0_140_s_3_500=6.39e-05 mcm4m1d_cc_w_0_140_s_3_500=1.65e-12 mcm4m1d_cf_w_0_140_s_3_500=4.50e-11
+  mcm4m1d_ca_w_1_120_s_0_140=6.39e-05 mcm4m1d_cc_w_1_120_s_0_140=1.41e-10 mcm4m1d_cf_w_1_120_s_0_140=3.56e-12
+  mcm4m1d_ca_w_1_120_s_0_175=6.39e-05 mcm4m1d_cc_w_1_120_s_0_175=1.35e-10 mcm4m1d_cf_w_1_120_s_0_175=4.66e-12
+  mcm4m1d_ca_w_1_120_s_0_210=6.39e-05 mcm4m1d_cc_w_1_120_s_0_210=1.26e-10 mcm4m1d_cf_w_1_120_s_0_210=5.76e-12
+  mcm4m1d_ca_w_1_120_s_0_280=6.39e-05 mcm4m1d_cc_w_1_120_s_0_280=1.06e-10 mcm4m1d_cf_w_1_120_s_0_280=7.91e-12
+  mcm4m1d_ca_w_1_120_s_0_350=6.39e-05 mcm4m1d_cc_w_1_120_s_0_350=8.97e-11 mcm4m1d_cf_w_1_120_s_0_350=1.00e-11
+  mcm4m1d_ca_w_1_120_s_0_420=6.39e-05 mcm4m1d_cc_w_1_120_s_0_420=7.63e-11 mcm4m1d_cf_w_1_120_s_0_420=1.21e-11
+  mcm4m1d_ca_w_1_120_s_0_560=6.39e-05 mcm4m1d_cc_w_1_120_s_0_560=5.76e-11 mcm4m1d_cf_w_1_120_s_0_560=1.60e-11
+  mcm4m1d_ca_w_1_120_s_0_840=6.39e-05 mcm4m1d_cc_w_1_120_s_0_840=3.71e-11 mcm4m1d_cf_w_1_120_s_0_840=2.30e-11
+  mcm4m1d_ca_w_1_120_s_1_540=6.39e-05 mcm4m1d_cc_w_1_120_s_1_540=1.56e-11 mcm4m1d_cf_w_1_120_s_1_540=3.54e-11
+  mcm4m1d_ca_w_1_120_s_3_500=6.39e-05 mcm4m1d_cc_w_1_120_s_3_500=1.96e-12 mcm4m1d_cf_w_1_120_s_3_500=4.72e-11
+  mcm4m1p1_ca_w_0_140_s_0_140=9.17e-05 mcm4m1p1_cc_w_0_140_s_0_140=1.23e-10 mcm4m1p1_cf_w_0_140_s_0_140=4.94e-12
+  mcm4m1p1_ca_w_0_140_s_0_175=9.17e-05 mcm4m1p1_cc_w_0_140_s_0_175=1.17e-10 mcm4m1p1_cf_w_0_140_s_0_175=6.53e-12
+  mcm4m1p1_ca_w_0_140_s_0_210=9.17e-05 mcm4m1p1_cc_w_0_140_s_0_210=1.09e-10 mcm4m1p1_cf_w_0_140_s_0_210=8.11e-12
+  mcm4m1p1_ca_w_0_140_s_0_280=9.17e-05 mcm4m1p1_cc_w_0_140_s_0_280=9.16e-11 mcm4m1p1_cf_w_0_140_s_0_280=1.11e-11
+  mcm4m1p1_ca_w_0_140_s_0_350=9.17e-05 mcm4m1p1_cc_w_0_140_s_0_350=7.65e-11 mcm4m1p1_cf_w_0_140_s_0_350=1.41e-11
+  mcm4m1p1_ca_w_0_140_s_0_420=9.17e-05 mcm4m1p1_cc_w_0_140_s_0_420=6.38e-11 mcm4m1p1_cf_w_0_140_s_0_420=1.69e-11
+  mcm4m1p1_ca_w_0_140_s_0_560=9.17e-05 mcm4m1p1_cc_w_0_140_s_0_560=4.67e-11 mcm4m1p1_cf_w_0_140_s_0_560=2.20e-11
+  mcm4m1p1_ca_w_0_140_s_0_840=9.17e-05 mcm4m1p1_cc_w_0_140_s_0_840=2.84e-11 mcm4m1p1_cf_w_0_140_s_0_840=3.06e-11
+  mcm4m1p1_ca_w_0_140_s_1_540=9.17e-05 mcm4m1p1_cc_w_0_140_s_1_540=1.02e-11 mcm4m1p1_cf_w_0_140_s_1_540=4.35e-11
+  mcm4m1p1_ca_w_0_140_s_3_500=9.17e-05 mcm4m1p1_cc_w_0_140_s_3_500=9.45e-13 mcm4m1p1_cf_w_0_140_s_3_500=5.22e-11
+  mcm4m1p1_ca_w_1_120_s_0_140=9.17e-05 mcm4m1p1_cc_w_1_120_s_0_140=1.35e-10 mcm4m1p1_cf_w_1_120_s_0_140=5.22e-12
+  mcm4m1p1_ca_w_1_120_s_0_175=9.17e-05 mcm4m1p1_cc_w_1_120_s_0_175=1.29e-10 mcm4m1p1_cf_w_1_120_s_0_175=6.81e-12
+  mcm4m1p1_ca_w_1_120_s_0_210=9.17e-05 mcm4m1p1_cc_w_1_120_s_0_210=1.20e-10 mcm4m1p1_cf_w_1_120_s_0_210=8.35e-12
+  mcm4m1p1_ca_w_1_120_s_0_280=9.17e-05 mcm4m1p1_cc_w_1_120_s_0_280=1.00e-10 mcm4m1p1_cf_w_1_120_s_0_280=1.14e-11
+  mcm4m1p1_ca_w_1_120_s_0_350=9.17e-05 mcm4m1p1_cc_w_1_120_s_0_350=8.38e-11 mcm4m1p1_cf_w_1_120_s_0_350=1.43e-11
+  mcm4m1p1_ca_w_1_120_s_0_420=9.17e-05 mcm4m1p1_cc_w_1_120_s_0_420=7.04e-11 mcm4m1p1_cf_w_1_120_s_0_420=1.71e-11
+  mcm4m1p1_ca_w_1_120_s_0_560=9.17e-05 mcm4m1p1_cc_w_1_120_s_0_560=5.19e-11 mcm4m1p1_cf_w_1_120_s_0_560=2.23e-11
+  mcm4m1p1_ca_w_1_120_s_0_840=9.17e-05 mcm4m1p1_cc_w_1_120_s_0_840=3.18e-11 mcm4m1p1_cf_w_1_120_s_0_840=3.10e-11
+  mcm4m1p1_ca_w_1_120_s_1_540=9.17e-05 mcm4m1p1_cc_w_1_120_s_1_540=1.20e-11 mcm4m1p1_cf_w_1_120_s_1_540=4.46e-11
+  mcm4m1p1_ca_w_1_120_s_3_500=9.17e-05 mcm4m1p1_cc_w_1_120_s_3_500=1.16e-12 mcm4m1p1_cf_w_1_120_s_3_500=5.46e-11
+  mcm4m1l1_ca_w_0_140_s_0_140=2.34e-04 mcm4m1l1_cc_w_0_140_s_0_140=1.13e-10 mcm4m1l1_cf_w_0_140_s_0_140=1.16e-11
+  mcm4m1l1_ca_w_0_140_s_0_175=2.34e-04 mcm4m1l1_cc_w_0_140_s_0_175=1.07e-10 mcm4m1l1_cf_w_0_140_s_0_175=1.57e-11
+  mcm4m1l1_ca_w_0_140_s_0_210=2.34e-04 mcm4m1l1_cc_w_0_140_s_0_210=9.86e-11 mcm4m1l1_cf_w_0_140_s_0_210=1.95e-11
+  mcm4m1l1_ca_w_0_140_s_0_280=2.34e-04 mcm4m1l1_cc_w_0_140_s_0_280=8.04e-11 mcm4m1l1_cf_w_0_140_s_0_280=2.64e-11
+  mcm4m1l1_ca_w_0_140_s_0_350=2.34e-04 mcm4m1l1_cc_w_0_140_s_0_350=6.49e-11 mcm4m1l1_cf_w_0_140_s_0_350=3.26e-11
+  mcm4m1l1_ca_w_0_140_s_0_420=2.34e-04 mcm4m1l1_cc_w_0_140_s_0_420=5.25e-11 mcm4m1l1_cf_w_0_140_s_0_420=3.80e-11
+  mcm4m1l1_ca_w_0_140_s_0_560=2.34e-04 mcm4m1l1_cc_w_0_140_s_0_560=3.64e-11 mcm4m1l1_cf_w_0_140_s_0_560=4.68e-11
+  mcm4m1l1_ca_w_0_140_s_0_840=2.34e-04 mcm4m1l1_cc_w_0_140_s_0_840=1.97e-11 mcm4m1l1_cf_w_0_140_s_0_840=5.85e-11
+  mcm4m1l1_ca_w_0_140_s_1_540=2.34e-04 mcm4m1l1_cc_w_0_140_s_1_540=5.78e-12 mcm4m1l1_cf_w_0_140_s_1_540=7.14e-11
+  mcm4m1l1_ca_w_0_140_s_3_500=2.34e-04 mcm4m1l1_cc_w_0_140_s_3_500=4.15e-13 mcm4m1l1_cf_w_0_140_s_3_500=7.74e-11
+  mcm4m1l1_ca_w_1_120_s_0_140=2.34e-04 mcm4m1l1_cc_w_1_120_s_0_140=1.23e-10 mcm4m1l1_cf_w_1_120_s_0_140=1.19e-11
+  mcm4m1l1_ca_w_1_120_s_0_175=2.34e-04 mcm4m1l1_cc_w_1_120_s_0_175=1.17e-10 mcm4m1l1_cf_w_1_120_s_0_175=1.59e-11
+  mcm4m1l1_ca_w_1_120_s_0_210=2.34e-04 mcm4m1l1_cc_w_1_120_s_0_210=1.07e-10 mcm4m1l1_cf_w_1_120_s_0_210=1.97e-11
+  mcm4m1l1_ca_w_1_120_s_0_280=2.34e-04 mcm4m1l1_cc_w_1_120_s_0_280=8.80e-11 mcm4m1l1_cf_w_1_120_s_0_280=2.66e-11
+  mcm4m1l1_ca_w_1_120_s_0_350=2.34e-04 mcm4m1l1_cc_w_1_120_s_0_350=7.17e-11 mcm4m1l1_cf_w_1_120_s_0_350=3.28e-11
+  mcm4m1l1_ca_w_1_120_s_0_420=2.34e-04 mcm4m1l1_cc_w_1_120_s_0_420=5.88e-11 mcm4m1l1_cf_w_1_120_s_0_420=3.82e-11
+  mcm4m1l1_ca_w_1_120_s_0_560=2.34e-04 mcm4m1l1_cc_w_1_120_s_0_560=4.10e-11 mcm4m1l1_cf_w_1_120_s_0_560=4.70e-11
+  mcm4m1l1_ca_w_1_120_s_0_840=2.34e-04 mcm4m1l1_cc_w_1_120_s_0_840=2.30e-11 mcm4m1l1_cf_w_1_120_s_0_840=5.90e-11
+  mcm4m1l1_ca_w_1_120_s_1_540=2.34e-04 mcm4m1l1_cc_w_1_120_s_1_540=7.40e-12 mcm4m1l1_cf_w_1_120_s_1_540=7.27e-11
+  mcm4m1l1_ca_w_1_120_s_3_500=2.34e-04 mcm4m1l1_cc_w_1_120_s_3_500=5.60e-13 mcm4m1l1_cf_w_1_120_s_3_500=8.01e-11
+  mcm5m1f_ca_w_0_140_s_0_140=4.68e-05 mcm5m1f_cc_w_0_140_s_0_140=1.29e-10 mcm5m1f_cf_w_0_140_s_0_140=2.54e-12
+  mcm5m1f_ca_w_0_140_s_0_175=4.68e-05 mcm5m1f_cc_w_0_140_s_0_175=1.23e-10 mcm5m1f_cf_w_0_140_s_0_175=3.35e-12
+  mcm5m1f_ca_w_0_140_s_0_210=4.68e-05 mcm5m1f_cc_w_0_140_s_0_210=1.15e-10 mcm5m1f_cf_w_0_140_s_0_210=4.16e-12
+  mcm5m1f_ca_w_0_140_s_0_280=4.68e-05 mcm5m1f_cc_w_0_140_s_0_280=9.86e-11 mcm5m1f_cf_w_0_140_s_0_280=5.76e-12
+  mcm5m1f_ca_w_0_140_s_0_350=4.68e-05 mcm5m1f_cc_w_0_140_s_0_350=8.39e-11 mcm5m1f_cf_w_0_140_s_0_350=7.32e-12
+  mcm5m1f_ca_w_0_140_s_0_420=4.68e-05 mcm5m1f_cc_w_0_140_s_0_420=7.17e-11 mcm5m1f_cf_w_0_140_s_0_420=8.91e-12
+  mcm5m1f_ca_w_0_140_s_0_560=4.68e-05 mcm5m1f_cc_w_0_140_s_0_560=5.53e-11 mcm5m1f_cf_w_0_140_s_0_560=1.18e-11
+  mcm5m1f_ca_w_0_140_s_0_840=4.68e-05 mcm5m1f_cc_w_0_140_s_0_840=3.76e-11 mcm5m1f_cf_w_0_140_s_0_840=1.72e-11
+  mcm5m1f_ca_w_0_140_s_1_540=4.68e-05 mcm5m1f_cc_w_0_140_s_1_540=1.82e-11 mcm5m1f_cf_w_0_140_s_1_540=2.74e-11
+  mcm5m1f_ca_w_0_140_s_3_500=4.68e-05 mcm5m1f_cc_w_0_140_s_3_500=3.63e-12 mcm5m1f_cf_w_0_140_s_3_500=3.91e-11
+  mcm5m1f_ca_w_1_120_s_0_140=4.68e-05 mcm5m1f_cc_w_1_120_s_0_140=1.47e-10 mcm5m1f_cf_w_1_120_s_0_140=2.62e-12
+  mcm5m1f_ca_w_1_120_s_0_175=4.68e-05 mcm5m1f_cc_w_1_120_s_0_175=1.41e-10 mcm5m1f_cf_w_1_120_s_0_175=3.44e-12
+  mcm5m1f_ca_w_1_120_s_0_210=4.68e-05 mcm5m1f_cc_w_1_120_s_0_210=1.33e-10 mcm5m1f_cf_w_1_120_s_0_210=4.25e-12
+  mcm5m1f_ca_w_1_120_s_0_280=4.68e-05 mcm5m1f_cc_w_1_120_s_0_280=1.13e-10 mcm5m1f_cf_w_1_120_s_0_280=5.84e-12
+  mcm5m1f_ca_w_1_120_s_0_350=4.68e-05 mcm5m1f_cc_w_1_120_s_0_350=9.62e-11 mcm5m1f_cf_w_1_120_s_0_350=7.41e-12
+  mcm5m1f_ca_w_1_120_s_0_420=4.68e-05 mcm5m1f_cc_w_1_120_s_0_420=8.32e-11 mcm5m1f_cf_w_1_120_s_0_420=8.94e-12
+  mcm5m1f_ca_w_1_120_s_0_560=4.68e-05 mcm5m1f_cc_w_1_120_s_0_560=6.45e-11 mcm5m1f_cf_w_1_120_s_0_560=1.19e-11
+  mcm5m1f_ca_w_1_120_s_0_840=4.68e-05 mcm5m1f_cc_w_1_120_s_0_840=4.40e-11 mcm5m1f_cf_w_1_120_s_0_840=1.74e-11
+  mcm5m1f_ca_w_1_120_s_1_540=4.68e-05 mcm5m1f_cc_w_1_120_s_1_540=2.18e-11 mcm5m1f_cf_w_1_120_s_1_540=2.80e-11
+  mcm5m1f_ca_w_1_120_s_3_500=4.68e-05 mcm5m1f_cc_w_1_120_s_3_500=4.61e-12 mcm5m1f_cf_w_1_120_s_3_500=4.14e-11
+  mcm5m1d_ca_w_0_140_s_0_140=5.66e-05 mcm5m1d_cc_w_0_140_s_0_140=1.28e-10 mcm5m1d_cf_w_0_140_s_0_140=3.06e-12
+  mcm5m1d_ca_w_0_140_s_0_175=5.66e-05 mcm5m1d_cc_w_0_140_s_0_175=1.22e-10 mcm5m1d_cf_w_0_140_s_0_175=4.04e-12
+  mcm5m1d_ca_w_0_140_s_0_210=5.66e-05 mcm5m1d_cc_w_0_140_s_0_210=1.14e-10 mcm5m1d_cf_w_0_140_s_0_210=5.03e-12
+  mcm5m1d_ca_w_0_140_s_0_280=5.66e-05 mcm5m1d_cc_w_0_140_s_0_280=9.68e-11 mcm5m1d_cf_w_0_140_s_0_280=6.94e-12
+  mcm5m1d_ca_w_0_140_s_0_350=5.66e-05 mcm5m1d_cc_w_0_140_s_0_350=8.22e-11 mcm5m1d_cf_w_0_140_s_0_350=8.81e-12
+  mcm5m1d_ca_w_0_140_s_0_420=5.66e-05 mcm5m1d_cc_w_0_140_s_0_420=6.99e-11 mcm5m1d_cf_w_0_140_s_0_420=1.07e-11
+  mcm5m1d_ca_w_0_140_s_0_560=5.66e-05 mcm5m1d_cc_w_0_140_s_0_560=5.32e-11 mcm5m1d_cf_w_0_140_s_0_560=1.41e-11
+  mcm5m1d_ca_w_0_140_s_0_840=5.66e-05 mcm5m1d_cc_w_0_140_s_0_840=3.53e-11 mcm5m1d_cf_w_0_140_s_0_840=2.03e-11
+  mcm5m1d_ca_w_0_140_s_1_540=5.66e-05 mcm5m1d_cc_w_0_140_s_1_540=1.62e-11 mcm5m1d_cf_w_0_140_s_1_540=3.14e-11
+  mcm5m1d_ca_w_0_140_s_3_500=5.66e-05 mcm5m1d_cc_w_0_140_s_3_500=2.85e-12 mcm5m1d_cf_w_0_140_s_3_500=4.26e-11
+  mcm5m1d_ca_w_1_120_s_0_140=5.66e-05 mcm5m1d_cc_w_1_120_s_0_140=1.44e-10 mcm5m1d_cf_w_1_120_s_0_140=3.19e-12
+  mcm5m1d_ca_w_1_120_s_0_175=5.66e-05 mcm5m1d_cc_w_1_120_s_0_175=1.38e-10 mcm5m1d_cf_w_1_120_s_0_175=4.16e-12
+  mcm5m1d_ca_w_1_120_s_0_210=5.66e-05 mcm5m1d_cc_w_1_120_s_0_210=1.30e-10 mcm5m1d_cf_w_1_120_s_0_210=5.13e-12
+  mcm5m1d_ca_w_1_120_s_0_280=5.66e-05 mcm5m1d_cc_w_1_120_s_0_280=1.10e-10 mcm5m1d_cf_w_1_120_s_0_280=7.05e-12
+  mcm5m1d_ca_w_1_120_s_0_350=5.66e-05 mcm5m1d_cc_w_1_120_s_0_350=9.34e-11 mcm5m1d_cf_w_1_120_s_0_350=8.93e-12
+  mcm5m1d_ca_w_1_120_s_0_420=5.66e-05 mcm5m1d_cc_w_1_120_s_0_420=8.04e-11 mcm5m1d_cf_w_1_120_s_0_420=1.08e-11
+  mcm5m1d_ca_w_1_120_s_0_560=5.66e-05 mcm5m1d_cc_w_1_120_s_0_560=6.16e-11 mcm5m1d_cf_w_1_120_s_0_560=1.43e-11
+  mcm5m1d_ca_w_1_120_s_0_840=5.66e-05 mcm5m1d_cc_w_1_120_s_0_840=4.12e-11 mcm5m1d_cf_w_1_120_s_0_840=2.06e-11
+  mcm5m1d_ca_w_1_120_s_1_540=5.66e-05 mcm5m1d_cc_w_1_120_s_1_540=1.94e-11 mcm5m1d_cf_w_1_120_s_1_540=3.21e-11
+  mcm5m1d_ca_w_1_120_s_3_500=5.66e-05 mcm5m1d_cc_w_1_120_s_3_500=3.76e-12 mcm5m1d_cf_w_1_120_s_3_500=4.51e-11
+  mcm5m1p1_ca_w_0_140_s_0_140=8.43e-05 mcm5m1p1_cc_w_0_140_s_0_140=1.23e-10 mcm5m1p1_cf_w_0_140_s_0_140=4.55e-12
+  mcm5m1p1_ca_w_0_140_s_0_175=8.43e-05 mcm5m1p1_cc_w_0_140_s_0_175=1.19e-10 mcm5m1p1_cf_w_0_140_s_0_175=6.02e-12
+  mcm5m1p1_ca_w_0_140_s_0_210=8.43e-05 mcm5m1p1_cc_w_0_140_s_0_210=1.10e-10 mcm5m1p1_cf_w_0_140_s_0_210=7.47e-12
+  mcm5m1p1_ca_w_0_140_s_0_280=8.43e-05 mcm5m1p1_cc_w_0_140_s_0_280=9.29e-11 mcm5m1p1_cf_w_0_140_s_0_280=1.03e-11
+  mcm5m1p1_ca_w_0_140_s_0_350=8.43e-05 mcm5m1p1_cc_w_0_140_s_0_350=7.79e-11 mcm5m1p1_cf_w_0_140_s_0_350=1.30e-11
+  mcm5m1p1_ca_w_0_140_s_0_420=8.43e-05 mcm5m1p1_cc_w_0_140_s_0_420=6.55e-11 mcm5m1p1_cf_w_0_140_s_0_420=1.56e-11
+  mcm5m1p1_ca_w_0_140_s_0_560=8.43e-05 mcm5m1p1_cc_w_0_140_s_0_560=4.85e-11 mcm5m1p1_cf_w_0_140_s_0_560=2.03e-11
+  mcm5m1p1_ca_w_0_140_s_0_840=8.43e-05 mcm5m1p1_cc_w_0_140_s_0_840=3.07e-11 mcm5m1p1_cf_w_0_140_s_0_840=2.83e-11
+  mcm5m1p1_ca_w_0_140_s_1_540=8.43e-05 mcm5m1p1_cc_w_0_140_s_1_540=1.25e-11 mcm5m1p1_cf_w_0_140_s_1_540=4.07e-11
+  mcm5m1p1_ca_w_0_140_s_3_500=8.43e-05 mcm5m1p1_cc_w_0_140_s_3_500=1.84e-12 mcm5m1p1_cf_w_0_140_s_3_500=5.04e-11
+  mcm5m1p1_ca_w_1_120_s_0_140=8.43e-05 mcm5m1p1_cc_w_1_120_s_0_140=1.39e-10 mcm5m1p1_cf_w_1_120_s_0_140=4.85e-12
+  mcm5m1p1_ca_w_1_120_s_0_175=8.43e-05 mcm5m1p1_cc_w_1_120_s_0_175=1.33e-10 mcm5m1p1_cf_w_1_120_s_0_175=6.32e-12
+  mcm5m1p1_ca_w_1_120_s_0_210=8.43e-05 mcm5m1p1_cc_w_1_120_s_0_210=1.24e-10 mcm5m1p1_cf_w_1_120_s_0_210=7.76e-12
+  mcm5m1p1_ca_w_1_120_s_0_280=8.43e-05 mcm5m1p1_cc_w_1_120_s_0_280=1.04e-10 mcm5m1p1_cf_w_1_120_s_0_280=1.05e-11
+  mcm5m1p1_ca_w_1_120_s_0_350=8.43e-05 mcm5m1p1_cc_w_1_120_s_0_350=8.75e-11 mcm5m1p1_cf_w_1_120_s_0_350=1.32e-11
+  mcm5m1p1_ca_w_1_120_s_0_420=8.43e-05 mcm5m1p1_cc_w_1_120_s_0_420=7.44e-11 mcm5m1p1_cf_w_1_120_s_0_420=1.58e-11
+  mcm5m1p1_ca_w_1_120_s_0_560=8.43e-05 mcm5m1p1_cc_w_1_120_s_0_560=5.58e-11 mcm5m1p1_cf_w_1_120_s_0_560=2.06e-11
+  mcm5m1p1_ca_w_1_120_s_0_840=8.43e-05 mcm5m1p1_cc_w_1_120_s_0_840=3.58e-11 mcm5m1p1_cf_w_1_120_s_0_840=2.87e-11
+  mcm5m1p1_ca_w_1_120_s_1_540=8.43e-05 mcm5m1p1_cc_w_1_120_s_1_540=1.55e-11 mcm5m1p1_cf_w_1_120_s_1_540=4.18e-11
+  mcm5m1p1_ca_w_1_120_s_3_500=8.43e-05 mcm5m1p1_cc_w_1_120_s_3_500=2.57e-12 mcm5m1p1_cf_w_1_120_s_3_500=5.33e-11
+  mcm5m1l1_ca_w_0_140_s_0_140=2.26e-04 mcm5m1l1_cc_w_0_140_s_0_140=1.13e-10 mcm5m1l1_cf_w_0_140_s_0_140=1.12e-11
+  mcm5m1l1_ca_w_0_140_s_0_175=2.26e-04 mcm5m1l1_cc_w_0_140_s_0_175=1.08e-10 mcm5m1l1_cf_w_0_140_s_0_175=1.52e-11
+  mcm5m1l1_ca_w_0_140_s_0_210=2.26e-04 mcm5m1l1_cc_w_0_140_s_0_210=9.95e-11 mcm5m1l1_cf_w_0_140_s_0_210=1.88e-11
+  mcm5m1l1_ca_w_0_140_s_0_280=2.26e-04 mcm5m1l1_cc_w_0_140_s_0_280=8.17e-11 mcm5m1l1_cf_w_0_140_s_0_280=2.55e-11
+  mcm5m1l1_ca_w_0_140_s_0_350=2.26e-04 mcm5m1l1_cc_w_0_140_s_0_350=6.65e-11 mcm5m1l1_cf_w_0_140_s_0_350=3.15e-11
+  mcm5m1l1_ca_w_0_140_s_0_420=2.26e-04 mcm5m1l1_cc_w_0_140_s_0_420=5.42e-11 mcm5m1l1_cf_w_0_140_s_0_420=3.67e-11
+  mcm5m1l1_ca_w_0_140_s_0_560=2.26e-04 mcm5m1l1_cc_w_0_140_s_0_560=3.83e-11 mcm5m1l1_cf_w_0_140_s_0_560=4.52e-11
+  mcm5m1l1_ca_w_0_140_s_0_840=2.26e-04 mcm5m1l1_cc_w_0_140_s_0_840=2.18e-11 mcm5m1l1_cf_w_0_140_s_0_840=5.65e-11
+  mcm5m1l1_ca_w_0_140_s_1_540=2.26e-04 mcm5m1l1_cc_w_0_140_s_1_540=7.45e-12 mcm5m1l1_cf_w_0_140_s_1_540=6.93e-11
+  mcm5m1l1_ca_w_0_140_s_3_500=2.26e-04 mcm5m1l1_cc_w_0_140_s_3_500=9.65e-13 mcm5m1l1_cf_w_0_140_s_3_500=7.65e-11
+  mcm5m1l1_ca_w_1_120_s_0_140=2.26e-04 mcm5m1l1_cc_w_1_120_s_0_140=1.26e-10 mcm5m1l1_cf_w_1_120_s_0_140=1.15e-11
+  mcm5m1l1_ca_w_1_120_s_0_175=2.26e-04 mcm5m1l1_cc_w_1_120_s_0_175=1.20e-10 mcm5m1l1_cf_w_1_120_s_0_175=1.55e-11
+  mcm5m1l1_ca_w_1_120_s_0_210=2.26e-04 mcm5m1l1_cc_w_1_120_s_0_210=1.11e-10 mcm5m1l1_cf_w_1_120_s_0_210=1.91e-11
+  mcm5m1l1_ca_w_1_120_s_0_280=2.26e-04 mcm5m1l1_cc_w_1_120_s_0_280=9.14e-11 mcm5m1l1_cf_w_1_120_s_0_280=2.58e-11
+  mcm5m1l1_ca_w_1_120_s_0_350=2.26e-04 mcm5m1l1_cc_w_1_120_s_0_350=7.51e-11 mcm5m1l1_cf_w_1_120_s_0_350=3.17e-11
+  mcm5m1l1_ca_w_1_120_s_0_420=2.26e-04 mcm5m1l1_cc_w_1_120_s_0_420=6.25e-11 mcm5m1l1_cf_w_1_120_s_0_420=3.69e-11
+  mcm5m1l1_ca_w_1_120_s_0_560=2.26e-04 mcm5m1l1_cc_w_1_120_s_0_560=4.48e-11 mcm5m1l1_cf_w_1_120_s_0_560=4.54e-11
+  mcm5m1l1_ca_w_1_120_s_0_840=2.26e-04 mcm5m1l1_cc_w_1_120_s_0_840=2.68e-11 mcm5m1l1_cf_w_1_120_s_0_840=5.70e-11
+  mcm5m1l1_ca_w_1_120_s_1_540=2.26e-04 mcm5m1l1_cc_w_1_120_s_1_540=1.04e-11 mcm5m1l1_cf_w_1_120_s_1_540=7.09e-11
+  mcm5m1l1_ca_w_1_120_s_3_500=2.26e-04 mcm5m1l1_cc_w_1_120_s_3_500=1.49e-12 mcm5m1l1_cf_w_1_120_s_3_500=8.01e-11
+  mcrdlm1f_ca_w_0_140_s_0_140=3.97e-05 mcrdlm1f_cc_w_0_140_s_0_140=1.31e-10 mcrdlm1f_cf_w_0_140_s_0_140=2.15e-12
+  mcrdlm1f_ca_w_0_140_s_0_175=3.97e-05 mcrdlm1f_cc_w_0_140_s_0_175=1.24e-10 mcrdlm1f_cf_w_0_140_s_0_175=2.84e-12
+  mcrdlm1f_ca_w_0_140_s_0_210=3.97e-05 mcrdlm1f_cc_w_0_140_s_0_210=1.16e-10 mcrdlm1f_cf_w_0_140_s_0_210=3.53e-12
+  mcrdlm1f_ca_w_0_140_s_0_280=3.97e-05 mcrdlm1f_cc_w_0_140_s_0_280=9.93e-11 mcrdlm1f_cf_w_0_140_s_0_280=4.89e-12
+  mcrdlm1f_ca_w_0_140_s_0_350=3.97e-05 mcrdlm1f_cc_w_0_140_s_0_350=8.49e-11 mcrdlm1f_cf_w_0_140_s_0_350=6.21e-12
+  mcrdlm1f_ca_w_0_140_s_0_420=3.97e-05 mcrdlm1f_cc_w_0_140_s_0_420=7.33e-11 mcrdlm1f_cf_w_0_140_s_0_420=7.54e-12
+  mcrdlm1f_ca_w_0_140_s_0_560=3.97e-05 mcrdlm1f_cc_w_0_140_s_0_560=5.75e-11 mcrdlm1f_cf_w_0_140_s_0_560=1.00e-11
+  mcrdlm1f_ca_w_0_140_s_0_840=3.97e-05 mcrdlm1f_cc_w_0_140_s_0_840=4.01e-11 mcrdlm1f_cf_w_0_140_s_0_840=1.46e-11
+  mcrdlm1f_ca_w_0_140_s_1_540=3.97e-05 mcrdlm1f_cc_w_0_140_s_1_540=2.17e-11 mcrdlm1f_cf_w_0_140_s_1_540=2.36e-11
+  mcrdlm1f_ca_w_0_140_s_3_500=3.97e-05 mcrdlm1f_cc_w_0_140_s_3_500=6.40e-12 mcrdlm1f_cf_w_0_140_s_3_500=3.55e-11
+  mcrdlm1f_ca_w_1_120_s_0_140=3.97e-05 mcrdlm1f_cc_w_1_120_s_0_140=1.51e-10 mcrdlm1f_cf_w_1_120_s_0_140=2.24e-12
+  mcrdlm1f_ca_w_1_120_s_0_175=3.97e-05 mcrdlm1f_cc_w_1_120_s_0_175=1.44e-10 mcrdlm1f_cf_w_1_120_s_0_175=2.93e-12
+  mcrdlm1f_ca_w_1_120_s_0_210=3.97e-05 mcrdlm1f_cc_w_1_120_s_0_210=1.36e-10 mcrdlm1f_cf_w_1_120_s_0_210=3.62e-12
+  mcrdlm1f_ca_w_1_120_s_0_280=3.97e-05 mcrdlm1f_cc_w_1_120_s_0_280=1.17e-10 mcrdlm1f_cf_w_1_120_s_0_280=4.96e-12
+  mcrdlm1f_ca_w_1_120_s_0_350=3.97e-05 mcrdlm1f_cc_w_1_120_s_0_350=1.00e-10 mcrdlm1f_cf_w_1_120_s_0_350=6.29e-12
+  mcrdlm1f_ca_w_1_120_s_0_420=3.97e-05 mcrdlm1f_cc_w_1_120_s_0_420=8.74e-11 mcrdlm1f_cf_w_1_120_s_0_420=7.60e-12
+  mcrdlm1f_ca_w_1_120_s_0_560=3.97e-05 mcrdlm1f_cc_w_1_120_s_0_560=6.89e-11 mcrdlm1f_cf_w_1_120_s_0_560=1.01e-11
+  mcrdlm1f_ca_w_1_120_s_0_840=3.97e-05 mcrdlm1f_cc_w_1_120_s_0_840=4.91e-11 mcrdlm1f_cf_w_1_120_s_0_840=1.48e-11
+  mcrdlm1f_ca_w_1_120_s_1_540=3.97e-05 mcrdlm1f_cc_w_1_120_s_1_540=2.75e-11 mcrdlm1f_cf_w_1_120_s_1_540=2.42e-11
+  mcrdlm1f_ca_w_1_120_s_3_500=3.97e-05 mcrdlm1f_cc_w_1_120_s_3_500=9.07e-12 mcrdlm1f_cf_w_1_120_s_3_500=3.77e-11
+  mcrdlm1d_ca_w_0_140_s_0_140=4.95e-05 mcrdlm1d_cc_w_0_140_s_0_140=1.29e-10 mcrdlm1d_cf_w_0_140_s_0_140=2.67e-12
+  mcrdlm1d_ca_w_0_140_s_0_175=4.95e-05 mcrdlm1d_cc_w_0_140_s_0_175=1.22e-10 mcrdlm1d_cf_w_0_140_s_0_175=3.53e-12
+  mcrdlm1d_ca_w_0_140_s_0_210=4.95e-05 mcrdlm1d_cc_w_0_140_s_0_210=1.15e-10 mcrdlm1d_cf_w_0_140_s_0_210=4.39e-12
+  mcrdlm1d_ca_w_0_140_s_0_280=4.95e-05 mcrdlm1d_cc_w_0_140_s_0_280=9.78e-11 mcrdlm1d_cf_w_0_140_s_0_280=6.06e-12
+  mcrdlm1d_ca_w_0_140_s_0_350=4.95e-05 mcrdlm1d_cc_w_0_140_s_0_350=8.32e-11 mcrdlm1d_cf_w_0_140_s_0_350=7.69e-12
+  mcrdlm1d_ca_w_0_140_s_0_420=4.95e-05 mcrdlm1d_cc_w_0_140_s_0_420=7.13e-11 mcrdlm1d_cf_w_0_140_s_0_420=9.32e-12
+  mcrdlm1d_ca_w_0_140_s_0_560=4.95e-05 mcrdlm1d_cc_w_0_140_s_0_560=5.54e-11 mcrdlm1d_cf_w_0_140_s_0_560=1.23e-11
+  mcrdlm1d_ca_w_0_140_s_0_840=4.95e-05 mcrdlm1d_cc_w_0_140_s_0_840=3.79e-11 mcrdlm1d_cf_w_0_140_s_0_840=1.77e-11
+  mcrdlm1d_ca_w_0_140_s_1_540=4.95e-05 mcrdlm1d_cc_w_0_140_s_1_540=1.95e-11 mcrdlm1d_cf_w_0_140_s_1_540=2.78e-11
+  mcrdlm1d_ca_w_0_140_s_3_500=4.95e-05 mcrdlm1d_cc_w_0_140_s_3_500=5.28e-12 mcrdlm1d_cf_w_0_140_s_3_500=3.96e-11
+  mcrdlm1d_ca_w_1_120_s_0_140=4.95e-05 mcrdlm1d_cc_w_1_120_s_0_140=1.48e-10 mcrdlm1d_cf_w_1_120_s_0_140=2.78e-12
+  mcrdlm1d_ca_w_1_120_s_0_175=4.95e-05 mcrdlm1d_cc_w_1_120_s_0_175=1.42e-10 mcrdlm1d_cf_w_1_120_s_0_175=3.65e-12
+  mcrdlm1d_ca_w_1_120_s_0_210=4.95e-05 mcrdlm1d_cc_w_1_120_s_0_210=1.34e-10 mcrdlm1d_cf_w_1_120_s_0_210=4.50e-12
+  mcrdlm1d_ca_w_1_120_s_0_280=4.95e-05 mcrdlm1d_cc_w_1_120_s_0_280=1.14e-10 mcrdlm1d_cf_w_1_120_s_0_280=6.17e-12
+  mcrdlm1d_ca_w_1_120_s_0_350=4.95e-05 mcrdlm1d_cc_w_1_120_s_0_350=9.72e-11 mcrdlm1d_cf_w_1_120_s_0_350=7.81e-12
+  mcrdlm1d_ca_w_1_120_s_0_420=4.95e-05 mcrdlm1d_cc_w_1_120_s_0_420=8.44e-11 mcrdlm1d_cf_w_1_120_s_0_420=9.41e-12
+  mcrdlm1d_ca_w_1_120_s_0_560=4.95e-05 mcrdlm1d_cc_w_1_120_s_0_560=6.60e-11 mcrdlm1d_cf_w_1_120_s_0_560=1.24e-11
+  mcrdlm1d_ca_w_1_120_s_0_840=4.95e-05 mcrdlm1d_cc_w_1_120_s_0_840=4.63e-11 mcrdlm1d_cf_w_1_120_s_0_840=1.80e-11
+  mcrdlm1d_ca_w_1_120_s_1_540=4.95e-05 mcrdlm1d_cc_w_1_120_s_1_540=2.51e-11 mcrdlm1d_cf_w_1_120_s_1_540=2.85e-11
+  mcrdlm1d_ca_w_1_120_s_3_500=4.95e-05 mcrdlm1d_cc_w_1_120_s_3_500=7.77e-12 mcrdlm1d_cf_w_1_120_s_3_500=4.21e-11
+  mcrdlm1p1_ca_w_0_140_s_0_140=7.72e-05 mcrdlm1p1_cc_w_0_140_s_0_140=1.24e-10 mcrdlm1p1_cf_w_0_140_s_0_140=4.15e-12
+  mcrdlm1p1_ca_w_0_140_s_0_175=7.72e-05 mcrdlm1p1_cc_w_0_140_s_0_175=1.19e-10 mcrdlm1p1_cf_w_0_140_s_0_175=5.50e-12
+  mcrdlm1p1_ca_w_0_140_s_0_210=7.72e-05 mcrdlm1p1_cc_w_0_140_s_0_210=1.11e-10 mcrdlm1p1_cf_w_0_140_s_0_210=6.83e-12
+  mcrdlm1p1_ca_w_0_140_s_0_280=7.72e-05 mcrdlm1p1_cc_w_0_140_s_0_280=9.40e-11 mcrdlm1p1_cf_w_0_140_s_0_280=9.40e-12
+  mcrdlm1p1_ca_w_0_140_s_0_350=7.72e-05 mcrdlm1p1_cc_w_0_140_s_0_350=7.86e-11 mcrdlm1p1_cf_w_0_140_s_0_350=1.18e-11
+  mcrdlm1p1_ca_w_0_140_s_0_420=7.72e-05 mcrdlm1p1_cc_w_0_140_s_0_420=6.68e-11 mcrdlm1p1_cf_w_0_140_s_0_420=1.43e-11
+  mcrdlm1p1_ca_w_0_140_s_0_560=7.72e-05 mcrdlm1p1_cc_w_0_140_s_0_560=5.05e-11 mcrdlm1p1_cf_w_0_140_s_0_560=1.85e-11
+  mcrdlm1p1_ca_w_0_140_s_0_840=7.72e-05 mcrdlm1p1_cc_w_0_140_s_0_840=3.31e-11 mcrdlm1p1_cf_w_0_140_s_0_840=2.59e-11
+  mcrdlm1p1_ca_w_0_140_s_1_540=7.72e-05 mcrdlm1p1_cc_w_0_140_s_1_540=1.54e-11 mcrdlm1p1_cf_w_0_140_s_1_540=3.76e-11
+  mcrdlm1p1_ca_w_0_140_s_3_500=7.72e-05 mcrdlm1p1_cc_w_0_140_s_3_500=3.65e-12 mcrdlm1p1_cf_w_0_140_s_3_500=4.83e-11
+  mcrdlm1p1_ca_w_1_120_s_0_140=7.72e-05 mcrdlm1p1_cc_w_1_120_s_0_140=1.42e-10 mcrdlm1p1_cf_w_1_120_s_0_140=4.45e-12
+  mcrdlm1p1_ca_w_1_120_s_0_175=7.72e-05 mcrdlm1p1_cc_w_1_120_s_0_175=1.35e-10 mcrdlm1p1_cf_w_1_120_s_0_175=5.76e-12
+  mcrdlm1p1_ca_w_1_120_s_0_210=7.72e-05 mcrdlm1p1_cc_w_1_120_s_0_210=1.28e-10 mcrdlm1p1_cf_w_1_120_s_0_210=7.10e-12
+  mcrdlm1p1_ca_w_1_120_s_0_280=7.72e-05 mcrdlm1p1_cc_w_1_120_s_0_280=1.08e-10 mcrdlm1p1_cf_w_1_120_s_0_280=9.64e-12
+  mcrdlm1p1_ca_w_1_120_s_0_350=7.72e-05 mcrdlm1p1_cc_w_1_120_s_0_350=9.14e-11 mcrdlm1p1_cf_w_1_120_s_0_350=1.21e-11
+  mcrdlm1p1_ca_w_1_120_s_0_420=7.72e-05 mcrdlm1p1_cc_w_1_120_s_0_420=7.83e-11 mcrdlm1p1_cf_w_1_120_s_0_420=1.45e-11
+  mcrdlm1p1_ca_w_1_120_s_0_560=7.72e-05 mcrdlm1p1_cc_w_1_120_s_0_560=6.04e-11 mcrdlm1p1_cf_w_1_120_s_0_560=1.87e-11
+  mcrdlm1p1_ca_w_1_120_s_0_840=7.72e-05 mcrdlm1p1_cc_w_1_120_s_0_840=4.09e-11 mcrdlm1p1_cf_w_1_120_s_0_840=2.61e-11
+  mcrdlm1p1_ca_w_1_120_s_1_540=7.72e-05 mcrdlm1p1_cc_w_1_120_s_1_540=2.08e-11 mcrdlm1p1_cf_w_1_120_s_1_540=3.85e-11
+  mcrdlm1p1_ca_w_1_120_s_3_500=7.72e-05 mcrdlm1p1_cc_w_1_120_s_3_500=5.92e-12 mcrdlm1p1_cf_w_1_120_s_3_500=5.14e-11
+  mcrdlm1l1_ca_w_0_140_s_0_140=2.19e-04 mcrdlm1l1_cc_w_0_140_s_0_140=1.14e-10 mcrdlm1l1_cf_w_0_140_s_0_140=1.08e-11
+  mcrdlm1l1_ca_w_0_140_s_0_175=2.19e-04 mcrdlm1l1_cc_w_0_140_s_0_175=1.09e-10 mcrdlm1l1_cf_w_0_140_s_0_175=1.46e-11
+  mcrdlm1l1_ca_w_0_140_s_0_210=2.19e-04 mcrdlm1l1_cc_w_0_140_s_0_210=1.01e-10 mcrdlm1l1_cf_w_0_140_s_0_210=1.82e-11
+  mcrdlm1l1_ca_w_0_140_s_0_280=2.19e-04 mcrdlm1l1_cc_w_0_140_s_0_280=8.30e-11 mcrdlm1l1_cf_w_0_140_s_0_280=2.47e-11
+  mcrdlm1l1_ca_w_0_140_s_0_350=2.19e-04 mcrdlm1l1_cc_w_0_140_s_0_350=6.77e-11 mcrdlm1l1_cf_w_0_140_s_0_350=3.03e-11
+  mcrdlm1l1_ca_w_0_140_s_0_420=2.19e-04 mcrdlm1l1_cc_w_0_140_s_0_420=5.58e-11 mcrdlm1l1_cf_w_0_140_s_0_420=3.54e-11
+  mcrdlm1l1_ca_w_0_140_s_0_560=2.19e-04 mcrdlm1l1_cc_w_0_140_s_0_560=3.99e-11 mcrdlm1l1_cf_w_0_140_s_0_560=4.34e-11
+  mcrdlm1l1_ca_w_0_140_s_0_840=2.19e-04 mcrdlm1l1_cc_w_0_140_s_0_840=2.41e-11 mcrdlm1l1_cf_w_0_140_s_0_840=5.43e-11
+  mcrdlm1l1_ca_w_0_140_s_1_540=2.19e-04 mcrdlm1l1_cc_w_0_140_s_1_540=9.72e-12 mcrdlm1l1_cf_w_0_140_s_1_540=6.73e-11
+  mcrdlm1l1_ca_w_0_140_s_3_500=2.19e-04 mcrdlm1l1_cc_w_0_140_s_3_500=2.05e-12 mcrdlm1l1_cf_w_0_140_s_3_500=7.53e-11
+  mcrdlm1l1_ca_w_1_120_s_0_140=2.19e-04 mcrdlm1l1_cc_w_1_120_s_0_140=1.30e-10 mcrdlm1l1_cf_w_1_120_s_0_140=1.11e-11
+  mcrdlm1l1_ca_w_1_120_s_0_175=2.19e-04 mcrdlm1l1_cc_w_1_120_s_0_175=1.23e-10 mcrdlm1l1_cf_w_1_120_s_0_175=1.49e-11
+  mcrdlm1l1_ca_w_1_120_s_0_210=2.19e-04 mcrdlm1l1_cc_w_1_120_s_0_210=1.14e-10 mcrdlm1l1_cf_w_1_120_s_0_210=1.85e-11
+  mcrdlm1l1_ca_w_1_120_s_0_280=2.19e-04 mcrdlm1l1_cc_w_1_120_s_0_280=9.50e-11 mcrdlm1l1_cf_w_1_120_s_0_280=2.49e-11
+  mcrdlm1l1_ca_w_1_120_s_0_350=2.19e-04 mcrdlm1l1_cc_w_1_120_s_0_350=7.92e-11 mcrdlm1l1_cf_w_1_120_s_0_350=3.07e-11
+  mcrdlm1l1_ca_w_1_120_s_0_420=2.19e-04 mcrdlm1l1_cc_w_1_120_s_0_420=6.66e-11 mcrdlm1l1_cf_w_1_120_s_0_420=3.56e-11
+  mcrdlm1l1_ca_w_1_120_s_0_560=2.19e-04 mcrdlm1l1_cc_w_1_120_s_0_560=4.94e-11 mcrdlm1l1_cf_w_1_120_s_0_560=4.36e-11
+  mcrdlm1l1_ca_w_1_120_s_0_840=2.19e-04 mcrdlm1l1_cc_w_1_120_s_0_840=3.17e-11 mcrdlm1l1_cf_w_1_120_s_0_840=5.47e-11
+  mcrdlm1l1_ca_w_1_120_s_1_540=2.19e-04 mcrdlm1l1_cc_w_1_120_s_1_540=1.50e-11 mcrdlm1l1_cf_w_1_120_s_1_540=6.88e-11
+  mcrdlm1l1_ca_w_1_120_s_3_500=2.19e-04 mcrdlm1l1_cc_w_1_120_s_3_500=3.93e-12 mcrdlm1l1_cf_w_1_120_s_3_500=7.98e-11
+  mcm3m2f_ca_w_0_140_s_0_140=1.55e-04 mcm3m2f_cc_w_0_140_s_0_140=1.18e-10 mcm3m2f_cf_w_0_140_s_0_140=7.85e-12
+  mcm3m2f_ca_w_0_140_s_0_175=1.55e-04 mcm3m2f_cc_w_0_140_s_0_175=1.11e-10 mcm3m2f_cf_w_0_140_s_0_175=1.02e-11
+  mcm3m2f_ca_w_0_140_s_0_210=1.55e-04 mcm3m2f_cc_w_0_140_s_0_210=1.03e-10 mcm3m2f_cf_w_0_140_s_0_210=1.25e-11
+  mcm3m2f_ca_w_0_140_s_0_280=1.55e-04 mcm3m2f_cc_w_0_140_s_0_280=8.50e-11 mcm3m2f_cf_w_0_140_s_0_280=1.67e-11
+  mcm3m2f_ca_w_0_140_s_0_350=1.55e-04 mcm3m2f_cc_w_0_140_s_0_350=7.00e-11 mcm3m2f_cf_w_0_140_s_0_350=2.07e-11
+  mcm3m2f_ca_w_0_140_s_0_420=1.55e-04 mcm3m2f_cc_w_0_140_s_0_420=5.74e-11 mcm3m2f_cf_w_0_140_s_0_420=2.46e-11
+  mcm3m2f_ca_w_0_140_s_0_560=1.55e-04 mcm3m2f_cc_w_0_140_s_0_560=4.03e-11 mcm3m2f_cf_w_0_140_s_0_560=3.10e-11
+  mcm3m2f_ca_w_0_140_s_0_840=1.55e-04 mcm3m2f_cc_w_0_140_s_0_840=2.25e-11 mcm3m2f_cf_w_0_140_s_0_840=4.10e-11
+  mcm3m2f_ca_w_0_140_s_1_540=1.55e-04 mcm3m2f_cc_w_0_140_s_1_540=6.71e-12 mcm3m2f_cf_w_0_140_s_1_540=5.34e-11
+  mcm3m2f_ca_w_0_140_s_3_500=1.55e-04 mcm3m2f_cc_w_0_140_s_3_500=3.90e-13 mcm3m2f_cf_w_0_140_s_3_500=5.96e-11
+  mcm3m2f_ca_w_1_120_s_0_140=1.55e-04 mcm3m2f_cc_w_1_120_s_0_140=1.26e-10 mcm3m2f_cf_w_1_120_s_0_140=7.88e-12
+  mcm3m2f_ca_w_1_120_s_0_175=1.55e-04 mcm3m2f_cc_w_1_120_s_0_175=1.20e-10 mcm3m2f_cf_w_1_120_s_0_175=1.02e-11
+  mcm3m2f_ca_w_1_120_s_0_210=1.55e-04 mcm3m2f_cc_w_1_120_s_0_210=1.11e-10 mcm3m2f_cf_w_1_120_s_0_210=1.25e-11
+  mcm3m2f_ca_w_1_120_s_0_280=1.55e-04 mcm3m2f_cc_w_1_120_s_0_280=9.18e-11 mcm3m2f_cf_w_1_120_s_0_280=1.68e-11
+  mcm3m2f_ca_w_1_120_s_0_350=1.55e-04 mcm3m2f_cc_w_1_120_s_0_350=7.51e-11 mcm3m2f_cf_w_1_120_s_0_350=2.08e-11
+  mcm3m2f_ca_w_1_120_s_0_420=1.55e-04 mcm3m2f_cc_w_1_120_s_0_420=6.19e-11 mcm3m2f_cf_w_1_120_s_0_420=2.45e-11
+  mcm3m2f_ca_w_1_120_s_0_560=1.55e-04 mcm3m2f_cc_w_1_120_s_0_560=4.37e-11 mcm3m2f_cf_w_1_120_s_0_560=3.11e-11
+  mcm3m2f_ca_w_1_120_s_0_840=1.55e-04 mcm3m2f_cc_w_1_120_s_0_840=2.49e-11 mcm3m2f_cf_w_1_120_s_0_840=4.11e-11
+  mcm3m2f_ca_w_1_120_s_1_540=1.55e-04 mcm3m2f_cc_w_1_120_s_1_540=7.78e-12 mcm3m2f_cf_w_1_120_s_1_540=5.42e-11
+  mcm3m2f_ca_w_1_120_s_3_500=1.55e-04 mcm3m2f_cc_w_1_120_s_3_500=4.70e-13 mcm3m2f_cf_w_1_120_s_3_500=6.13e-11
+  mcm3m2d_ca_w_0_140_s_0_140=1.59e-04 mcm3m2d_cc_w_0_140_s_0_140=1.18e-10 mcm3m2d_cf_w_0_140_s_0_140=8.06e-12
+  mcm3m2d_ca_w_0_140_s_0_175=1.59e-04 mcm3m2d_cc_w_0_140_s_0_175=1.10e-10 mcm3m2d_cf_w_0_140_s_0_175=1.05e-11
+  mcm3m2d_ca_w_0_140_s_0_210=1.59e-04 mcm3m2d_cc_w_0_140_s_0_210=1.03e-10 mcm3m2d_cf_w_0_140_s_0_210=1.28e-11
+  mcm3m2d_ca_w_0_140_s_0_280=1.59e-04 mcm3m2d_cc_w_0_140_s_0_280=8.44e-11 mcm3m2d_cf_w_0_140_s_0_280=1.72e-11
+  mcm3m2d_ca_w_0_140_s_0_350=1.59e-04 mcm3m2d_cc_w_0_140_s_0_350=6.92e-11 mcm3m2d_cf_w_0_140_s_0_350=2.13e-11
+  mcm3m2d_ca_w_0_140_s_0_420=1.59e-04 mcm3m2d_cc_w_0_140_s_0_420=5.66e-11 mcm3m2d_cf_w_0_140_s_0_420=2.53e-11
+  mcm3m2d_ca_w_0_140_s_0_560=1.59e-04 mcm3m2d_cc_w_0_140_s_0_560=3.93e-11 mcm3m2d_cf_w_0_140_s_0_560=3.19e-11
+  mcm3m2d_ca_w_0_140_s_0_840=1.59e-04 mcm3m2d_cc_w_0_140_s_0_840=2.15e-11 mcm3m2d_cf_w_0_140_s_0_840=4.22e-11
+  mcm3m2d_ca_w_0_140_s_1_540=1.59e-04 mcm3m2d_cc_w_0_140_s_1_540=5.95e-12 mcm3m2d_cf_w_0_140_s_1_540=5.45e-11
+  mcm3m2d_ca_w_0_140_s_3_500=1.59e-04 mcm3m2d_cc_w_0_140_s_3_500=2.95e-13 mcm3m2d_cf_w_0_140_s_3_500=6.02e-11
+  mcm3m2d_ca_w_1_120_s_0_140=1.59e-04 mcm3m2d_cc_w_1_120_s_0_140=1.25e-10 mcm3m2d_cf_w_1_120_s_0_140=8.09e-12
+  mcm3m2d_ca_w_1_120_s_0_175=1.59e-04 mcm3m2d_cc_w_1_120_s_0_175=1.19e-10 mcm3m2d_cf_w_1_120_s_0_175=1.05e-11
+  mcm3m2d_ca_w_1_120_s_0_210=1.59e-04 mcm3m2d_cc_w_1_120_s_0_210=1.09e-10 mcm3m2d_cf_w_1_120_s_0_210=1.28e-11
+  mcm3m2d_ca_w_1_120_s_0_280=1.59e-04 mcm3m2d_cc_w_1_120_s_0_280=9.03e-11 mcm3m2d_cf_w_1_120_s_0_280=1.73e-11
+  mcm3m2d_ca_w_1_120_s_0_350=1.59e-04 mcm3m2d_cc_w_1_120_s_0_350=7.35e-11 mcm3m2d_cf_w_1_120_s_0_350=2.14e-11
+  mcm3m2d_ca_w_1_120_s_0_420=1.59e-04 mcm3m2d_cc_w_1_120_s_0_420=6.03e-11 mcm3m2d_cf_w_1_120_s_0_420=2.53e-11
+  mcm3m2d_ca_w_1_120_s_0_560=1.59e-04 mcm3m2d_cc_w_1_120_s_0_560=4.22e-11 mcm3m2d_cf_w_1_120_s_0_560=3.20e-11
+  mcm3m2d_ca_w_1_120_s_0_840=1.59e-04 mcm3m2d_cc_w_1_120_s_0_840=2.33e-11 mcm3m2d_cf_w_1_120_s_0_840=4.24e-11
+  mcm3m2d_ca_w_1_120_s_1_540=1.59e-04 mcm3m2d_cc_w_1_120_s_1_540=6.68e-12 mcm3m2d_cf_w_1_120_s_1_540=5.53e-11
+  mcm3m2d_ca_w_1_120_s_3_500=1.59e-04 mcm3m2d_cc_w_1_120_s_3_500=3.55e-13 mcm3m2d_cf_w_1_120_s_3_500=6.17e-11
+  mcm3m2p1_ca_w_0_140_s_0_140=1.67e-04 mcm3m2p1_cc_w_0_140_s_0_140=1.17e-10 mcm3m2p1_cf_w_0_140_s_0_140=8.50e-12
+  mcm3m2p1_ca_w_0_140_s_0_175=1.67e-04 mcm3m2p1_cc_w_0_140_s_0_175=1.09e-10 mcm3m2p1_cf_w_0_140_s_0_175=1.11e-11
+  mcm3m2p1_ca_w_0_140_s_0_210=1.67e-04 mcm3m2p1_cc_w_0_140_s_0_210=1.02e-10 mcm3m2p1_cf_w_0_140_s_0_210=1.35e-11
+  mcm3m2p1_ca_w_0_140_s_0_280=1.67e-04 mcm3m2p1_cc_w_0_140_s_0_280=8.31e-11 mcm3m2p1_cf_w_0_140_s_0_280=1.82e-11
+  mcm3m2p1_ca_w_0_140_s_0_350=1.67e-04 mcm3m2p1_cc_w_0_140_s_0_350=6.77e-11 mcm3m2p1_cf_w_0_140_s_0_350=2.25e-11
+  mcm3m2p1_ca_w_0_140_s_0_420=1.67e-04 mcm3m2p1_cc_w_0_140_s_0_420=5.46e-11 mcm3m2p1_cf_w_0_140_s_0_420=2.67e-11
+  mcm3m2p1_ca_w_0_140_s_0_560=1.67e-04 mcm3m2p1_cc_w_0_140_s_0_560=3.74e-11 mcm3m2p1_cf_w_0_140_s_0_560=3.38e-11
+  mcm3m2p1_ca_w_0_140_s_0_840=1.67e-04 mcm3m2p1_cc_w_0_140_s_0_840=1.96e-11 mcm3m2p1_cf_w_0_140_s_0_840=4.45e-11
+  mcm3m2p1_ca_w_0_140_s_1_540=1.67e-04 mcm3m2p1_cc_w_0_140_s_1_540=4.66e-12 mcm3m2p1_cf_w_0_140_s_1_540=5.69e-11
+  mcm3m2p1_ca_w_0_140_s_3_500=1.67e-04 mcm3m2p1_cc_w_0_140_s_3_500=1.95e-13 mcm3m2p1_cf_w_0_140_s_3_500=6.15e-11
+  mcm3m2p1_ca_w_1_120_s_0_140=1.67e-04 mcm3m2p1_cc_w_1_120_s_0_140=1.23e-10 mcm3m2p1_cf_w_1_120_s_0_140=8.56e-12
+  mcm3m2p1_ca_w_1_120_s_0_175=1.67e-04 mcm3m2p1_cc_w_1_120_s_0_175=1.16e-10 mcm3m2p1_cf_w_1_120_s_0_175=1.11e-11
+  mcm3m2p1_ca_w_1_120_s_0_210=1.67e-04 mcm3m2p1_cc_w_1_120_s_0_210=1.06e-10 mcm3m2p1_cf_w_1_120_s_0_210=1.36e-11
+  mcm3m2p1_ca_w_1_120_s_0_280=1.67e-04 mcm3m2p1_cc_w_1_120_s_0_280=8.71e-11 mcm3m2p1_cf_w_1_120_s_0_280=1.83e-11
+  mcm3m2p1_ca_w_1_120_s_0_350=1.67e-04 mcm3m2p1_cc_w_1_120_s_0_350=7.08e-11 mcm3m2p1_cf_w_1_120_s_0_350=2.26e-11
+  mcm3m2p1_ca_w_1_120_s_0_420=1.67e-04 mcm3m2p1_cc_w_1_120_s_0_420=5.77e-11 mcm3m2p1_cf_w_1_120_s_0_420=2.68e-11
+  mcm3m2p1_ca_w_1_120_s_0_560=1.67e-04 mcm3m2p1_cc_w_1_120_s_0_560=3.93e-11 mcm3m2p1_cf_w_1_120_s_0_560=3.39e-11
+  mcm3m2p1_ca_w_1_120_s_0_840=1.67e-04 mcm3m2p1_cc_w_1_120_s_0_840=2.06e-11 mcm3m2p1_cf_w_1_120_s_0_840=4.47e-11
+  mcm3m2p1_ca_w_1_120_s_1_540=1.67e-04 mcm3m2p1_cc_w_1_120_s_1_540=5.01e-12 mcm3m2p1_cf_w_1_120_s_1_540=5.74e-11
+  mcm3m2p1_ca_w_1_120_s_3_500=1.67e-04 mcm3m2p1_cc_w_1_120_s_3_500=1.80e-13 mcm3m2p1_cf_w_1_120_s_3_500=6.25e-11
+  mcm3m2l1_ca_w_0_140_s_0_140=1.83e-04 mcm3m2l1_cc_w_0_140_s_0_140=1.13e-10 mcm3m2l1_cf_w_0_140_s_0_140=9.36e-12
+  mcm3m2l1_ca_w_0_140_s_0_175=1.83e-04 mcm3m2l1_cc_w_0_140_s_0_175=1.08e-10 mcm3m2l1_cf_w_0_140_s_0_175=1.22e-11
+  mcm3m2l1_ca_w_0_140_s_0_210=1.83e-04 mcm3m2l1_cc_w_0_140_s_0_210=9.95e-11 mcm3m2l1_cf_w_0_140_s_0_210=1.49e-11
+  mcm3m2l1_ca_w_0_140_s_0_280=1.83e-04 mcm3m2l1_cc_w_0_140_s_0_280=8.10e-11 mcm3m2l1_cf_w_0_140_s_0_280=2.01e-11
+  mcm3m2l1_ca_w_0_140_s_0_350=1.83e-04 mcm3m2l1_cc_w_0_140_s_0_350=6.51e-11 mcm3m2l1_cf_w_0_140_s_0_350=2.50e-11
+  mcm3m2l1_ca_w_0_140_s_0_420=1.83e-04 mcm3m2l1_cc_w_0_140_s_0_420=5.18e-11 mcm3m2l1_cf_w_0_140_s_0_420=2.96e-11
+  mcm3m2l1_ca_w_0_140_s_0_560=1.83e-04 mcm3m2l1_cc_w_0_140_s_0_560=3.43e-11 mcm3m2l1_cf_w_0_140_s_0_560=3.75e-11
+  mcm3m2l1_ca_w_0_140_s_0_840=1.83e-04 mcm3m2l1_cc_w_0_140_s_0_840=1.65e-11 mcm3m2l1_cf_w_0_140_s_0_840=4.90e-11
+  mcm3m2l1_ca_w_0_140_s_1_540=1.83e-04 mcm3m2l1_cc_w_0_140_s_1_540=3.03e-12 mcm3m2l1_cf_w_0_140_s_1_540=6.07e-11
+  mcm3m2l1_ca_w_0_140_s_3_500=1.83e-04 mcm3m2l1_cc_w_0_140_s_3_500=1.10e-13 mcm3m2l1_cf_w_0_140_s_3_500=6.42e-11
+  mcm3m2l1_ca_w_1_120_s_0_140=1.83e-04 mcm3m2l1_cc_w_1_120_s_0_140=1.18e-10 mcm3m2l1_cf_w_1_120_s_0_140=9.39e-12
+  mcm3m2l1_ca_w_1_120_s_0_175=1.83e-04 mcm3m2l1_cc_w_1_120_s_0_175=1.12e-10 mcm3m2l1_cf_w_1_120_s_0_175=1.22e-11
+  mcm3m2l1_ca_w_1_120_s_0_210=1.83e-04 mcm3m2l1_cc_w_1_120_s_0_210=1.02e-10 mcm3m2l1_cf_w_1_120_s_0_210=1.50e-11
+  mcm3m2l1_ca_w_1_120_s_0_280=1.83e-04 mcm3m2l1_cc_w_1_120_s_0_280=8.27e-11 mcm3m2l1_cf_w_1_120_s_0_280=2.02e-11
+  mcm3m2l1_ca_w_1_120_s_0_350=1.83e-04 mcm3m2l1_cc_w_1_120_s_0_350=6.66e-11 mcm3m2l1_cf_w_1_120_s_0_350=2.51e-11
+  mcm3m2l1_ca_w_1_120_s_0_420=1.83e-04 mcm3m2l1_cc_w_1_120_s_0_420=5.33e-11 mcm3m2l1_cf_w_1_120_s_0_420=2.97e-11
+  mcm3m2l1_ca_w_1_120_s_0_560=1.83e-04 mcm3m2l1_cc_w_1_120_s_0_560=3.51e-11 mcm3m2l1_cf_w_1_120_s_0_560=3.76e-11
+  mcm3m2l1_ca_w_1_120_s_0_840=1.83e-04 mcm3m2l1_cc_w_1_120_s_0_840=1.70e-11 mcm3m2l1_cf_w_1_120_s_0_840=4.92e-11
+  mcm3m2l1_ca_w_1_120_s_1_540=1.83e-04 mcm3m2l1_cc_w_1_120_s_1_540=3.15e-12 mcm3m2l1_cf_w_1_120_s_1_540=6.14e-11
+  mcm3m2l1_ca_w_1_120_s_3_500=1.83e-04 mcm3m2l1_cc_w_1_120_s_3_500=5.00e-14 mcm3m2l1_cf_w_1_120_s_3_500=6.47e-11
+  mcm3m2m1_ca_w_0_140_s_0_140=4.44e-04 mcm3m2m1_cc_w_0_140_s_0_140=9.86e-11 mcm3m2m1_cf_w_0_140_s_0_140=2.11e-11
+  mcm3m2m1_ca_w_0_140_s_0_175=4.44e-04 mcm3m2m1_cc_w_0_140_s_0_175=9.13e-11 mcm3m2m1_cf_w_0_140_s_0_175=2.84e-11
+  mcm3m2m1_ca_w_0_140_s_0_210=4.44e-04 mcm3m2m1_cc_w_0_140_s_0_210=8.25e-11 mcm3m2m1_cf_w_0_140_s_0_210=3.51e-11
+  mcm3m2m1_ca_w_0_140_s_0_280=4.44e-04 mcm3m2m1_cc_w_0_140_s_0_280=6.39e-11 mcm3m2m1_cf_w_0_140_s_0_280=4.70e-11
+  mcm3m2m1_ca_w_0_140_s_0_350=4.44e-04 mcm3m2m1_cc_w_0_140_s_0_350=4.79e-11 mcm3m2m1_cf_w_0_140_s_0_350=5.73e-11
+  mcm3m2m1_ca_w_0_140_s_0_420=4.44e-04 mcm3m2m1_cc_w_0_140_s_0_420=3.54e-11 mcm3m2m1_cf_w_0_140_s_0_420=6.59e-11
+  mcm3m2m1_ca_w_0_140_s_0_560=4.44e-04 mcm3m2m1_cc_w_0_140_s_0_560=1.95e-11 mcm3m2m1_cf_w_0_140_s_0_560=7.87e-11
+  mcm3m2m1_ca_w_0_140_s_0_840=4.44e-04 mcm3m2m1_cc_w_0_140_s_0_840=6.23e-12 mcm3m2m1_cf_w_0_140_s_0_840=9.19e-11
+  mcm3m2m1_ca_w_0_140_s_1_540=4.44e-04 mcm3m2m1_cc_w_0_140_s_1_540=4.70e-13 mcm3m2m1_cf_w_0_140_s_1_540=9.97e-11
+  mcm3m2m1_ca_w_0_140_s_3_500=4.44e-04 mcm3m2m1_cc_w_0_140_s_3_500=0.00e+00 mcm3m2m1_cf_w_0_140_s_3_500=1.01e-10
+  mcm3m2m1_ca_w_1_120_s_0_140=4.44e-04 mcm3m2m1_cc_w_1_120_s_0_140=9.87e-11 mcm3m2m1_cf_w_1_120_s_0_140=2.10e-11
+  mcm3m2m1_ca_w_1_120_s_0_175=4.44e-04 mcm3m2m1_cc_w_1_120_s_0_175=9.22e-11 mcm3m2m1_cf_w_1_120_s_0_175=2.84e-11
+  mcm3m2m1_ca_w_1_120_s_0_210=4.44e-04 mcm3m2m1_cc_w_1_120_s_0_210=8.34e-11 mcm3m2m1_cf_w_1_120_s_0_210=3.52e-11
+  mcm3m2m1_ca_w_1_120_s_0_280=4.44e-04 mcm3m2m1_cc_w_1_120_s_0_280=6.39e-11 mcm3m2m1_cf_w_1_120_s_0_280=4.71e-11
+  mcm3m2m1_ca_w_1_120_s_0_350=4.44e-04 mcm3m2m1_cc_w_1_120_s_0_350=4.83e-11 mcm3m2m1_cf_w_1_120_s_0_350=5.73e-11
+  mcm3m2m1_ca_w_1_120_s_0_420=4.44e-04 mcm3m2m1_cc_w_1_120_s_0_420=3.57e-11 mcm3m2m1_cf_w_1_120_s_0_420=6.60e-11
+  mcm3m2m1_ca_w_1_120_s_0_560=4.44e-04 mcm3m2m1_cc_w_1_120_s_0_560=1.97e-11 mcm3m2m1_cf_w_1_120_s_0_560=7.87e-11
+  mcm3m2m1_ca_w_1_120_s_0_840=4.44e-04 mcm3m2m1_cc_w_1_120_s_0_840=6.30e-12 mcm3m2m1_cf_w_1_120_s_0_840=9.22e-11
+  mcm3m2m1_ca_w_1_120_s_1_540=4.44e-04 mcm3m2m1_cc_w_1_120_s_1_540=5.00e-13 mcm3m2m1_cf_w_1_120_s_1_540=9.97e-11
+  mcm3m2m1_ca_w_1_120_s_3_500=4.44e-04 mcm3m2m1_cc_w_1_120_s_3_500=5.00e-14 mcm3m2m1_cf_w_1_120_s_3_500=1.02e-10
+  mcm4m2f_ca_w_0_140_s_0_140=4.88e-05 mcm4m2f_cc_w_0_140_s_0_140=1.28e-10 mcm4m2f_cf_w_0_140_s_0_140=2.64e-12
+  mcm4m2f_ca_w_0_140_s_0_175=4.88e-05 mcm4m2f_cc_w_0_140_s_0_175=1.21e-10 mcm4m2f_cf_w_0_140_s_0_175=3.47e-12
+  mcm4m2f_ca_w_0_140_s_0_210=4.88e-05 mcm4m2f_cc_w_0_140_s_0_210=1.15e-10 mcm4m2f_cf_w_0_140_s_0_210=4.32e-12
+  mcm4m2f_ca_w_0_140_s_0_280=4.88e-05 mcm4m2f_cc_w_0_140_s_0_280=9.71e-11 mcm4m2f_cf_w_0_140_s_0_280=5.96e-12
+  mcm4m2f_ca_w_0_140_s_0_350=4.88e-05 mcm4m2f_cc_w_0_140_s_0_350=8.25e-11 mcm4m2f_cf_w_0_140_s_0_350=7.57e-12
+  mcm4m2f_ca_w_0_140_s_0_420=4.88e-05 mcm4m2f_cc_w_0_140_s_0_420=7.01e-11 mcm4m2f_cf_w_0_140_s_0_420=9.22e-12
+  mcm4m2f_ca_w_0_140_s_0_560=4.88e-05 mcm4m2f_cc_w_0_140_s_0_560=5.35e-11 mcm4m2f_cf_w_0_140_s_0_560=1.22e-11
+  mcm4m2f_ca_w_0_140_s_0_840=4.88e-05 mcm4m2f_cc_w_0_140_s_0_840=3.54e-11 mcm4m2f_cf_w_0_140_s_0_840=1.78e-11
+  mcm4m2f_ca_w_0_140_s_1_540=4.88e-05 mcm4m2f_cc_w_0_140_s_1_540=1.59e-11 mcm4m2f_cf_w_0_140_s_1_540=2.82e-11
+  mcm4m2f_ca_w_0_140_s_3_500=4.88e-05 mcm4m2f_cc_w_0_140_s_3_500=2.31e-12 mcm4m2f_cf_w_0_140_s_3_500=3.93e-11
+  mcm4m2f_ca_w_1_120_s_0_140=4.88e-05 mcm4m2f_cc_w_1_120_s_0_140=1.44e-10 mcm4m2f_cf_w_1_120_s_0_140=2.68e-12
+  mcm4m2f_ca_w_1_120_s_0_175=4.88e-05 mcm4m2f_cc_w_1_120_s_0_175=1.37e-10 mcm4m2f_cf_w_1_120_s_0_175=3.52e-12
+  mcm4m2f_ca_w_1_120_s_0_210=4.88e-05 mcm4m2f_cc_w_1_120_s_0_210=1.29e-10 mcm4m2f_cf_w_1_120_s_0_210=4.35e-12
+  mcm4m2f_ca_w_1_120_s_0_280=4.88e-05 mcm4m2f_cc_w_1_120_s_0_280=1.09e-10 mcm4m2f_cf_w_1_120_s_0_280=5.99e-12
+  mcm4m2f_ca_w_1_120_s_0_350=4.88e-05 mcm4m2f_cc_w_1_120_s_0_350=9.22e-11 mcm4m2f_cf_w_1_120_s_0_350=7.63e-12
+  mcm4m2f_ca_w_1_120_s_0_420=4.88e-05 mcm4m2f_cc_w_1_120_s_0_420=7.88e-11 mcm4m2f_cf_w_1_120_s_0_420=9.23e-12
+  mcm4m2f_ca_w_1_120_s_0_560=4.88e-05 mcm4m2f_cc_w_1_120_s_0_560=6.03e-11 mcm4m2f_cf_w_1_120_s_0_560=1.23e-11
+  mcm4m2f_ca_w_1_120_s_0_840=4.88e-05 mcm4m2f_cc_w_1_120_s_0_840=3.98e-11 mcm4m2f_cf_w_1_120_s_0_840=1.79e-11
+  mcm4m2f_ca_w_1_120_s_1_540=4.88e-05 mcm4m2f_cc_w_1_120_s_1_540=1.81e-11 mcm4m2f_cf_w_1_120_s_1_540=2.89e-11
+  mcm4m2f_ca_w_1_120_s_3_500=4.88e-05 mcm4m2f_cc_w_1_120_s_3_500=2.66e-12 mcm4m2f_cf_w_1_120_s_3_500=4.13e-11
+  mcm4m2d_ca_w_0_140_s_0_140=5.26e-05 mcm4m2d_cc_w_0_140_s_0_140=1.28e-10 mcm4m2d_cf_w_0_140_s_0_140=2.85e-12
+  mcm4m2d_ca_w_0_140_s_0_175=5.26e-05 mcm4m2d_cc_w_0_140_s_0_175=1.21e-10 mcm4m2d_cf_w_0_140_s_0_175=3.75e-12
+  mcm4m2d_ca_w_0_140_s_0_210=5.26e-05 mcm4m2d_cc_w_0_140_s_0_210=1.14e-10 mcm4m2d_cf_w_0_140_s_0_210=4.66e-12
+  mcm4m2d_ca_w_0_140_s_0_280=5.26e-05 mcm4m2d_cc_w_0_140_s_0_280=9.65e-11 mcm4m2d_cf_w_0_140_s_0_280=6.43e-12
+  mcm4m2d_ca_w_0_140_s_0_350=5.26e-05 mcm4m2d_cc_w_0_140_s_0_350=8.18e-11 mcm4m2d_cf_w_0_140_s_0_350=8.17e-12
+  mcm4m2d_ca_w_0_140_s_0_420=5.26e-05 mcm4m2d_cc_w_0_140_s_0_420=6.93e-11 mcm4m2d_cf_w_0_140_s_0_420=9.93e-12
+  mcm4m2d_ca_w_0_140_s_0_560=5.26e-05 mcm4m2d_cc_w_0_140_s_0_560=5.25e-11 mcm4m2d_cf_w_0_140_s_0_560=1.32e-11
+  mcm4m2d_ca_w_0_140_s_0_840=5.26e-05 mcm4m2d_cc_w_0_140_s_0_840=3.42e-11 mcm4m2d_cf_w_0_140_s_0_840=1.91e-11
+  mcm4m2d_ca_w_0_140_s_1_540=5.26e-05 mcm4m2d_cc_w_0_140_s_1_540=1.48e-11 mcm4m2d_cf_w_0_140_s_1_540=3.00e-11
+  mcm4m2d_ca_w_0_140_s_3_500=5.26e-05 mcm4m2d_cc_w_0_140_s_3_500=1.90e-12 mcm4m2d_cf_w_0_140_s_3_500=4.08e-11
+  mcm4m2d_ca_w_1_120_s_0_140=5.26e-05 mcm4m2d_cc_w_1_120_s_0_140=1.42e-10 mcm4m2d_cf_w_1_120_s_0_140=2.89e-12
+  mcm4m2d_ca_w_1_120_s_0_175=5.26e-05 mcm4m2d_cc_w_1_120_s_0_175=1.36e-10 mcm4m2d_cf_w_1_120_s_0_175=3.79e-12
+  mcm4m2d_ca_w_1_120_s_0_210=5.26e-05 mcm4m2d_cc_w_1_120_s_0_210=1.27e-10 mcm4m2d_cf_w_1_120_s_0_210=4.70e-12
+  mcm4m2d_ca_w_1_120_s_0_280=5.26e-05 mcm4m2d_cc_w_1_120_s_0_280=1.07e-10 mcm4m2d_cf_w_1_120_s_0_280=6.47e-12
+  mcm4m2d_ca_w_1_120_s_0_350=5.26e-05 mcm4m2d_cc_w_1_120_s_0_350=9.06e-11 mcm4m2d_cf_w_1_120_s_0_350=8.25e-12
+  mcm4m2d_ca_w_1_120_s_0_420=5.26e-05 mcm4m2d_cc_w_1_120_s_0_420=7.71e-11 mcm4m2d_cf_w_1_120_s_0_420=9.96e-12
+  mcm4m2d_ca_w_1_120_s_0_560=5.26e-05 mcm4m2d_cc_w_1_120_s_0_560=5.87e-11 mcm4m2d_cf_w_1_120_s_0_560=1.33e-11
+  mcm4m2d_ca_w_1_120_s_0_840=5.26e-05 mcm4m2d_cc_w_1_120_s_0_840=3.82e-11 mcm4m2d_cf_w_1_120_s_0_840=1.93e-11
+  mcm4m2d_ca_w_1_120_s_1_540=5.26e-05 mcm4m2d_cc_w_1_120_s_1_540=1.66e-11 mcm4m2d_cf_w_1_120_s_1_540=3.07e-11
+  mcm4m2d_ca_w_1_120_s_3_500=5.26e-05 mcm4m2d_cc_w_1_120_s_3_500=2.16e-12 mcm4m2d_cf_w_1_120_s_3_500=4.26e-11
+  mcm4m2p1_ca_w_0_140_s_0_140=6.08e-05 mcm4m2p1_cc_w_0_140_s_0_140=1.28e-10 mcm4m2p1_cf_w_0_140_s_0_140=3.30e-12
+  mcm4m2p1_ca_w_0_140_s_0_175=6.08e-05 mcm4m2p1_cc_w_0_140_s_0_175=1.20e-10 mcm4m2p1_cf_w_0_140_s_0_175=4.34e-12
+  mcm4m2p1_ca_w_0_140_s_0_210=6.08e-05 mcm4m2p1_cc_w_0_140_s_0_210=1.13e-10 mcm4m2p1_cf_w_0_140_s_0_210=5.39e-12
+  mcm4m2p1_ca_w_0_140_s_0_280=6.08e-05 mcm4m2p1_cc_w_0_140_s_0_280=9.50e-11 mcm4m2p1_cf_w_0_140_s_0_280=7.44e-12
+  mcm4m2p1_ca_w_0_140_s_0_350=6.08e-05 mcm4m2p1_cc_w_0_140_s_0_350=8.03e-11 mcm4m2p1_cf_w_0_140_s_0_350=9.44e-12
+  mcm4m2p1_ca_w_0_140_s_0_420=6.08e-05 mcm4m2p1_cc_w_0_140_s_0_420=6.76e-11 mcm4m2p1_cf_w_0_140_s_0_420=1.15e-11
+  mcm4m2p1_ca_w_0_140_s_0_560=6.08e-05 mcm4m2p1_cc_w_0_140_s_0_560=5.07e-11 mcm4m2p1_cf_w_0_140_s_0_560=1.51e-11
+  mcm4m2p1_ca_w_0_140_s_0_840=6.08e-05 mcm4m2p1_cc_w_0_140_s_0_840=3.21e-11 mcm4m2p1_cf_w_0_140_s_0_840=2.18e-11
+  mcm4m2p1_ca_w_0_140_s_1_540=6.08e-05 mcm4m2p1_cc_w_0_140_s_1_540=1.29e-11 mcm4m2p1_cf_w_0_140_s_1_540=3.34e-11
+  mcm4m2p1_ca_w_0_140_s_3_500=6.08e-05 mcm4m2p1_cc_w_0_140_s_3_500=1.32e-12 mcm4m2p1_cf_w_0_140_s_3_500=4.35e-11
+  mcm4m2p1_ca_w_1_120_s_0_140=6.08e-05 mcm4m2p1_cc_w_1_120_s_0_140=1.39e-10 mcm4m2p1_cf_w_1_120_s_0_140=3.38e-12
+  mcm4m2p1_ca_w_1_120_s_0_175=6.08e-05 mcm4m2p1_cc_w_1_120_s_0_175=1.33e-10 mcm4m2p1_cf_w_1_120_s_0_175=4.44e-12
+  mcm4m2p1_ca_w_1_120_s_0_210=6.08e-05 mcm4m2p1_cc_w_1_120_s_0_210=1.24e-10 mcm4m2p1_cf_w_1_120_s_0_210=5.48e-12
+  mcm4m2p1_ca_w_1_120_s_0_280=6.08e-05 mcm4m2p1_cc_w_1_120_s_0_280=1.04e-10 mcm4m2p1_cf_w_1_120_s_0_280=7.50e-12
+  mcm4m2p1_ca_w_1_120_s_0_350=6.08e-05 mcm4m2p1_cc_w_1_120_s_0_350=8.74e-11 mcm4m2p1_cf_w_1_120_s_0_350=9.53e-12
+  mcm4m2p1_ca_w_1_120_s_0_420=6.08e-05 mcm4m2p1_cc_w_1_120_s_0_420=7.45e-11 mcm4m2p1_cf_w_1_120_s_0_420=1.15e-11
+  mcm4m2p1_ca_w_1_120_s_0_560=6.08e-05 mcm4m2p1_cc_w_1_120_s_0_560=5.57e-11 mcm4m2p1_cf_w_1_120_s_0_560=1.53e-11
+  mcm4m2p1_ca_w_1_120_s_0_840=6.08e-05 mcm4m2p1_cc_w_1_120_s_0_840=3.54e-11 mcm4m2p1_cf_w_1_120_s_0_840=2.21e-11
+  mcm4m2p1_ca_w_1_120_s_1_540=6.08e-05 mcm4m2p1_cc_w_1_120_s_1_540=1.43e-11 mcm4m2p1_cf_w_1_120_s_1_540=3.42e-11
+  mcm4m2p1_ca_w_1_120_s_3_500=6.08e-05 mcm4m2p1_cc_w_1_120_s_3_500=1.51e-12 mcm4m2p1_cf_w_1_120_s_3_500=4.52e-11
+  mcm4m2l1_ca_w_0_140_s_0_140=7.75e-05 mcm4m2l1_cc_w_0_140_s_0_140=1.24e-10 mcm4m2l1_cf_w_0_140_s_0_140=4.15e-12
+  mcm4m2l1_ca_w_0_140_s_0_175=7.75e-05 mcm4m2l1_cc_w_0_140_s_0_175=1.19e-10 mcm4m2l1_cf_w_0_140_s_0_175=5.49e-12
+  mcm4m2l1_ca_w_0_140_s_0_210=7.75e-05 mcm4m2l1_cc_w_0_140_s_0_210=1.11e-10 mcm4m2l1_cf_w_0_140_s_0_210=6.81e-12
+  mcm4m2l1_ca_w_0_140_s_0_280=7.75e-05 mcm4m2l1_cc_w_0_140_s_0_280=9.28e-11 mcm4m2l1_cf_w_0_140_s_0_280=9.40e-12
+  mcm4m2l1_ca_w_0_140_s_0_350=7.75e-05 mcm4m2l1_cc_w_0_140_s_0_350=7.76e-11 mcm4m2l1_cf_w_0_140_s_0_350=1.19e-11
+  mcm4m2l1_ca_w_0_140_s_0_420=7.75e-05 mcm4m2l1_cc_w_0_140_s_0_420=6.50e-11 mcm4m2l1_cf_w_0_140_s_0_420=1.44e-11
+  mcm4m2l1_ca_w_0_140_s_0_560=7.75e-05 mcm4m2l1_cc_w_0_140_s_0_560=4.75e-11 mcm4m2l1_cf_w_0_140_s_0_560=1.89e-11
+  mcm4m2l1_ca_w_0_140_s_0_840=7.75e-05 mcm4m2l1_cc_w_0_140_s_0_840=2.89e-11 mcm4m2l1_cf_w_0_140_s_0_840=2.68e-11
+  mcm4m2l1_ca_w_0_140_s_1_540=7.75e-05 mcm4m2l1_cc_w_0_140_s_1_540=1.02e-11 mcm4m2l1_cf_w_0_140_s_1_540=3.93e-11
+  mcm4m2l1_ca_w_0_140_s_3_500=7.75e-05 mcm4m2l1_cc_w_0_140_s_3_500=8.00e-13 mcm4m2l1_cf_w_0_140_s_3_500=4.80e-11
+  mcm4m2l1_ca_w_1_120_s_0_140=7.75e-05 mcm4m2l1_cc_w_1_120_s_0_140=1.35e-10 mcm4m2l1_cf_w_1_120_s_0_140=4.19e-12
+  mcm4m2l1_ca_w_1_120_s_0_175=7.75e-05 mcm4m2l1_cc_w_1_120_s_0_175=1.29e-10 mcm4m2l1_cf_w_1_120_s_0_175=5.54e-12
+  mcm4m2l1_ca_w_1_120_s_0_210=7.75e-05 mcm4m2l1_cc_w_1_120_s_0_210=1.20e-10 mcm4m2l1_cf_w_1_120_s_0_210=6.86e-12
+  mcm4m2l1_ca_w_1_120_s_0_280=7.75e-05 mcm4m2l1_cc_w_1_120_s_0_280=1.00e-10 mcm4m2l1_cf_w_1_120_s_0_280=9.44e-12
+  mcm4m2l1_ca_w_1_120_s_0_350=7.75e-05 mcm4m2l1_cc_w_1_120_s_0_350=8.37e-11 mcm4m2l1_cf_w_1_120_s_0_350=1.20e-11
+  mcm4m2l1_ca_w_1_120_s_0_420=7.75e-05 mcm4m2l1_cc_w_1_120_s_0_420=7.02e-11 mcm4m2l1_cf_w_1_120_s_0_420=1.44e-11
+  mcm4m2l1_ca_w_1_120_s_0_560=7.75e-05 mcm4m2l1_cc_w_1_120_s_0_560=5.16e-11 mcm4m2l1_cf_w_1_120_s_0_560=1.90e-11
+  mcm4m2l1_ca_w_1_120_s_0_840=7.75e-05 mcm4m2l1_cc_w_1_120_s_0_840=3.14e-11 mcm4m2l1_cf_w_1_120_s_0_840=2.71e-11
+  mcm4m2l1_ca_w_1_120_s_1_540=7.75e-05 mcm4m2l1_cc_w_1_120_s_1_540=1.14e-11 mcm4m2l1_cf_w_1_120_s_1_540=4.01e-11
+  mcm4m2l1_ca_w_1_120_s_3_500=7.75e-05 mcm4m2l1_cc_w_1_120_s_3_500=9.05e-13 mcm4m2l1_cf_w_1_120_s_3_500=4.97e-11
+  mcm4m2m1_ca_w_0_140_s_0_140=3.38e-04 mcm4m2m1_cc_w_0_140_s_0_140=1.08e-10 mcm4m2m1_cf_w_0_140_s_0_140=1.59e-11
+  mcm4m2m1_ca_w_0_140_s_0_175=3.38e-04 mcm4m2m1_cc_w_0_140_s_0_175=1.02e-10 mcm4m2m1_cf_w_0_140_s_0_175=2.17e-11
+  mcm4m2m1_ca_w_0_140_s_0_210=3.38e-04 mcm4m2m1_cc_w_0_140_s_0_210=9.34e-11 mcm4m2m1_cf_w_0_140_s_0_210=2.70e-11
+  mcm4m2m1_ca_w_0_140_s_0_280=3.38e-04 mcm4m2m1_cc_w_0_140_s_0_280=7.52e-11 mcm4m2m1_cf_w_0_140_s_0_280=3.63e-11
+  mcm4m2m1_ca_w_0_140_s_0_350=3.38e-04 mcm4m2m1_cc_w_0_140_s_0_350=6.02e-11 mcm4m2m1_cf_w_0_140_s_0_350=4.42e-11
+  mcm4m2m1_ca_w_0_140_s_0_420=3.38e-04 mcm4m2m1_cc_w_0_140_s_0_420=4.81e-11 mcm4m2m1_cf_w_0_140_s_0_420=5.09e-11
+  mcm4m2m1_ca_w_0_140_s_0_560=3.38e-04 mcm4m2m1_cc_w_0_140_s_0_560=3.20e-11 mcm4m2m1_cf_w_0_140_s_0_560=6.12e-11
+  mcm4m2m1_ca_w_0_140_s_0_840=3.38e-04 mcm4m2m1_cc_w_0_140_s_0_840=1.62e-11 mcm4m2m1_cf_w_0_140_s_0_840=7.40e-11
+  mcm4m2m1_ca_w_0_140_s_1_540=3.38e-04 mcm4m2m1_cc_w_0_140_s_1_540=3.96e-12 mcm4m2m1_cf_w_0_140_s_1_540=8.62e-11
+  mcm4m2m1_ca_w_0_140_s_3_500=3.38e-04 mcm4m2m1_cc_w_0_140_s_3_500=2.30e-13 mcm4m2m1_cf_w_0_140_s_3_500=9.13e-11
+  mcm4m2m1_ca_w_1_120_s_0_140=3.38e-04 mcm4m2m1_cc_w_1_120_s_0_140=1.17e-10 mcm4m2m1_cf_w_1_120_s_0_140=1.59e-11
+  mcm4m2m1_ca_w_1_120_s_0_175=3.38e-04 mcm4m2m1_cc_w_1_120_s_0_175=1.10e-10 mcm4m2m1_cf_w_1_120_s_0_175=2.17e-11
+  mcm4m2m1_ca_w_1_120_s_0_210=3.38e-04 mcm4m2m1_cc_w_1_120_s_0_210=9.99e-11 mcm4m2m1_cf_w_1_120_s_0_210=2.69e-11
+  mcm4m2m1_ca_w_1_120_s_0_280=3.38e-04 mcm4m2m1_cc_w_1_120_s_0_280=8.10e-11 mcm4m2m1_cf_w_1_120_s_0_280=3.63e-11
+  mcm4m2m1_ca_w_1_120_s_0_350=3.38e-04 mcm4m2m1_cc_w_1_120_s_0_350=6.50e-11 mcm4m2m1_cf_w_1_120_s_0_350=4.42e-11
+  mcm4m2m1_ca_w_1_120_s_0_420=3.38e-04 mcm4m2m1_cc_w_1_120_s_0_420=5.26e-11 mcm4m2m1_cf_w_1_120_s_0_420=5.09e-11
+  mcm4m2m1_ca_w_1_120_s_0_560=3.38e-04 mcm4m2m1_cc_w_1_120_s_0_560=3.54e-11 mcm4m2m1_cf_w_1_120_s_0_560=6.12e-11
+  mcm4m2m1_ca_w_1_120_s_0_840=3.38e-04 mcm4m2m1_cc_w_1_120_s_0_840=1.84e-11 mcm4m2m1_cf_w_1_120_s_0_840=7.43e-11
+  mcm4m2m1_ca_w_1_120_s_1_540=3.38e-04 mcm4m2m1_cc_w_1_120_s_1_540=4.89e-12 mcm4m2m1_cf_w_1_120_s_1_540=8.76e-11
+  mcm4m2m1_ca_w_1_120_s_3_500=3.38e-04 mcm4m2m1_cc_w_1_120_s_3_500=2.85e-13 mcm4m2m1_cf_w_1_120_s_3_500=9.35e-11
+  mcm5m2f_ca_w_0_140_s_0_140=3.68e-05 mcm5m2f_cc_w_0_140_s_0_140=1.29e-10 mcm5m2f_cf_w_0_140_s_0_140=2.01e-12
+  mcm5m2f_ca_w_0_140_s_0_175=3.68e-05 mcm5m2f_cc_w_0_140_s_0_175=1.23e-10 mcm5m2f_cf_w_0_140_s_0_175=2.64e-12
+  mcm5m2f_ca_w_0_140_s_0_210=3.68e-05 mcm5m2f_cc_w_0_140_s_0_210=1.16e-10 mcm5m2f_cf_w_0_140_s_0_210=3.28e-12
+  mcm5m2f_ca_w_0_140_s_0_280=3.68e-05 mcm5m2f_cc_w_0_140_s_0_280=9.92e-11 mcm5m2f_cf_w_0_140_s_0_280=4.55e-12
+  mcm5m2f_ca_w_0_140_s_0_350=3.68e-05 mcm5m2f_cc_w_0_140_s_0_350=8.49e-11 mcm5m2f_cf_w_0_140_s_0_350=5.79e-12
+  mcm5m2f_ca_w_0_140_s_0_420=3.68e-05 mcm5m2f_cc_w_0_140_s_0_420=7.29e-11 mcm5m2f_cf_w_0_140_s_0_420=7.07e-12
+  mcm5m2f_ca_w_0_140_s_0_560=3.68e-05 mcm5m2f_cc_w_0_140_s_0_560=5.65e-11 mcm5m2f_cf_w_0_140_s_0_560=9.42e-12
+  mcm5m2f_ca_w_0_140_s_0_840=3.68e-05 mcm5m2f_cc_w_0_140_s_0_840=3.90e-11 mcm5m2f_cf_w_0_140_s_0_840=1.38e-11
+  mcm5m2f_ca_w_0_140_s_1_540=3.68e-05 mcm5m2f_cc_w_0_140_s_1_540=1.99e-11 mcm5m2f_cf_w_0_140_s_1_540=2.27e-11
+  mcm5m2f_ca_w_0_140_s_3_500=3.68e-05 mcm5m2f_cc_w_0_140_s_3_500=4.43e-12 mcm5m2f_cf_w_0_140_s_3_500=3.44e-11
+  mcm5m2f_ca_w_1_120_s_0_140=3.68e-05 mcm5m2f_cc_w_1_120_s_0_140=1.49e-10 mcm5m2f_cf_w_1_120_s_0_140=2.05e-12
+  mcm5m2f_ca_w_1_120_s_0_175=3.68e-05 mcm5m2f_cc_w_1_120_s_0_175=1.42e-10 mcm5m2f_cf_w_1_120_s_0_175=2.69e-12
+  mcm5m2f_ca_w_1_120_s_0_210=3.68e-05 mcm5m2f_cc_w_1_120_s_0_210=1.34e-10 mcm5m2f_cf_w_1_120_s_0_210=3.33e-12
+  mcm5m2f_ca_w_1_120_s_0_280=3.68e-05 mcm5m2f_cc_w_1_120_s_0_280=1.14e-10 mcm5m2f_cf_w_1_120_s_0_280=4.59e-12
+  mcm5m2f_ca_w_1_120_s_0_350=3.68e-05 mcm5m2f_cc_w_1_120_s_0_350=9.75e-11 mcm5m2f_cf_w_1_120_s_0_350=5.85e-12
+  mcm5m2f_ca_w_1_120_s_0_420=3.68e-05 mcm5m2f_cc_w_1_120_s_0_420=8.46e-11 mcm5m2f_cf_w_1_120_s_0_420=7.05e-12
+  mcm5m2f_ca_w_1_120_s_0_560=3.68e-05 mcm5m2f_cc_w_1_120_s_0_560=6.59e-11 mcm5m2f_cf_w_1_120_s_0_560=9.47e-12
+  mcm5m2f_ca_w_1_120_s_0_840=3.68e-05 mcm5m2f_cc_w_1_120_s_0_840=4.56e-11 mcm5m2f_cf_w_1_120_s_0_840=1.40e-11
+  mcm5m2f_ca_w_1_120_s_1_540=3.68e-05 mcm5m2f_cc_w_1_120_s_1_540=2.35e-11 mcm5m2f_cf_w_1_120_s_1_540=2.32e-11
+  mcm5m2f_ca_w_1_120_s_3_500=3.68e-05 mcm5m2f_cc_w_1_120_s_3_500=5.42e-12 mcm5m2f_cf_w_1_120_s_3_500=3.64e-11
+  mcm5m2d_ca_w_0_140_s_0_140=4.07e-05 mcm5m2d_cc_w_0_140_s_0_140=1.29e-10 mcm5m2d_cf_w_0_140_s_0_140=2.22e-12
+  mcm5m2d_ca_w_0_140_s_0_175=4.07e-05 mcm5m2d_cc_w_0_140_s_0_175=1.22e-10 mcm5m2d_cf_w_0_140_s_0_175=2.92e-12
+  mcm5m2d_ca_w_0_140_s_0_210=4.07e-05 mcm5m2d_cc_w_0_140_s_0_210=1.15e-10 mcm5m2d_cf_w_0_140_s_0_210=3.63e-12
+  mcm5m2d_ca_w_0_140_s_0_280=4.07e-05 mcm5m2d_cc_w_0_140_s_0_280=9.85e-11 mcm5m2d_cf_w_0_140_s_0_280=5.03e-12
+  mcm5m2d_ca_w_0_140_s_0_350=4.07e-05 mcm5m2d_cc_w_0_140_s_0_350=8.38e-11 mcm5m2d_cf_w_0_140_s_0_350=6.38e-12
+  mcm5m2d_ca_w_0_140_s_0_420=4.07e-05 mcm5m2d_cc_w_0_140_s_0_420=7.21e-11 mcm5m2d_cf_w_0_140_s_0_420=7.79e-12
+  mcm5m2d_ca_w_0_140_s_0_560=4.07e-05 mcm5m2d_cc_w_0_140_s_0_560=5.56e-11 mcm5m2d_cf_w_0_140_s_0_560=1.04e-11
+  mcm5m2d_ca_w_0_140_s_0_840=4.07e-05 mcm5m2d_cc_w_0_140_s_0_840=3.79e-11 mcm5m2d_cf_w_0_140_s_0_840=1.51e-11
+  mcm5m2d_ca_w_0_140_s_1_540=4.07e-05 mcm5m2d_cc_w_0_140_s_1_540=1.87e-11 mcm5m2d_cf_w_0_140_s_1_540=2.46e-11
+  mcm5m2d_ca_w_0_140_s_3_500=4.07e-05 mcm5m2d_cc_w_0_140_s_3_500=3.80e-12 mcm5m2d_cf_w_0_140_s_3_500=3.62e-11
+  mcm5m2d_ca_w_1_120_s_0_140=4.07e-05 mcm5m2d_cc_w_1_120_s_0_140=1.47e-10 mcm5m2d_cf_w_1_120_s_0_140=2.28e-12
+  mcm5m2d_ca_w_1_120_s_0_175=4.07e-05 mcm5m2d_cc_w_1_120_s_0_175=1.41e-10 mcm5m2d_cf_w_1_120_s_0_175=2.97e-12
+  mcm5m2d_ca_w_1_120_s_0_210=4.07e-05 mcm5m2d_cc_w_1_120_s_0_210=1.32e-10 mcm5m2d_cf_w_1_120_s_0_210=3.67e-12
+  mcm5m2d_ca_w_1_120_s_0_280=4.07e-05 mcm5m2d_cc_w_1_120_s_0_280=1.13e-10 mcm5m2d_cf_w_1_120_s_0_280=5.06e-12
+  mcm5m2d_ca_w_1_120_s_0_350=4.07e-05 mcm5m2d_cc_w_1_120_s_0_350=9.59e-11 mcm5m2d_cf_w_1_120_s_0_350=6.45e-12
+  mcm5m2d_ca_w_1_120_s_0_420=4.07e-05 mcm5m2d_cc_w_1_120_s_0_420=8.30e-11 mcm5m2d_cf_w_1_120_s_0_420=7.79e-12
+  mcm5m2d_ca_w_1_120_s_0_560=4.07e-05 mcm5m2d_cc_w_1_120_s_0_560=6.44e-11 mcm5m2d_cf_w_1_120_s_0_560=1.04e-11
+  mcm5m2d_ca_w_1_120_s_0_840=4.07e-05 mcm5m2d_cc_w_1_120_s_0_840=4.41e-11 mcm5m2d_cf_w_1_120_s_0_840=1.53e-11
+  mcm5m2d_ca_w_1_120_s_1_540=4.07e-05 mcm5m2d_cc_w_1_120_s_1_540=2.20e-11 mcm5m2d_cf_w_1_120_s_1_540=2.52e-11
+  mcm5m2d_ca_w_1_120_s_3_500=4.07e-05 mcm5m2d_cc_w_1_120_s_3_500=4.67e-12 mcm5m2d_cf_w_1_120_s_3_500=3.82e-11
+  mcm5m2p1_ca_w_0_140_s_0_140=4.89e-05 mcm5m2p1_cc_w_0_140_s_0_140=1.29e-10 mcm5m2p1_cf_w_0_140_s_0_140=2.66e-12
+  mcm5m2p1_ca_w_0_140_s_0_175=4.89e-05 mcm5m2p1_cc_w_0_140_s_0_175=1.22e-10 mcm5m2p1_cf_w_0_140_s_0_175=3.51e-12
+  mcm5m2p1_ca_w_0_140_s_0_210=4.89e-05 mcm5m2p1_cc_w_0_140_s_0_210=1.14e-10 mcm5m2p1_cf_w_0_140_s_0_210=4.36e-12
+  mcm5m2p1_ca_w_0_140_s_0_280=4.89e-05 mcm5m2p1_cc_w_0_140_s_0_280=9.72e-11 mcm5m2p1_cf_w_0_140_s_0_280=6.02e-12
+  mcm5m2p1_ca_w_0_140_s_0_350=4.89e-05 mcm5m2p1_cc_w_0_140_s_0_350=8.19e-11 mcm5m2p1_cf_w_0_140_s_0_350=7.66e-12
+  mcm5m2p1_ca_w_0_140_s_0_420=4.89e-05 mcm5m2p1_cc_w_0_140_s_0_420=7.05e-11 mcm5m2p1_cf_w_0_140_s_0_420=9.31e-12
+  mcm5m2p1_ca_w_0_140_s_0_560=4.89e-05 mcm5m2p1_cc_w_0_140_s_0_560=5.36e-11 mcm5m2p1_cf_w_0_140_s_0_560=1.23e-11
+  mcm5m2p1_ca_w_0_140_s_0_840=4.89e-05 mcm5m2p1_cc_w_0_140_s_0_840=3.57e-11 mcm5m2p1_cf_w_0_140_s_0_840=1.79e-11
+  mcm5m2p1_ca_w_0_140_s_1_540=4.89e-05 mcm5m2p1_cc_w_0_140_s_1_540=1.66e-11 mcm5m2p1_cf_w_0_140_s_1_540=2.83e-11
+  mcm5m2p1_ca_w_0_140_s_3_500=4.89e-05 mcm5m2p1_cc_w_0_140_s_3_500=2.93e-12 mcm5m2p1_cf_w_0_140_s_3_500=3.95e-11
+  mcm5m2p1_ca_w_1_120_s_0_140=4.89e-05 mcm5m2p1_cc_w_1_120_s_0_140=1.44e-10 mcm5m2p1_cf_w_1_120_s_0_140=2.75e-12
+  mcm5m2p1_ca_w_1_120_s_0_175=4.89e-05 mcm5m2p1_cc_w_1_120_s_0_175=1.38e-10 mcm5m2p1_cf_w_1_120_s_0_175=3.61e-12
+  mcm5m2p1_ca_w_1_120_s_0_210=4.89e-05 mcm5m2p1_cc_w_1_120_s_0_210=1.29e-10 mcm5m2p1_cf_w_1_120_s_0_210=4.46e-12
+  mcm5m2p1_ca_w_1_120_s_0_280=4.89e-05 mcm5m2p1_cc_w_1_120_s_0_280=1.10e-10 mcm5m2p1_cf_w_1_120_s_0_280=6.12e-12
+  mcm5m2p1_ca_w_1_120_s_0_350=4.89e-05 mcm5m2p1_cc_w_1_120_s_0_350=9.31e-11 mcm5m2p1_cf_w_1_120_s_0_350=7.77e-12
+  mcm5m2p1_ca_w_1_120_s_0_420=4.89e-05 mcm5m2p1_cc_w_1_120_s_0_420=7.99e-11 mcm5m2p1_cf_w_1_120_s_0_420=9.36e-12
+  mcm5m2p1_ca_w_1_120_s_0_560=4.89e-05 mcm5m2p1_cc_w_1_120_s_0_560=6.13e-11 mcm5m2p1_cf_w_1_120_s_0_560=1.24e-11
+  mcm5m2p1_ca_w_1_120_s_0_840=4.89e-05 mcm5m2p1_cc_w_1_120_s_0_840=4.10e-11 mcm5m2p1_cf_w_1_120_s_0_840=1.81e-11
+  mcm5m2p1_ca_w_1_120_s_1_540=4.89e-05 mcm5m2p1_cc_w_1_120_s_1_540=1.95e-11 mcm5m2p1_cf_w_1_120_s_1_540=2.89e-11
+  mcm5m2p1_ca_w_1_120_s_3_500=4.89e-05 mcm5m2p1_cc_w_1_120_s_3_500=3.59e-12 mcm5m2p1_cf_w_1_120_s_3_500=4.17e-11
+  mcm5m2l1_ca_w_0_140_s_0_140=6.56e-05 mcm5m2l1_cc_w_0_140_s_0_140=1.25e-10 mcm5m2l1_cf_w_0_140_s_0_140=3.52e-12
+  mcm5m2l1_ca_w_0_140_s_0_175=6.56e-05 mcm5m2l1_cc_w_0_140_s_0_175=1.20e-10 mcm5m2l1_cf_w_0_140_s_0_175=4.65e-12
+  mcm5m2l1_ca_w_0_140_s_0_210=6.56e-05 mcm5m2l1_cc_w_0_140_s_0_210=1.12e-10 mcm5m2l1_cf_w_0_140_s_0_210=5.79e-12
+  mcm5m2l1_ca_w_0_140_s_0_280=6.56e-05 mcm5m2l1_cc_w_0_140_s_0_280=9.48e-11 mcm5m2l1_cf_w_0_140_s_0_280=7.99e-12
+  mcm5m2l1_ca_w_0_140_s_0_350=6.56e-05 mcm5m2l1_cc_w_0_140_s_0_350=7.91e-11 mcm5m2l1_cf_w_0_140_s_0_350=1.01e-11
+  mcm5m2l1_ca_w_0_140_s_0_420=6.56e-05 mcm5m2l1_cc_w_0_140_s_0_420=6.75e-11 mcm5m2l1_cf_w_0_140_s_0_420=1.23e-11
+  mcm5m2l1_ca_w_0_140_s_0_560=6.56e-05 mcm5m2l1_cc_w_0_140_s_0_560=5.06e-11 mcm5m2l1_cf_w_0_140_s_0_560=1.62e-11
+  mcm5m2l1_ca_w_0_140_s_0_840=6.56e-05 mcm5m2l1_cc_w_0_140_s_0_840=3.24e-11 mcm5m2l1_cf_w_0_140_s_0_840=2.31e-11
+  mcm5m2l1_ca_w_0_140_s_1_540=6.56e-05 mcm5m2l1_cc_w_0_140_s_1_540=1.37e-11 mcm5m2l1_cf_w_0_140_s_1_540=3.46e-11
+  mcm5m2l1_ca_w_0_140_s_3_500=6.56e-05 mcm5m2l1_cc_w_0_140_s_3_500=1.98e-12 mcm5m2l1_cf_w_0_140_s_3_500=4.49e-11
+  mcm5m2l1_ca_w_1_120_s_0_140=6.56e-05 mcm5m2l1_cc_w_1_120_s_0_140=1.40e-10 mcm5m2l1_cf_w_1_120_s_0_140=3.57e-12
+  mcm5m2l1_ca_w_1_120_s_0_175=6.56e-05 mcm5m2l1_cc_w_1_120_s_0_175=1.34e-10 mcm5m2l1_cf_w_1_120_s_0_175=4.70e-12
+  mcm5m2l1_ca_w_1_120_s_0_210=6.56e-05 mcm5m2l1_cc_w_1_120_s_0_210=1.25e-10 mcm5m2l1_cf_w_1_120_s_0_210=5.83e-12
+  mcm5m2l1_ca_w_1_120_s_0_280=6.56e-05 mcm5m2l1_cc_w_1_120_s_0_280=1.05e-10 mcm5m2l1_cf_w_1_120_s_0_280=8.04e-12
+  mcm5m2l1_ca_w_1_120_s_0_350=6.56e-05 mcm5m2l1_cc_w_1_120_s_0_350=8.89e-11 mcm5m2l1_cf_w_1_120_s_0_350=1.02e-11
+  mcm5m2l1_ca_w_1_120_s_0_420=6.56e-05 mcm5m2l1_cc_w_1_120_s_0_420=7.56e-11 mcm5m2l1_cf_w_1_120_s_0_420=1.23e-11
+  mcm5m2l1_ca_w_1_120_s_0_560=6.56e-05 mcm5m2l1_cc_w_1_120_s_0_560=5.71e-11 mcm5m2l1_cf_w_1_120_s_0_560=1.62e-11
+  mcm5m2l1_ca_w_1_120_s_0_840=6.56e-05 mcm5m2l1_cc_w_1_120_s_0_840=3.71e-11 mcm5m2l1_cf_w_1_120_s_0_840=2.32e-11
+  mcm5m2l1_ca_w_1_120_s_1_540=6.56e-05 mcm5m2l1_cc_w_1_120_s_1_540=1.63e-11 mcm5m2l1_cf_w_1_120_s_1_540=3.53e-11
+  mcm5m2l1_ca_w_1_120_s_3_500=6.56e-05 mcm5m2l1_cc_w_1_120_s_3_500=2.62e-12 mcm5m2l1_cf_w_1_120_s_3_500=4.72e-11
+  mcm5m2m1_ca_w_0_140_s_0_140=3.26e-04 mcm5m2m1_cc_w_0_140_s_0_140=1.09e-10 mcm5m2m1_cf_w_0_140_s_0_140=1.53e-11
+  mcm5m2m1_ca_w_0_140_s_0_175=3.26e-04 mcm5m2m1_cc_w_0_140_s_0_175=1.03e-10 mcm5m2m1_cf_w_0_140_s_0_175=2.09e-11
+  mcm5m2m1_ca_w_0_140_s_0_210=3.26e-04 mcm5m2m1_cc_w_0_140_s_0_210=9.50e-11 mcm5m2m1_cf_w_0_140_s_0_210=2.59e-11
+  mcm5m2m1_ca_w_0_140_s_0_280=3.26e-04 mcm5m2m1_cc_w_0_140_s_0_280=7.74e-11 mcm5m2m1_cf_w_0_140_s_0_280=3.49e-11
+  mcm5m2m1_ca_w_0_140_s_0_350=3.26e-04 mcm5m2m1_cc_w_0_140_s_0_350=6.26e-11 mcm5m2m1_cf_w_0_140_s_0_350=4.24e-11
+  mcm5m2m1_ca_w_0_140_s_0_420=3.26e-04 mcm5m2m1_cc_w_0_140_s_0_420=5.06e-11 mcm5m2m1_cf_w_0_140_s_0_420=4.89e-11
+  mcm5m2m1_ca_w_0_140_s_0_560=3.26e-04 mcm5m2m1_cc_w_0_140_s_0_560=3.49e-11 mcm5m2m1_cf_w_0_140_s_0_560=5.87e-11
+  mcm5m2m1_ca_w_0_140_s_0_840=3.26e-04 mcm5m2m1_cc_w_0_140_s_0_840=1.92e-11 mcm5m2m1_cf_w_0_140_s_0_840=7.08e-11
+  mcm5m2m1_ca_w_0_140_s_1_540=3.26e-04 mcm5m2m1_cc_w_0_140_s_1_540=6.18e-12 mcm5m2m1_cf_w_0_140_s_1_540=8.38e-11
+  mcm5m2m1_ca_w_0_140_s_3_500=3.26e-04 mcm5m2m1_cc_w_0_140_s_3_500=6.25e-13 mcm5m2m1_cf_w_0_140_s_3_500=9.02e-11
+  mcm5m2m1_ca_w_1_120_s_0_140=3.26e-04 mcm5m2m1_cc_w_1_120_s_0_140=1.21e-10 mcm5m2m1_cf_w_1_120_s_0_140=1.52e-11
+  mcm5m2m1_ca_w_1_120_s_0_175=3.26e-04 mcm5m2m1_cc_w_1_120_s_0_175=1.14e-10 mcm5m2m1_cf_w_1_120_s_0_175=2.08e-11
+  mcm5m2m1_ca_w_1_120_s_0_210=3.26e-04 mcm5m2m1_cc_w_1_120_s_0_210=1.05e-10 mcm5m2m1_cf_w_1_120_s_0_210=2.59e-11
+  mcm5m2m1_ca_w_1_120_s_0_280=3.26e-04 mcm5m2m1_cc_w_1_120_s_0_280=8.62e-11 mcm5m2m1_cf_w_1_120_s_0_280=3.49e-11
+  mcm5m2m1_ca_w_1_120_s_0_350=3.26e-04 mcm5m2m1_cc_w_1_120_s_0_350=7.04e-11 mcm5m2m1_cf_w_1_120_s_0_350=4.24e-11
+  mcm5m2m1_ca_w_1_120_s_0_420=3.26e-04 mcm5m2m1_cc_w_1_120_s_0_420=5.81e-11 mcm5m2m1_cf_w_1_120_s_0_420=4.87e-11
+  mcm5m2m1_ca_w_1_120_s_0_560=3.26e-04 mcm5m2m1_cc_w_1_120_s_0_560=4.07e-11 mcm5m2m1_cf_w_1_120_s_0_560=5.86e-11
+  mcm5m2m1_ca_w_1_120_s_0_840=3.26e-04 mcm5m2m1_cc_w_1_120_s_0_840=2.38e-11 mcm5m2m1_cf_w_1_120_s_0_840=7.11e-11
+  mcm5m2m1_ca_w_1_120_s_1_540=3.26e-04 mcm5m2m1_cc_w_1_120_s_1_540=8.55e-12 mcm5m2m1_cf_w_1_120_s_1_540=8.52e-11
+  mcm5m2m1_ca_w_1_120_s_3_500=3.26e-04 mcm5m2m1_cc_w_1_120_s_3_500=1.00e-12 mcm5m2m1_cf_w_1_120_s_3_500=9.37e-11
+  mcrdlm2f_ca_w_0_140_s_0_140=2.78e-05 mcrdlm2f_cc_w_0_140_s_0_140=1.32e-10 mcrdlm2f_cf_w_0_140_s_0_140=1.52e-12
+  mcrdlm2f_ca_w_0_140_s_0_175=2.78e-05 mcrdlm2f_cc_w_0_140_s_0_175=1.25e-10 mcrdlm2f_cf_w_0_140_s_0_175=2.00e-12
+  mcrdlm2f_ca_w_0_140_s_0_210=2.78e-05 mcrdlm2f_cc_w_0_140_s_0_210=1.17e-10 mcrdlm2f_cf_w_0_140_s_0_210=2.49e-12
+  mcrdlm2f_ca_w_0_140_s_0_280=2.78e-05 mcrdlm2f_cc_w_0_140_s_0_280=1.00e-10 mcrdlm2f_cf_w_0_140_s_0_280=3.45e-12
+  mcrdlm2f_ca_w_0_140_s_0_350=2.78e-05 mcrdlm2f_cc_w_0_140_s_0_350=8.60e-11 mcrdlm2f_cf_w_0_140_s_0_350=4.39e-12
+  mcrdlm2f_ca_w_0_140_s_0_420=2.78e-05 mcrdlm2f_cc_w_0_140_s_0_420=7.45e-11 mcrdlm2f_cf_w_0_140_s_0_420=5.36e-12
+  mcrdlm2f_ca_w_0_140_s_0_560=2.78e-05 mcrdlm2f_cc_w_0_140_s_0_560=5.92e-11 mcrdlm2f_cf_w_0_140_s_0_560=7.15e-12
+  mcrdlm2f_ca_w_0_140_s_0_840=2.78e-05 mcrdlm2f_cc_w_0_140_s_0_840=4.24e-11 mcrdlm2f_cf_w_0_140_s_0_840=1.06e-11
+  mcrdlm2f_ca_w_0_140_s_1_540=2.78e-05 mcrdlm2f_cc_w_0_140_s_1_540=2.44e-11 mcrdlm2f_cf_w_0_140_s_1_540=1.77e-11
+  mcrdlm2f_ca_w_0_140_s_3_500=2.78e-05 mcrdlm2f_cc_w_0_140_s_3_500=8.34e-12 mcrdlm2f_cf_w_0_140_s_3_500=2.90e-11
+  mcrdlm2f_ca_w_1_120_s_0_140=2.78e-05 mcrdlm2f_cc_w_1_120_s_0_140=1.53e-10 mcrdlm2f_cf_w_1_120_s_0_140=1.56e-12
+  mcrdlm2f_ca_w_1_120_s_0_175=2.78e-05 mcrdlm2f_cc_w_1_120_s_0_175=1.46e-10 mcrdlm2f_cf_w_1_120_s_0_175=2.05e-12
+  mcrdlm2f_ca_w_1_120_s_0_210=2.78e-05 mcrdlm2f_cc_w_1_120_s_0_210=1.38e-10 mcrdlm2f_cf_w_1_120_s_0_210=2.54e-12
+  mcrdlm2f_ca_w_1_120_s_0_280=2.78e-05 mcrdlm2f_cc_w_1_120_s_0_280=1.19e-10 mcrdlm2f_cf_w_1_120_s_0_280=3.48e-12
+  mcrdlm2f_ca_w_1_120_s_0_350=2.78e-05 mcrdlm2f_cc_w_1_120_s_0_350=1.03e-10 mcrdlm2f_cf_w_1_120_s_0_350=4.43e-12
+  mcrdlm2f_ca_w_1_120_s_0_420=2.78e-05 mcrdlm2f_cc_w_1_120_s_0_420=8.97e-11 mcrdlm2f_cf_w_1_120_s_0_420=5.36e-12
+  mcrdlm2f_ca_w_1_120_s_0_560=2.78e-05 mcrdlm2f_cc_w_1_120_s_0_560=7.16e-11 mcrdlm2f_cf_w_1_120_s_0_560=7.19e-12
+  mcrdlm2f_ca_w_1_120_s_0_840=2.78e-05 mcrdlm2f_cc_w_1_120_s_0_840=5.21e-11 mcrdlm2f_cf_w_1_120_s_0_840=1.07e-11
+  mcrdlm2f_ca_w_1_120_s_1_540=2.78e-05 mcrdlm2f_cc_w_1_120_s_1_540=3.07e-11 mcrdlm2f_cf_w_1_120_s_1_540=1.81e-11
+  mcrdlm2f_ca_w_1_120_s_3_500=2.78e-05 mcrdlm2f_cc_w_1_120_s_3_500=1.13e-11 mcrdlm2f_cf_w_1_120_s_3_500=3.08e-11
+  mcrdlm2d_ca_w_0_140_s_0_140=3.17e-05 mcrdlm2d_cc_w_0_140_s_0_140=1.31e-10 mcrdlm2d_cf_w_0_140_s_0_140=1.73e-12
+  mcrdlm2d_ca_w_0_140_s_0_175=3.17e-05 mcrdlm2d_cc_w_0_140_s_0_175=1.24e-10 mcrdlm2d_cf_w_0_140_s_0_175=2.28e-12
+  mcrdlm2d_ca_w_0_140_s_0_210=3.17e-05 mcrdlm2d_cc_w_0_140_s_0_210=1.17e-10 mcrdlm2d_cf_w_0_140_s_0_210=2.83e-12
+  mcrdlm2d_ca_w_0_140_s_0_280=3.17e-05 mcrdlm2d_cc_w_0_140_s_0_280=9.97e-11 mcrdlm2d_cf_w_0_140_s_0_280=3.92e-12
+  mcrdlm2d_ca_w_0_140_s_0_350=3.17e-05 mcrdlm2d_cc_w_0_140_s_0_350=8.53e-11 mcrdlm2d_cf_w_0_140_s_0_350=4.99e-12
+  mcrdlm2d_ca_w_0_140_s_0_420=3.17e-05 mcrdlm2d_cc_w_0_140_s_0_420=7.37e-11 mcrdlm2d_cf_w_0_140_s_0_420=6.08e-12
+  mcrdlm2d_ca_w_0_140_s_0_560=3.17e-05 mcrdlm2d_cc_w_0_140_s_0_560=5.82e-11 mcrdlm2d_cf_w_0_140_s_0_560=8.11e-12
+  mcrdlm2d_ca_w_0_140_s_0_840=3.17e-05 mcrdlm2d_cc_w_0_140_s_0_840=4.12e-11 mcrdlm2d_cf_w_0_140_s_0_840=1.19e-11
+  mcrdlm2d_ca_w_0_140_s_1_540=3.17e-05 mcrdlm2d_cc_w_0_140_s_1_540=2.31e-11 mcrdlm2d_cf_w_0_140_s_1_540=1.97e-11
+  mcrdlm2d_ca_w_0_140_s_3_500=3.17e-05 mcrdlm2d_cc_w_0_140_s_3_500=7.44e-12 mcrdlm2d_cf_w_0_140_s_3_500=3.13e-11
+  mcrdlm2d_ca_w_1_120_s_0_140=3.17e-05 mcrdlm2d_cc_w_1_120_s_0_140=1.51e-10 mcrdlm2d_cf_w_1_120_s_0_140=1.78e-12
+  mcrdlm2d_ca_w_1_120_s_0_175=3.17e-05 mcrdlm2d_cc_w_1_120_s_0_175=1.45e-10 mcrdlm2d_cf_w_1_120_s_0_175=2.33e-12
+  mcrdlm2d_ca_w_1_120_s_0_210=3.17e-05 mcrdlm2d_cc_w_1_120_s_0_210=1.37e-10 mcrdlm2d_cf_w_1_120_s_0_210=2.88e-12
+  mcrdlm2d_ca_w_1_120_s_0_280=3.17e-05 mcrdlm2d_cc_w_1_120_s_0_280=1.18e-10 mcrdlm2d_cf_w_1_120_s_0_280=3.97e-12
+  mcrdlm2d_ca_w_1_120_s_0_350=3.17e-05 mcrdlm2d_cc_w_1_120_s_0_350=1.01e-10 mcrdlm2d_cf_w_1_120_s_0_350=5.04e-12
+  mcrdlm2d_ca_w_1_120_s_0_420=3.17e-05 mcrdlm2d_cc_w_1_120_s_0_420=8.81e-11 mcrdlm2d_cf_w_1_120_s_0_420=6.10e-12
+  mcrdlm2d_ca_w_1_120_s_0_560=3.17e-05 mcrdlm2d_cc_w_1_120_s_0_560=7.00e-11 mcrdlm2d_cf_w_1_120_s_0_560=8.16e-12
+  mcrdlm2d_ca_w_1_120_s_0_840=3.17e-05 mcrdlm2d_cc_w_1_120_s_0_840=5.04e-11 mcrdlm2d_cf_w_1_120_s_0_840=1.20e-11
+  mcrdlm2d_ca_w_1_120_s_1_540=3.17e-05 mcrdlm2d_cc_w_1_120_s_1_540=2.91e-11 mcrdlm2d_cf_w_1_120_s_1_540=2.01e-11
+  mcrdlm2d_ca_w_1_120_s_3_500=3.17e-05 mcrdlm2d_cc_w_1_120_s_3_500=1.01e-11 mcrdlm2d_cf_w_1_120_s_3_500=3.31e-11
+  mcrdlm2p1_ca_w_0_140_s_0_140=3.98e-05 mcrdlm2p1_cc_w_0_140_s_0_140=1.30e-10 mcrdlm2p1_cf_w_0_140_s_0_140=2.17e-12
+  mcrdlm2p1_ca_w_0_140_s_0_175=3.98e-05 mcrdlm2p1_cc_w_0_140_s_0_175=1.23e-10 mcrdlm2p1_cf_w_0_140_s_0_175=2.87e-12
+  mcrdlm2p1_ca_w_0_140_s_0_210=3.98e-05 mcrdlm2p1_cc_w_0_140_s_0_210=1.15e-10 mcrdlm2p1_cf_w_0_140_s_0_210=3.56e-12
+  mcrdlm2p1_ca_w_0_140_s_0_280=3.98e-05 mcrdlm2p1_cc_w_0_140_s_0_280=9.84e-11 mcrdlm2p1_cf_w_0_140_s_0_280=4.92e-12
+  mcrdlm2p1_ca_w_0_140_s_0_350=3.98e-05 mcrdlm2p1_cc_w_0_140_s_0_350=8.35e-11 mcrdlm2p1_cf_w_0_140_s_0_350=6.26e-12
+  mcrdlm2p1_ca_w_0_140_s_0_420=3.98e-05 mcrdlm2p1_cc_w_0_140_s_0_420=7.21e-11 mcrdlm2p1_cf_w_0_140_s_0_420=7.60e-12
+  mcrdlm2p1_ca_w_0_140_s_0_560=3.98e-05 mcrdlm2p1_cc_w_0_140_s_0_560=5.61e-11 mcrdlm2p1_cf_w_0_140_s_0_560=1.01e-11
+  mcrdlm2p1_ca_w_0_140_s_0_840=3.98e-05 mcrdlm2p1_cc_w_0_140_s_0_840=3.91e-11 mcrdlm2p1_cf_w_0_140_s_0_840=1.47e-11
+  mcrdlm2p1_ca_w_0_140_s_1_540=3.98e-05 mcrdlm2p1_cc_w_0_140_s_1_540=2.08e-11 mcrdlm2p1_cf_w_0_140_s_1_540=2.37e-11
+  mcrdlm2p1_ca_w_0_140_s_3_500=3.98e-05 mcrdlm2p1_cc_w_0_140_s_3_500=6.03e-12 mcrdlm2p1_cf_w_0_140_s_3_500=3.52e-11
+  mcrdlm2p1_ca_w_1_120_s_0_140=3.98e-05 mcrdlm2p1_cc_w_1_120_s_0_140=1.49e-10 mcrdlm2p1_cf_w_1_120_s_0_140=2.28e-12
+  mcrdlm2p1_ca_w_1_120_s_0_175=3.98e-05 mcrdlm2p1_cc_w_1_120_s_0_175=1.42e-10 mcrdlm2p1_cf_w_1_120_s_0_175=2.98e-12
+  mcrdlm2p1_ca_w_1_120_s_0_210=3.98e-05 mcrdlm2p1_cc_w_1_120_s_0_210=1.34e-10 mcrdlm2p1_cf_w_1_120_s_0_210=3.67e-12
+  mcrdlm2p1_ca_w_1_120_s_0_280=3.98e-05 mcrdlm2p1_cc_w_1_120_s_0_280=1.15e-10 mcrdlm2p1_cf_w_1_120_s_0_280=5.00e-12
+  mcrdlm2p1_ca_w_1_120_s_0_350=3.98e-05 mcrdlm2p1_cc_w_1_120_s_0_350=9.80e-11 mcrdlm2p1_cf_w_1_120_s_0_350=6.34e-12
+  mcrdlm2p1_ca_w_1_120_s_0_420=3.98e-05 mcrdlm2p1_cc_w_1_120_s_0_420=8.50e-11 mcrdlm2p1_cf_w_1_120_s_0_420=7.65e-12
+  mcrdlm2p1_ca_w_1_120_s_0_560=3.98e-05 mcrdlm2p1_cc_w_1_120_s_0_560=6.72e-11 mcrdlm2p1_cf_w_1_120_s_0_560=1.02e-11
+  mcrdlm2p1_ca_w_1_120_s_0_840=3.98e-05 mcrdlm2p1_cc_w_1_120_s_0_840=4.74e-11 mcrdlm2p1_cf_w_1_120_s_0_840=1.48e-11
+  mcrdlm2p1_ca_w_1_120_s_1_540=3.98e-05 mcrdlm2p1_cc_w_1_120_s_1_540=2.64e-11 mcrdlm2p1_cf_w_1_120_s_1_540=2.41e-11
+  mcrdlm2p1_ca_w_1_120_s_3_500=3.98e-05 mcrdlm2p1_cc_w_1_120_s_3_500=8.63e-12 mcrdlm2p1_cf_w_1_120_s_3_500=3.74e-11
+  mcrdlm2l1_ca_w_0_140_s_0_140=5.66e-05 mcrdlm2l1_cc_w_0_140_s_0_140=1.26e-10 mcrdlm2l1_cf_w_0_140_s_0_140=3.03e-12
+  mcrdlm2l1_ca_w_0_140_s_0_175=5.66e-05 mcrdlm2l1_cc_w_0_140_s_0_175=1.21e-10 mcrdlm2l1_cf_w_0_140_s_0_175=4.01e-12
+  mcrdlm2l1_ca_w_0_140_s_0_210=5.66e-05 mcrdlm2l1_cc_w_0_140_s_0_210=1.13e-10 mcrdlm2l1_cf_w_0_140_s_0_210=4.99e-12
+  mcrdlm2l1_ca_w_0_140_s_0_280=5.66e-05 mcrdlm2l1_cc_w_0_140_s_0_280=9.63e-11 mcrdlm2l1_cf_w_0_140_s_0_280=6.90e-12
+  mcrdlm2l1_ca_w_0_140_s_0_350=5.66e-05 mcrdlm2l1_cc_w_0_140_s_0_350=8.08e-11 mcrdlm2l1_cf_w_0_140_s_0_350=8.74e-12
+  mcrdlm2l1_ca_w_0_140_s_0_420=5.66e-05 mcrdlm2l1_cc_w_0_140_s_0_420=6.93e-11 mcrdlm2l1_cf_w_0_140_s_0_420=1.06e-11
+  mcrdlm2l1_ca_w_0_140_s_0_560=5.66e-05 mcrdlm2l1_cc_w_0_140_s_0_560=5.28e-11 mcrdlm2l1_cf_w_0_140_s_0_560=1.39e-11
+  mcrdlm2l1_ca_w_0_140_s_0_840=5.66e-05 mcrdlm2l1_cc_w_0_140_s_0_840=3.55e-11 mcrdlm2l1_cf_w_0_140_s_0_840=1.98e-11
+  mcrdlm2l1_ca_w_0_140_s_1_540=5.66e-05 mcrdlm2l1_cc_w_0_140_s_1_540=1.76e-11 mcrdlm2l1_cf_w_0_140_s_1_540=3.04e-11
+  mcrdlm2l1_ca_w_0_140_s_3_500=5.66e-05 mcrdlm2l1_cc_w_0_140_s_3_500=4.50e-12 mcrdlm2l1_cf_w_0_140_s_3_500=4.16e-11
+  mcrdlm2l1_ca_w_1_120_s_0_140=5.66e-05 mcrdlm2l1_cc_w_1_120_s_0_140=1.45e-10 mcrdlm2l1_cf_w_1_120_s_0_140=3.08e-12
+  mcrdlm2l1_ca_w_1_120_s_0_175=5.66e-05 mcrdlm2l1_cc_w_1_120_s_0_175=1.38e-10 mcrdlm2l1_cf_w_1_120_s_0_175=4.07e-12
+  mcrdlm2l1_ca_w_1_120_s_0_210=5.66e-05 mcrdlm2l1_cc_w_1_120_s_0_210=1.30e-10 mcrdlm2l1_cf_w_1_120_s_0_210=5.05e-12
+  mcrdlm2l1_ca_w_1_120_s_0_280=5.66e-05 mcrdlm2l1_cc_w_1_120_s_0_280=1.10e-10 mcrdlm2l1_cf_w_1_120_s_0_280=6.94e-12
+  mcrdlm2l1_ca_w_1_120_s_0_350=5.66e-05 mcrdlm2l1_cc_w_1_120_s_0_350=9.39e-11 mcrdlm2l1_cf_w_1_120_s_0_350=8.78e-12
+  mcrdlm2l1_ca_w_1_120_s_0_420=5.66e-05 mcrdlm2l1_cc_w_1_120_s_0_420=8.12e-11 mcrdlm2l1_cf_w_1_120_s_0_420=1.06e-11
+  mcrdlm2l1_ca_w_1_120_s_0_560=5.66e-05 mcrdlm2l1_cc_w_1_120_s_0_560=6.30e-11 mcrdlm2l1_cf_w_1_120_s_0_560=1.40e-11
+  mcrdlm2l1_ca_w_1_120_s_0_840=5.66e-05 mcrdlm2l1_cc_w_1_120_s_0_840=4.34e-11 mcrdlm2l1_cf_w_1_120_s_0_840=2.00e-11
+  mcrdlm2l1_ca_w_1_120_s_1_540=5.66e-05 mcrdlm2l1_cc_w_1_120_s_1_540=2.29e-11 mcrdlm2l1_cf_w_1_120_s_1_540=3.10e-11
+  mcrdlm2l1_ca_w_1_120_s_3_500=5.66e-05 mcrdlm2l1_cc_w_1_120_s_3_500=6.86e-12 mcrdlm2l1_cf_w_1_120_s_3_500=4.41e-11
+  mcrdlm2m1_ca_w_0_140_s_0_140=3.17e-04 mcrdlm2m1_cc_w_0_140_s_0_140=1.10e-10 mcrdlm2m1_cf_w_0_140_s_0_140=1.48e-11
+  mcrdlm2m1_ca_w_0_140_s_0_175=3.17e-04 mcrdlm2m1_cc_w_0_140_s_0_175=1.04e-10 mcrdlm2m1_cf_w_0_140_s_0_175=2.02e-11
+  mcrdlm2m1_ca_w_0_140_s_0_210=3.17e-04 mcrdlm2m1_cc_w_0_140_s_0_210=9.63e-11 mcrdlm2m1_cf_w_0_140_s_0_210=2.51e-11
+  mcrdlm2m1_ca_w_0_140_s_0_280=3.17e-04 mcrdlm2m1_cc_w_0_140_s_0_280=7.89e-11 mcrdlm2m1_cf_w_0_140_s_0_280=3.38e-11
+  mcrdlm2m1_ca_w_0_140_s_0_350=3.17e-04 mcrdlm2m1_cc_w_0_140_s_0_350=6.41e-11 mcrdlm2m1_cf_w_0_140_s_0_350=4.10e-11
+  mcrdlm2m1_ca_w_0_140_s_0_420=3.17e-04 mcrdlm2m1_cc_w_0_140_s_0_420=5.25e-11 mcrdlm2m1_cf_w_0_140_s_0_420=4.71e-11
+  mcrdlm2m1_ca_w_0_140_s_0_560=3.17e-04 mcrdlm2m1_cc_w_0_140_s_0_560=3.71e-11 mcrdlm2m1_cf_w_0_140_s_0_560=5.64e-11
+  mcrdlm2m1_ca_w_0_140_s_0_840=3.17e-04 mcrdlm2m1_cc_w_0_140_s_0_840=2.20e-11 mcrdlm2m1_cf_w_0_140_s_0_840=6.82e-11
+  mcrdlm2m1_ca_w_0_140_s_1_540=3.17e-04 mcrdlm2m1_cc_w_0_140_s_1_540=8.59e-12 mcrdlm2m1_cf_w_0_140_s_1_540=8.12e-11
+  mcrdlm2m1_ca_w_0_140_s_3_500=3.17e-04 mcrdlm2m1_cc_w_0_140_s_3_500=1.76e-12 mcrdlm2m1_cf_w_0_140_s_3_500=8.90e-11
+  mcrdlm2m1_ca_w_1_120_s_0_140=3.17e-04 mcrdlm2m1_cc_w_1_120_s_0_140=1.27e-10 mcrdlm2m1_cf_w_1_120_s_0_140=1.47e-11
+  mcrdlm2m1_ca_w_1_120_s_0_175=3.17e-04 mcrdlm2m1_cc_w_1_120_s_0_175=1.19e-10 mcrdlm2m1_cf_w_1_120_s_0_175=2.02e-11
+  mcrdlm2m1_ca_w_1_120_s_0_210=3.17e-04 mcrdlm2m1_cc_w_1_120_s_0_210=1.10e-10 mcrdlm2m1_cf_w_1_120_s_0_210=2.52e-11
+  mcrdlm2m1_ca_w_1_120_s_0_280=3.17e-04 mcrdlm2m1_cc_w_1_120_s_0_280=9.08e-11 mcrdlm2m1_cf_w_1_120_s_0_280=3.38e-11
+  mcrdlm2m1_ca_w_1_120_s_0_350=3.17e-04 mcrdlm2m1_cc_w_1_120_s_0_350=7.54e-11 mcrdlm2m1_cf_w_1_120_s_0_350=4.11e-11
+  mcrdlm2m1_ca_w_1_120_s_0_420=3.17e-04 mcrdlm2m1_cc_w_1_120_s_0_420=6.32e-11 mcrdlm2m1_cf_w_1_120_s_0_420=4.70e-11
+  mcrdlm2m1_ca_w_1_120_s_0_560=3.17e-04 mcrdlm2m1_cc_w_1_120_s_0_560=4.65e-11 mcrdlm2m1_cf_w_1_120_s_0_560=5.63e-11
+  mcrdlm2m1_ca_w_1_120_s_0_840=3.17e-04 mcrdlm2m1_cc_w_1_120_s_0_840=2.96e-11 mcrdlm2m1_cf_w_1_120_s_0_840=6.85e-11
+  mcrdlm2m1_ca_w_1_120_s_1_540=3.17e-04 mcrdlm2m1_cc_w_1_120_s_1_540=1.38e-11 mcrdlm2m1_cf_w_1_120_s_1_540=8.28e-11
+  mcrdlm2m1_ca_w_1_120_s_3_500=3.17e-04 mcrdlm2m1_cc_w_1_120_s_3_500=3.56e-12 mcrdlm2m1_cf_w_1_120_s_3_500=9.36e-11
+  mcm4m3f_ca_w_0_300_s_0_300=2.08e-04 mcm4m3f_cc_w_0_300_s_0_300=1.00e-10 mcm4m3f_cf_w_0_300_s_0_300=1.90e-11
+  mcm4m3f_ca_w_0_300_s_0_360=2.08e-04 mcm4m3f_cc_w_0_300_s_0_360=9.01e-11 mcm4m3f_cf_w_0_300_s_0_360=2.26e-11
+  mcm4m3f_ca_w_0_300_s_0_450=2.08e-04 mcm4m3f_cc_w_0_300_s_0_450=7.72e-11 mcm4m3f_cf_w_0_300_s_0_450=2.75e-11
+  mcm4m3f_ca_w_0_300_s_0_600=2.08e-04 mcm4m3f_cc_w_0_300_s_0_600=6.06e-11 mcm4m3f_cf_w_0_300_s_0_600=3.45e-11
+  mcm4m3f_ca_w_0_300_s_0_800=2.08e-04 mcm4m3f_cc_w_0_300_s_0_800=4.48e-11 mcm4m3f_cf_w_0_300_s_0_800=4.19e-11
+  mcm4m3f_ca_w_0_300_s_1_000=2.08e-04 mcm4m3f_cc_w_0_300_s_1_000=3.37e-11 mcm4m3f_cf_w_0_300_s_1_000=4.81e-11
+  mcm4m3f_ca_w_0_300_s_1_200=2.08e-04 mcm4m3f_cc_w_0_300_s_1_200=2.57e-11 mcm4m3f_cf_w_0_300_s_1_200=5.27e-11
+  mcm4m3f_ca_w_0_300_s_2_100=2.08e-04 mcm4m3f_cc_w_0_300_s_2_100=8.98e-12 mcm4m3f_cf_w_0_300_s_2_100=6.53e-11
+  mcm4m3f_ca_w_0_300_s_3_300=2.08e-04 mcm4m3f_cc_w_0_300_s_3_300=2.57e-12 mcm4m3f_cf_w_0_300_s_3_300=7.13e-11
+  mcm4m3f_ca_w_0_300_s_9_000=2.08e-04 mcm4m3f_cc_w_0_300_s_9_000=3.50e-14 mcm4m3f_cf_w_0_300_s_9_000=7.39e-11
+  mcm4m3f_ca_w_2_400_s_0_300=2.08e-04 mcm4m3f_cc_w_2_400_s_0_300=1.07e-10 mcm4m3f_cf_w_2_400_s_0_300=1.90e-11
+  mcm4m3f_ca_w_2_400_s_0_360=2.08e-04 mcm4m3f_cc_w_2_400_s_0_360=9.54e-11 mcm4m3f_cf_w_2_400_s_0_360=2.26e-11
+  mcm4m3f_ca_w_2_400_s_0_450=2.08e-04 mcm4m3f_cc_w_2_400_s_0_450=8.19e-11 mcm4m3f_cf_w_2_400_s_0_450=2.75e-11
+  mcm4m3f_ca_w_2_400_s_0_600=2.08e-04 mcm4m3f_cc_w_2_400_s_0_600=6.47e-11 mcm4m3f_cf_w_2_400_s_0_600=3.44e-11
+  mcm4m3f_ca_w_2_400_s_0_800=2.08e-04 mcm4m3f_cc_w_2_400_s_0_800=4.80e-11 mcm4m3f_cf_w_2_400_s_0_800=4.19e-11
+  mcm4m3f_ca_w_2_400_s_1_000=2.08e-04 mcm4m3f_cc_w_2_400_s_1_000=3.63e-11 mcm4m3f_cf_w_2_400_s_1_000=4.81e-11
+  mcm4m3f_ca_w_2_400_s_1_200=2.08e-04 mcm4m3f_cc_w_2_400_s_1_200=2.79e-11 mcm4m3f_cf_w_2_400_s_1_200=5.29e-11
+  mcm4m3f_ca_w_2_400_s_2_100=2.08e-04 mcm4m3f_cc_w_2_400_s_2_100=1.01e-11 mcm4m3f_cf_w_2_400_s_2_100=6.61e-11
+  mcm4m3f_ca_w_2_400_s_3_300=2.08e-04 mcm4m3f_cc_w_2_400_s_3_300=3.01e-12 mcm4m3f_cf_w_2_400_s_3_300=7.25e-11
+  mcm4m3f_ca_w_2_400_s_9_000=2.08e-04 mcm4m3f_cc_w_2_400_s_9_000=1.50e-14 mcm4m3f_cf_w_2_400_s_9_000=7.55e-11
+  mcm4m3d_ca_w_0_300_s_0_300=2.09e-04 mcm4m3d_cc_w_0_300_s_0_300=9.97e-11 mcm4m3d_cf_w_0_300_s_0_300=1.92e-11
+  mcm4m3d_ca_w_0_300_s_0_360=2.09e-04 mcm4m3d_cc_w_0_300_s_0_360=8.96e-11 mcm4m3d_cf_w_0_300_s_0_360=2.29e-11
+  mcm4m3d_ca_w_0_300_s_0_450=2.09e-04 mcm4m3d_cc_w_0_300_s_0_450=7.68e-11 mcm4m3d_cf_w_0_300_s_0_450=2.78e-11
+  mcm4m3d_ca_w_0_300_s_0_600=2.09e-04 mcm4m3d_cc_w_0_300_s_0_600=5.99e-11 mcm4m3d_cf_w_0_300_s_0_600=3.49e-11
+  mcm4m3d_ca_w_0_300_s_0_800=2.09e-04 mcm4m3d_cc_w_0_300_s_0_800=4.41e-11 mcm4m3d_cf_w_0_300_s_0_800=4.25e-11
+  mcm4m3d_ca_w_0_300_s_1_000=2.09e-04 mcm4m3d_cc_w_0_300_s_1_000=3.30e-11 mcm4m3d_cf_w_0_300_s_1_000=4.86e-11
+  mcm4m3d_ca_w_0_300_s_1_200=2.09e-04 mcm4m3d_cc_w_0_300_s_1_200=2.51e-11 mcm4m3d_cf_w_0_300_s_1_200=5.35e-11
+  mcm4m3d_ca_w_0_300_s_2_100=2.09e-04 mcm4m3d_cc_w_0_300_s_2_100=8.34e-12 mcm4m3d_cf_w_0_300_s_2_100=6.61e-11
+  mcm4m3d_ca_w_0_300_s_3_300=2.09e-04 mcm4m3d_cc_w_0_300_s_3_300=2.30e-12 mcm4m3d_cf_w_0_300_s_3_300=7.19e-11
+  mcm4m3d_ca_w_0_300_s_9_000=2.09e-04 mcm4m3d_cc_w_0_300_s_9_000=6.00e-14 mcm4m3d_cf_w_0_300_s_9_000=7.42e-11
+  mcm4m3d_ca_w_2_400_s_0_300=2.09e-04 mcm4m3d_cc_w_2_400_s_0_300=1.06e-10 mcm4m3d_cf_w_2_400_s_0_300=1.93e-11
+  mcm4m3d_ca_w_2_400_s_0_360=2.09e-04 mcm4m3d_cc_w_2_400_s_0_360=9.43e-11 mcm4m3d_cf_w_2_400_s_0_360=2.29e-11
+  mcm4m3d_ca_w_2_400_s_0_450=2.09e-04 mcm4m3d_cc_w_2_400_s_0_450=8.09e-11 mcm4m3d_cf_w_2_400_s_0_450=2.78e-11
+  mcm4m3d_ca_w_2_400_s_0_600=2.09e-04 mcm4m3d_cc_w_2_400_s_0_600=6.36e-11 mcm4m3d_cf_w_2_400_s_0_600=3.48e-11
+  mcm4m3d_ca_w_2_400_s_0_800=2.09e-04 mcm4m3d_cc_w_2_400_s_0_800=4.69e-11 mcm4m3d_cf_w_2_400_s_0_800=4.25e-11
+  mcm4m3d_ca_w_2_400_s_1_000=2.09e-04 mcm4m3d_cc_w_2_400_s_1_000=3.52e-11 mcm4m3d_cf_w_2_400_s_1_000=4.88e-11
+  mcm4m3d_ca_w_2_400_s_1_200=2.09e-04 mcm4m3d_cc_w_2_400_s_1_200=2.69e-11 mcm4m3d_cf_w_2_400_s_1_200=5.37e-11
+  mcm4m3d_ca_w_2_400_s_2_100=2.09e-04 mcm4m3d_cc_w_2_400_s_2_100=9.28e-12 mcm4m3d_cf_w_2_400_s_2_100=6.69e-11
+  mcm4m3d_ca_w_2_400_s_3_300=2.09e-04 mcm4m3d_cc_w_2_400_s_3_300=2.58e-12 mcm4m3d_cf_w_2_400_s_3_300=7.30e-11
+  mcm4m3d_ca_w_2_400_s_9_000=2.09e-04 mcm4m3d_cc_w_2_400_s_9_000=7.00e-14 mcm4m3d_cf_w_2_400_s_9_000=7.56e-11
+  mcm4m3p1_ca_w_0_300_s_0_300=2.13e-04 mcm4m3p1_cc_w_0_300_s_0_300=9.89e-11 mcm4m3p1_cf_w_0_300_s_0_300=1.96e-11
+  mcm4m3p1_ca_w_0_300_s_0_360=2.13e-04 mcm4m3p1_cc_w_0_300_s_0_360=8.87e-11 mcm4m3p1_cf_w_0_300_s_0_360=2.34e-11
+  mcm4m3p1_ca_w_0_300_s_0_450=2.13e-04 mcm4m3p1_cc_w_0_300_s_0_450=7.58e-11 mcm4m3p1_cf_w_0_300_s_0_450=2.84e-11
+  mcm4m3p1_ca_w_0_300_s_0_600=2.13e-04 mcm4m3p1_cc_w_0_300_s_0_600=5.89e-11 mcm4m3p1_cf_w_0_300_s_0_600=3.57e-11
+  mcm4m3p1_ca_w_0_300_s_0_800=2.13e-04 mcm4m3p1_cc_w_0_300_s_0_800=4.30e-11 mcm4m3p1_cf_w_0_300_s_0_800=4.35e-11
+  mcm4m3p1_ca_w_0_300_s_1_000=2.13e-04 mcm4m3p1_cc_w_0_300_s_1_000=3.19e-11 mcm4m3p1_cf_w_0_300_s_1_000=4.99e-11
+  mcm4m3p1_ca_w_0_300_s_1_200=2.13e-04 mcm4m3p1_cc_w_0_300_s_1_200=2.38e-11 mcm4m3p1_cf_w_0_300_s_1_200=5.48e-11
+  mcm4m3p1_ca_w_0_300_s_2_100=2.13e-04 mcm4m3p1_cc_w_0_300_s_2_100=7.46e-12 mcm4m3p1_cf_w_0_300_s_2_100=6.75e-11
+  mcm4m3p1_ca_w_0_300_s_3_300=2.13e-04 mcm4m3p1_cc_w_0_300_s_3_300=1.83e-12 mcm4m3p1_cf_w_0_300_s_3_300=7.28e-11
+  mcm4m3p1_ca_w_0_300_s_9_000=2.13e-04 mcm4m3p1_cc_w_0_300_s_9_000=2.00e-14 mcm4m3p1_cf_w_0_300_s_9_000=7.47e-11
+  mcm4m3p1_ca_w_2_400_s_0_300=2.13e-04 mcm4m3p1_cc_w_2_400_s_0_300=1.03e-10 mcm4m3p1_cf_w_2_400_s_0_300=1.97e-11
+  mcm4m3p1_ca_w_2_400_s_0_360=2.13e-04 mcm4m3p1_cc_w_2_400_s_0_360=9.25e-11 mcm4m3p1_cf_w_2_400_s_0_360=2.34e-11
+  mcm4m3p1_ca_w_2_400_s_0_450=2.13e-04 mcm4m3p1_cc_w_2_400_s_0_450=7.92e-11 mcm4m3p1_cf_w_2_400_s_0_450=2.84e-11
+  mcm4m3p1_ca_w_2_400_s_0_600=2.13e-04 mcm4m3p1_cc_w_2_400_s_0_600=6.17e-11 mcm4m3p1_cf_w_2_400_s_0_600=3.57e-11
+  mcm4m3p1_ca_w_2_400_s_0_800=2.13e-04 mcm4m3p1_cc_w_2_400_s_0_800=4.52e-11 mcm4m3p1_cf_w_2_400_s_0_800=4.36e-11
+  mcm4m3p1_ca_w_2_400_s_1_000=2.13e-04 mcm4m3p1_cc_w_2_400_s_1_000=3.35e-11 mcm4m3p1_cf_w_2_400_s_1_000=5.00e-11
+  mcm4m3p1_ca_w_2_400_s_1_200=2.13e-04 mcm4m3p1_cc_w_2_400_s_1_200=2.52e-11 mcm4m3p1_cf_w_2_400_s_1_200=5.50e-11
+  mcm4m3p1_ca_w_2_400_s_2_100=2.13e-04 mcm4m3p1_cc_w_2_400_s_2_100=8.05e-12 mcm4m3p1_cf_w_2_400_s_2_100=6.82e-11
+  mcm4m3p1_ca_w_2_400_s_3_300=2.13e-04 mcm4m3p1_cc_w_2_400_s_3_300=2.03e-12 mcm4m3p1_cf_w_2_400_s_3_300=7.38e-11
+  mcm4m3p1_ca_w_2_400_s_9_000=2.13e-04 mcm4m3p1_cc_w_2_400_s_9_000=5.50e-14 mcm4m3p1_cf_w_2_400_s_9_000=7.59e-11
+  mcm4m3l1_ca_w_0_300_s_0_300=2.18e-04 mcm4m3l1_cc_w_0_300_s_0_300=9.77e-11 mcm4m3l1_cf_w_0_300_s_0_300=2.02e-11
+  mcm4m3l1_ca_w_0_300_s_0_360=2.18e-04 mcm4m3l1_cc_w_0_300_s_0_360=8.74e-11 mcm4m3l1_cf_w_0_300_s_0_360=2.41e-11
+  mcm4m3l1_ca_w_0_300_s_0_450=2.18e-04 mcm4m3l1_cc_w_0_300_s_0_450=7.45e-11 mcm4m3l1_cf_w_0_300_s_0_450=2.93e-11
+  mcm4m3l1_ca_w_0_300_s_0_600=2.18e-04 mcm4m3l1_cc_w_0_300_s_0_600=5.75e-11 mcm4m3l1_cf_w_0_300_s_0_600=3.69e-11
+  mcm4m3l1_ca_w_0_300_s_0_800=2.18e-04 mcm4m3l1_cc_w_0_300_s_0_800=4.14e-11 mcm4m3l1_cf_w_0_300_s_0_800=4.51e-11
+  mcm4m3l1_ca_w_0_300_s_1_000=2.18e-04 mcm4m3l1_cc_w_0_300_s_1_000=3.01e-11 mcm4m3l1_cf_w_0_300_s_1_000=5.16e-11
+  mcm4m3l1_ca_w_0_300_s_1_200=2.18e-04 mcm4m3l1_cc_w_0_300_s_1_200=2.23e-11 mcm4m3l1_cf_w_0_300_s_1_200=5.68e-11
+  mcm4m3l1_ca_w_0_300_s_2_100=2.18e-04 mcm4m3l1_cc_w_0_300_s_2_100=6.32e-12 mcm4m3l1_cf_w_0_300_s_2_100=6.94e-11
+  mcm4m3l1_ca_w_0_300_s_3_300=2.18e-04 mcm4m3l1_cc_w_0_300_s_3_300=1.38e-12 mcm4m3l1_cf_w_0_300_s_3_300=7.42e-11
+  mcm4m3l1_ca_w_0_300_s_9_000=2.18e-04 mcm4m3l1_cc_w_0_300_s_9_000=1.50e-14 mcm4m3l1_cf_w_0_300_s_9_000=7.57e-11
+  mcm4m3l1_ca_w_2_400_s_0_300=2.18e-04 mcm4m3l1_cc_w_2_400_s_0_300=1.01e-10 mcm4m3l1_cf_w_2_400_s_0_300=2.02e-11
+  mcm4m3l1_ca_w_2_400_s_0_360=2.18e-04 mcm4m3l1_cc_w_2_400_s_0_360=9.05e-11 mcm4m3l1_cf_w_2_400_s_0_360=2.41e-11
+  mcm4m3l1_ca_w_2_400_s_0_450=2.18e-04 mcm4m3l1_cc_w_2_400_s_0_450=7.69e-11 mcm4m3l1_cf_w_2_400_s_0_450=2.93e-11
+  mcm4m3l1_ca_w_2_400_s_0_600=2.18e-04 mcm4m3l1_cc_w_2_400_s_0_600=5.95e-11 mcm4m3l1_cf_w_2_400_s_0_600=3.69e-11
+  mcm4m3l1_ca_w_2_400_s_0_800=2.18e-04 mcm4m3l1_cc_w_2_400_s_0_800=4.28e-11 mcm4m3l1_cf_w_2_400_s_0_800=4.51e-11
+  mcm4m3l1_ca_w_2_400_s_1_000=2.18e-04 mcm4m3l1_cc_w_2_400_s_1_000=3.13e-11 mcm4m3l1_cf_w_2_400_s_1_000=5.17e-11
+  mcm4m3l1_ca_w_2_400_s_1_200=2.18e-04 mcm4m3l1_cc_w_2_400_s_1_200=2.31e-11 mcm4m3l1_cf_w_2_400_s_1_200=5.69e-11
+  mcm4m3l1_ca_w_2_400_s_2_100=2.18e-04 mcm4m3l1_cc_w_2_400_s_2_100=6.68e-12 mcm4m3l1_cf_w_2_400_s_2_100=6.99e-11
+  mcm4m3l1_ca_w_2_400_s_3_300=2.18e-04 mcm4m3l1_cc_w_2_400_s_3_300=1.45e-12 mcm4m3l1_cf_w_2_400_s_3_300=7.50e-11
+  mcm4m3l1_ca_w_2_400_s_9_000=2.18e-04 mcm4m3l1_cc_w_2_400_s_9_000=5.17e-26 mcm4m3l1_cf_w_2_400_s_9_000=7.65e-11
+  mcm4m3m1_ca_w_0_300_s_0_300=2.37e-04 mcm4m3m1_cc_w_0_300_s_0_300=9.39e-11 mcm4m3m1_cf_w_0_300_s_0_300=2.24e-11
+  mcm4m3m1_ca_w_0_300_s_0_360=2.37e-04 mcm4m3m1_cc_w_0_300_s_0_360=8.33e-11 mcm4m3m1_cf_w_0_300_s_0_360=2.67e-11
+  mcm4m3m1_ca_w_0_300_s_0_450=2.37e-04 mcm4m3m1_cc_w_0_300_s_0_450=7.01e-11 mcm4m3m1_cf_w_0_300_s_0_450=3.27e-11
+  mcm4m3m1_ca_w_0_300_s_0_600=2.37e-04 mcm4m3m1_cc_w_0_300_s_0_600=5.30e-11 mcm4m3m1_cf_w_0_300_s_0_600=4.12e-11
+  mcm4m3m1_ca_w_0_300_s_0_800=2.37e-04 mcm4m3m1_cc_w_0_300_s_0_800=3.69e-11 mcm4m3m1_cf_w_0_300_s_0_800=5.05e-11
+  mcm4m3m1_ca_w_0_300_s_1_000=2.37e-04 mcm4m3m1_cc_w_0_300_s_1_000=2.55e-11 mcm4m3m1_cf_w_0_300_s_1_000=5.78e-11
+  mcm4m3m1_ca_w_0_300_s_1_200=2.37e-04 mcm4m3m1_cc_w_0_300_s_1_200=1.79e-11 mcm4m3m1_cf_w_0_300_s_1_200=6.33e-11
+  mcm4m3m1_ca_w_0_300_s_2_100=2.37e-04 mcm4m3m1_cc_w_0_300_s_2_100=3.89e-12 mcm4m3m1_cf_w_0_300_s_2_100=7.53e-11
+  mcm4m3m1_ca_w_0_300_s_3_300=2.37e-04 mcm4m3m1_cc_w_0_300_s_3_300=5.95e-13 mcm4m3m1_cf_w_0_300_s_3_300=7.86e-11
+  mcm4m3m1_ca_w_0_300_s_9_000=2.37e-04 mcm4m3m1_cc_w_0_300_s_9_000=4.00e-14 mcm4m3m1_cf_w_0_300_s_9_000=7.92e-11
+  mcm4m3m1_ca_w_2_400_s_0_300=2.37e-04 mcm4m3m1_cc_w_2_400_s_0_300=9.55e-11 mcm4m3m1_cf_w_2_400_s_0_300=2.24e-11
+  mcm4m3m1_ca_w_2_400_s_0_360=2.37e-04 mcm4m3m1_cc_w_2_400_s_0_360=8.45e-11 mcm4m3m1_cf_w_2_400_s_0_360=2.67e-11
+  mcm4m3m1_ca_w_2_400_s_0_450=2.37e-04 mcm4m3m1_cc_w_2_400_s_0_450=7.10e-11 mcm4m3m1_cf_w_2_400_s_0_450=3.26e-11
+  mcm4m3m1_ca_w_2_400_s_0_600=2.37e-04 mcm4m3m1_cc_w_2_400_s_0_600=5.37e-11 mcm4m3m1_cf_w_2_400_s_0_600=4.12e-11
+  mcm4m3m1_ca_w_2_400_s_0_800=2.37e-04 mcm4m3m1_cc_w_2_400_s_0_800=3.73e-11 mcm4m3m1_cf_w_2_400_s_0_800=5.05e-11
+  mcm4m3m1_ca_w_2_400_s_1_000=2.37e-04 mcm4m3m1_cc_w_2_400_s_1_000=2.59e-11 mcm4m3m1_cf_w_2_400_s_1_000=5.78e-11
+  mcm4m3m1_ca_w_2_400_s_1_200=2.37e-04 mcm4m3m1_cc_w_2_400_s_1_200=1.81e-11 mcm4m3m1_cf_w_2_400_s_1_200=6.34e-11
+  mcm4m3m1_ca_w_2_400_s_2_100=2.37e-04 mcm4m3m1_cc_w_2_400_s_2_100=3.95e-12 mcm4m3m1_cf_w_2_400_s_2_100=7.56e-11
+  mcm4m3m1_ca_w_2_400_s_3_300=2.37e-04 mcm4m3m1_cc_w_2_400_s_3_300=6.00e-13 mcm4m3m1_cf_w_2_400_s_3_300=7.88e-11
+  mcm4m3m1_ca_w_2_400_s_9_000=2.37e-04 mcm4m3m1_cc_w_2_400_s_9_000=5.00e-14 mcm4m3m1_cf_w_2_400_s_9_000=7.95e-11
+  mcm4m3m2_ca_w_0_300_s_0_300=3.22e-04 mcm4m3m2_cc_w_0_300_s_0_300=8.37e-11 mcm4m3m2_cf_w_0_300_s_0_300=3.14e-11
+  mcm4m3m2_ca_w_0_300_s_0_360=3.22e-04 mcm4m3m2_cc_w_0_300_s_0_360=7.33e-11 mcm4m3m2_cf_w_0_300_s_0_360=3.73e-11
+  mcm4m3m2_ca_w_0_300_s_0_450=3.22e-04 mcm4m3m2_cc_w_0_300_s_0_450=6.01e-11 mcm4m3m2_cf_w_0_300_s_0_450=4.53e-11
+  mcm4m3m2_ca_w_0_300_s_0_600=3.22e-04 mcm4m3m2_cc_w_0_300_s_0_600=4.30e-11 mcm4m3m2_cf_w_0_300_s_0_600=5.65e-11
+  mcm4m3m2_ca_w_0_300_s_0_800=3.22e-04 mcm4m3m2_cc_w_0_300_s_0_800=2.77e-11 mcm4m3m2_cf_w_0_300_s_0_800=6.79e-11
+  mcm4m3m2_ca_w_0_300_s_1_000=3.22e-04 mcm4m3m2_cc_w_0_300_s_1_000=1.75e-11 mcm4m3m2_cf_w_0_300_s_1_000=7.63e-11
+  mcm4m3m2_ca_w_0_300_s_1_200=3.22e-04 mcm4m3m2_cc_w_0_300_s_1_200=1.09e-11 mcm4m3m2_cf_w_0_300_s_1_200=8.16e-11
+  mcm4m3m2_ca_w_0_300_s_2_100=3.22e-04 mcm4m3m2_cc_w_0_300_s_2_100=1.55e-12 mcm4m3m2_cf_w_0_300_s_2_100=9.09e-11
+  mcm4m3m2_ca_w_0_300_s_3_300=3.22e-04 mcm4m3m2_cc_w_0_300_s_3_300=2.00e-13 mcm4m3m2_cf_w_0_300_s_3_300=9.24e-11
+  mcm4m3m2_ca_w_0_300_s_9_000=3.22e-04 mcm4m3m2_cc_w_0_300_s_9_000=0.00e+00 mcm4m3m2_cf_w_0_300_s_9_000=9.26e-11
+  mcm4m3m2_ca_w_2_400_s_0_300=3.22e-04 mcm4m3m2_cc_w_2_400_s_0_300=8.39e-11 mcm4m3m2_cf_w_2_400_s_0_300=3.14e-11
+  mcm4m3m2_ca_w_2_400_s_0_360=3.22e-04 mcm4m3m2_cc_w_2_400_s_0_360=7.33e-11 mcm4m3m2_cf_w_2_400_s_0_360=3.74e-11
+  mcm4m3m2_ca_w_2_400_s_0_450=3.22e-04 mcm4m3m2_cc_w_2_400_s_0_450=5.99e-11 mcm4m3m2_cf_w_2_400_s_0_450=4.54e-11
+  mcm4m3m2_ca_w_2_400_s_0_600=3.22e-04 mcm4m3m2_cc_w_2_400_s_0_600=4.32e-11 mcm4m3m2_cf_w_2_400_s_0_600=5.65e-11
+  mcm4m3m2_ca_w_2_400_s_0_800=3.22e-04 mcm4m3m2_cc_w_2_400_s_0_800=2.77e-11 mcm4m3m2_cf_w_2_400_s_0_800=6.79e-11
+  mcm4m3m2_ca_w_2_400_s_1_000=3.22e-04 mcm4m3m2_cc_w_2_400_s_1_000=1.75e-11 mcm4m3m2_cf_w_2_400_s_1_000=7.66e-11
+  mcm4m3m2_ca_w_2_400_s_1_200=3.22e-04 mcm4m3m2_cc_w_2_400_s_1_200=1.09e-11 mcm4m3m2_cf_w_2_400_s_1_200=8.18e-11
+  mcm4m3m2_ca_w_2_400_s_2_100=3.22e-04 mcm4m3m2_cc_w_2_400_s_2_100=1.55e-12 mcm4m3m2_cf_w_2_400_s_2_100=9.09e-11
+  mcm4m3m2_ca_w_2_400_s_3_300=3.22e-04 mcm4m3m2_cc_w_2_400_s_3_300=2.00e-13 mcm4m3m2_cf_w_2_400_s_3_300=9.24e-11
+  mcm4m3m2_ca_w_2_400_s_9_000=3.22e-04 mcm4m3m2_cc_w_2_400_s_9_000=0.00e+00 mcm4m3m2_cf_w_2_400_s_9_000=9.27e-11
+  mcm5m3f_ca_w_0_300_s_0_300=4.08e-05 mcm5m3f_cc_w_0_300_s_0_300=1.18e-10 mcm5m3f_cf_w_0_300_s_0_300=4.99e-12
+  mcm5m3f_ca_w_0_300_s_0_360=4.08e-05 mcm5m3f_cc_w_0_300_s_0_360=1.08e-10 mcm5m3f_cf_w_0_300_s_0_360=6.15e-12
+  mcm5m3f_ca_w_0_300_s_0_450=4.08e-05 mcm5m3f_cc_w_0_300_s_0_450=9.44e-11 mcm5m3f_cf_w_0_300_s_0_450=7.88e-12
+  mcm5m3f_ca_w_0_300_s_0_600=4.08e-05 mcm5m3f_cc_w_0_300_s_0_600=7.77e-11 mcm5m3f_cf_w_0_300_s_0_600=1.07e-11
+  mcm5m3f_ca_w_0_300_s_0_800=4.08e-05 mcm5m3f_cc_w_0_300_s_0_800=6.14e-11 mcm5m3f_cf_w_0_300_s_0_800=1.41e-11
+  mcm5m3f_ca_w_0_300_s_1_000=4.08e-05 mcm5m3f_cc_w_0_300_s_1_000=4.92e-11 mcm5m3f_cf_w_0_300_s_1_000=1.75e-11
+  mcm5m3f_ca_w_0_300_s_1_200=4.08e-05 mcm5m3f_cc_w_0_300_s_1_200=4.03e-11 mcm5m3f_cf_w_0_300_s_1_200=2.05e-11
+  mcm5m3f_ca_w_0_300_s_2_100=4.08e-05 mcm5m3f_cc_w_0_300_s_2_100=1.90e-11 mcm5m3f_cf_w_0_300_s_2_100=3.16e-11
+  mcm5m3f_ca_w_0_300_s_3_300=4.08e-05 mcm5m3f_cc_w_0_300_s_3_300=7.81e-12 mcm5m3f_cf_w_0_300_s_3_300=4.00e-11
+  mcm5m3f_ca_w_0_300_s_9_000=4.08e-05 mcm5m3f_cc_w_0_300_s_9_000=1.55e-13 mcm5m3f_cf_w_0_300_s_9_000=4.71e-11
+  mcm5m3f_ca_w_2_400_s_0_300=4.08e-05 mcm5m3f_cc_w_2_400_s_0_300=1.28e-10 mcm5m3f_cf_w_2_400_s_0_300=5.05e-12
+  mcm5m3f_ca_w_2_400_s_0_360=4.08e-05 mcm5m3f_cc_w_2_400_s_0_360=1.17e-10 mcm5m3f_cf_w_2_400_s_0_360=6.20e-12
+  mcm5m3f_ca_w_2_400_s_0_450=4.08e-05 mcm5m3f_cc_w_2_400_s_0_450=1.02e-10 mcm5m3f_cf_w_2_400_s_0_450=7.90e-12
+  mcm5m3f_ca_w_2_400_s_0_600=4.08e-05 mcm5m3f_cc_w_2_400_s_0_600=8.40e-11 mcm5m3f_cf_w_2_400_s_0_600=1.07e-11
+  mcm5m3f_ca_w_2_400_s_0_800=4.08e-05 mcm5m3f_cc_w_2_400_s_0_800=6.61e-11 mcm5m3f_cf_w_2_400_s_0_800=1.42e-11
+  mcm5m3f_ca_w_2_400_s_1_000=4.08e-05 mcm5m3f_cc_w_2_400_s_1_000=5.32e-11 mcm5m3f_cf_w_2_400_s_1_000=1.76e-11
+  mcm5m3f_ca_w_2_400_s_1_200=4.08e-05 mcm5m3f_cc_w_2_400_s_1_200=4.36e-11 mcm5m3f_cf_w_2_400_s_1_200=2.08e-11
+  mcm5m3f_ca_w_2_400_s_2_100=4.08e-05 mcm5m3f_cc_w_2_400_s_2_100=2.06e-11 mcm5m3f_cf_w_2_400_s_2_100=3.22e-11
+  mcm5m3f_ca_w_2_400_s_3_300=4.08e-05 mcm5m3f_cc_w_2_400_s_3_300=8.60e-12 mcm5m3f_cf_w_2_400_s_3_300=4.12e-11
+  mcm5m3f_ca_w_2_400_s_9_000=4.08e-05 mcm5m3f_cc_w_2_400_s_9_000=1.55e-13 mcm5m3f_cf_w_2_400_s_9_000=4.90e-11
+  mcm5m3d_ca_w_0_300_s_0_300=4.26e-05 mcm5m3d_cc_w_0_300_s_0_300=1.17e-10 mcm5m3d_cf_w_0_300_s_0_300=5.21e-12
+  mcm5m3d_ca_w_0_300_s_0_360=4.26e-05 mcm5m3d_cc_w_0_300_s_0_360=1.07e-10 mcm5m3d_cf_w_0_300_s_0_360=6.41e-12
+  mcm5m3d_ca_w_0_300_s_0_450=4.26e-05 mcm5m3d_cc_w_0_300_s_0_450=9.39e-11 mcm5m3d_cf_w_0_300_s_0_450=8.22e-12
+  mcm5m3d_ca_w_0_300_s_0_600=4.26e-05 mcm5m3d_cc_w_0_300_s_0_600=7.71e-11 mcm5m3d_cf_w_0_300_s_0_600=1.11e-11
+  mcm5m3d_ca_w_0_300_s_0_800=4.26e-05 mcm5m3d_cc_w_0_300_s_0_800=6.08e-11 mcm5m3d_cf_w_0_300_s_0_800=1.47e-11
+  mcm5m3d_ca_w_0_300_s_1_000=4.26e-05 mcm5m3d_cc_w_0_300_s_1_000=4.86e-11 mcm5m3d_cf_w_0_300_s_1_000=1.82e-11
+  mcm5m3d_ca_w_0_300_s_1_200=4.26e-05 mcm5m3d_cc_w_0_300_s_1_200=3.96e-11 mcm5m3d_cf_w_0_300_s_1_200=2.14e-11
+  mcm5m3d_ca_w_0_300_s_2_100=4.26e-05 mcm5m3d_cc_w_0_300_s_2_100=1.82e-11 mcm5m3d_cf_w_0_300_s_2_100=3.27e-11
+  mcm5m3d_ca_w_0_300_s_3_300=4.26e-05 mcm5m3d_cc_w_0_300_s_3_300=7.23e-12 mcm5m3d_cf_w_0_300_s_3_300=4.11e-11
+  mcm5m3d_ca_w_0_300_s_9_000=4.26e-05 mcm5m3d_cc_w_0_300_s_9_000=1.70e-13 mcm5m3d_cf_w_0_300_s_9_000=4.77e-11
+  mcm5m3d_ca_w_2_400_s_0_300=4.26e-05 mcm5m3d_cc_w_2_400_s_0_300=1.26e-10 mcm5m3d_cf_w_2_400_s_0_300=5.28e-12
+  mcm5m3d_ca_w_2_400_s_0_360=4.26e-05 mcm5m3d_cc_w_2_400_s_0_360=1.15e-10 mcm5m3d_cf_w_2_400_s_0_360=6.48e-12
+  mcm5m3d_ca_w_2_400_s_0_450=4.26e-05 mcm5m3d_cc_w_2_400_s_0_450=1.01e-10 mcm5m3d_cf_w_2_400_s_0_450=8.25e-12
+  mcm5m3d_ca_w_2_400_s_0_600=4.26e-05 mcm5m3d_cc_w_2_400_s_0_600=8.29e-11 mcm5m3d_cf_w_2_400_s_0_600=1.11e-11
+  mcm5m3d_ca_w_2_400_s_0_800=4.26e-05 mcm5m3d_cc_w_2_400_s_0_800=6.50e-11 mcm5m3d_cf_w_2_400_s_0_800=1.48e-11
+  mcm5m3d_ca_w_2_400_s_1_000=4.26e-05 mcm5m3d_cc_w_2_400_s_1_000=5.21e-11 mcm5m3d_cf_w_2_400_s_1_000=1.84e-11
+  mcm5m3d_ca_w_2_400_s_1_200=4.26e-05 mcm5m3d_cc_w_2_400_s_1_200=4.25e-11 mcm5m3d_cf_w_2_400_s_1_200=2.16e-11
+  mcm5m3d_ca_w_2_400_s_2_100=4.26e-05 mcm5m3d_cc_w_2_400_s_2_100=1.96e-11 mcm5m3d_cf_w_2_400_s_2_100=3.33e-11
+  mcm5m3d_ca_w_2_400_s_3_300=4.26e-05 mcm5m3d_cc_w_2_400_s_3_300=7.83e-12 mcm5m3d_cf_w_2_400_s_3_300=4.23e-11
+  mcm5m3d_ca_w_2_400_s_9_000=4.26e-05 mcm5m3d_cc_w_2_400_s_9_000=1.55e-13 mcm5m3d_cf_w_2_400_s_9_000=4.94e-11
+  mcm5m3p1_ca_w_0_300_s_0_300=4.58e-05 mcm5m3p1_cc_w_0_300_s_0_300=1.16e-10 mcm5m3p1_cf_w_0_300_s_0_300=5.60e-12
+  mcm5m3p1_ca_w_0_300_s_0_360=4.58e-05 mcm5m3p1_cc_w_0_300_s_0_360=1.06e-10 mcm5m3p1_cf_w_0_300_s_0_360=6.90e-12
+  mcm5m3p1_ca_w_0_300_s_0_450=4.58e-05 mcm5m3p1_cc_w_0_300_s_0_450=9.30e-11 mcm5m3p1_cf_w_0_300_s_0_450=8.83e-12
+  mcm5m3p1_ca_w_0_300_s_0_600=4.58e-05 mcm5m3p1_cc_w_0_300_s_0_600=7.59e-11 mcm5m3p1_cf_w_0_300_s_0_600=1.19e-11
+  mcm5m3p1_ca_w_0_300_s_0_800=4.58e-05 mcm5m3p1_cc_w_0_300_s_0_800=5.96e-11 mcm5m3p1_cf_w_0_300_s_0_800=1.58e-11
+  mcm5m3p1_ca_w_0_300_s_1_000=4.58e-05 mcm5m3p1_cc_w_0_300_s_1_000=4.73e-11 mcm5m3p1_cf_w_0_300_s_1_000=1.95e-11
+  mcm5m3p1_ca_w_0_300_s_1_200=4.58e-05 mcm5m3p1_cc_w_0_300_s_1_200=3.83e-11 mcm5m3p1_cf_w_0_300_s_1_200=2.28e-11
+  mcm5m3p1_ca_w_0_300_s_2_100=4.58e-05 mcm5m3p1_cc_w_0_300_s_2_100=1.69e-11 mcm5m3p1_cf_w_0_300_s_2_100=3.46e-11
+  mcm5m3p1_ca_w_0_300_s_3_300=4.58e-05 mcm5m3p1_cc_w_0_300_s_3_300=6.36e-12 mcm5m3p1_cf_w_0_300_s_3_300=4.30e-11
+  mcm5m3p1_ca_w_0_300_s_9_000=4.58e-05 mcm5m3p1_cc_w_0_300_s_9_000=1.15e-13 mcm5m3p1_cf_w_0_300_s_9_000=4.89e-11
+  mcm5m3p1_ca_w_2_400_s_0_300=4.58e-05 mcm5m3p1_cc_w_2_400_s_0_300=1.25e-10 mcm5m3p1_cf_w_2_400_s_0_300=5.69e-12
+  mcm5m3p1_ca_w_2_400_s_0_360=4.58e-05 mcm5m3p1_cc_w_2_400_s_0_360=1.14e-10 mcm5m3p1_cf_w_2_400_s_0_360=6.99e-12
+  mcm5m3p1_ca_w_2_400_s_0_450=4.58e-05 mcm5m3p1_cc_w_2_400_s_0_450=9.94e-11 mcm5m3p1_cf_w_2_400_s_0_450=8.90e-12
+  mcm5m3p1_ca_w_2_400_s_0_600=4.58e-05 mcm5m3p1_cc_w_2_400_s_0_600=8.11e-11 mcm5m3p1_cf_w_2_400_s_0_600=1.20e-11
+  mcm5m3p1_ca_w_2_400_s_0_800=4.58e-05 mcm5m3p1_cc_w_2_400_s_0_800=6.32e-11 mcm5m3p1_cf_w_2_400_s_0_800=1.59e-11
+  mcm5m3p1_ca_w_2_400_s_1_000=4.58e-05 mcm5m3p1_cc_w_2_400_s_1_000=5.03e-11 mcm5m3p1_cf_w_2_400_s_1_000=1.97e-11
+  mcm5m3p1_ca_w_2_400_s_1_200=4.58e-05 mcm5m3p1_cc_w_2_400_s_1_200=4.07e-11 mcm5m3p1_cf_w_2_400_s_1_200=2.31e-11
+  mcm5m3p1_ca_w_2_400_s_2_100=4.58e-05 mcm5m3p1_cc_w_2_400_s_2_100=1.81e-11 mcm5m3p1_cf_w_2_400_s_2_100=3.52e-11
+  mcm5m3p1_ca_w_2_400_s_3_300=4.58e-05 mcm5m3p1_cc_w_2_400_s_3_300=6.84e-12 mcm5m3p1_cf_w_2_400_s_3_300=4.41e-11
+  mcm5m3p1_ca_w_2_400_s_9_000=4.58e-05 mcm5m3p1_cc_w_2_400_s_9_000=1.00e-13 mcm5m3p1_cf_w_2_400_s_9_000=5.04e-11
+  mcm5m3l1_ca_w_0_300_s_0_300=5.08e-05 mcm5m3l1_cc_w_0_300_s_0_300=1.15e-10 mcm5m3l1_cf_w_0_300_s_0_300=6.19e-12
+  mcm5m3l1_ca_w_0_300_s_0_360=5.08e-05 mcm5m3l1_cc_w_0_300_s_0_360=1.05e-10 mcm5m3l1_cf_w_0_300_s_0_360=7.62e-12
+  mcm5m3l1_ca_w_0_300_s_0_450=5.08e-05 mcm5m3l1_cc_w_0_300_s_0_450=9.15e-11 mcm5m3l1_cf_w_0_300_s_0_450=9.75e-12
+  mcm5m3l1_ca_w_0_300_s_0_600=5.08e-05 mcm5m3l1_cc_w_0_300_s_0_600=7.43e-11 mcm5m3l1_cf_w_0_300_s_0_600=1.31e-11
+  mcm5m3l1_ca_w_0_300_s_0_800=5.08e-05 mcm5m3l1_cc_w_0_300_s_0_800=5.80e-11 mcm5m3l1_cf_w_0_300_s_0_800=1.74e-11
+  mcm5m3l1_ca_w_0_300_s_1_000=5.08e-05 mcm5m3l1_cc_w_0_300_s_1_000=4.57e-11 mcm5m3l1_cf_w_0_300_s_1_000=2.13e-11
+  mcm5m3l1_ca_w_0_300_s_1_200=5.08e-05 mcm5m3l1_cc_w_0_300_s_1_200=3.65e-11 mcm5m3l1_cf_w_0_300_s_1_200=2.50e-11
+  mcm5m3l1_ca_w_0_300_s_2_100=5.08e-05 mcm5m3l1_cc_w_0_300_s_2_100=1.54e-11 mcm5m3l1_cf_w_0_300_s_2_100=3.73e-11
+  mcm5m3l1_ca_w_0_300_s_3_300=5.08e-05 mcm5m3l1_cc_w_0_300_s_3_300=5.36e-12 mcm5m3l1_cf_w_0_300_s_3_300=4.55e-11
+  mcm5m3l1_ca_w_0_300_s_9_000=5.08e-05 mcm5m3l1_cc_w_0_300_s_9_000=7.00e-14 mcm5m3l1_cf_w_0_300_s_9_000=5.06e-11
+  mcm5m3l1_ca_w_2_400_s_0_300=5.08e-05 mcm5m3l1_cc_w_2_400_s_0_300=1.22e-10 mcm5m3l1_cf_w_2_400_s_0_300=6.23e-12
+  mcm5m3l1_ca_w_2_400_s_0_360=5.08e-05 mcm5m3l1_cc_w_2_400_s_0_360=1.11e-10 mcm5m3l1_cf_w_2_400_s_0_360=7.66e-12
+  mcm5m3l1_ca_w_2_400_s_0_450=5.08e-05 mcm5m3l1_cc_w_2_400_s_0_450=9.70e-11 mcm5m3l1_cf_w_2_400_s_0_450=9.77e-12
+  mcm5m3l1_ca_w_2_400_s_0_600=5.08e-05 mcm5m3l1_cc_w_2_400_s_0_600=7.85e-11 mcm5m3l1_cf_w_2_400_s_0_600=1.31e-11
+  mcm5m3l1_ca_w_2_400_s_0_800=5.08e-05 mcm5m3l1_cc_w_2_400_s_0_800=6.10e-11 mcm5m3l1_cf_w_2_400_s_0_800=1.75e-11
+  mcm5m3l1_ca_w_2_400_s_1_000=5.08e-05 mcm5m3l1_cc_w_2_400_s_1_000=4.82e-11 mcm5m3l1_cf_w_2_400_s_1_000=2.15e-11
+  mcm5m3l1_ca_w_2_400_s_1_200=5.08e-05 mcm5m3l1_cc_w_2_400_s_1_200=3.86e-11 mcm5m3l1_cf_w_2_400_s_1_200=2.52e-11
+  mcm5m3l1_ca_w_2_400_s_2_100=5.08e-05 mcm5m3l1_cc_w_2_400_s_2_100=1.64e-11 mcm5m3l1_cf_w_2_400_s_2_100=3.79e-11
+  mcm5m3l1_ca_w_2_400_s_3_300=5.08e-05 mcm5m3l1_cc_w_2_400_s_3_300=5.70e-12 mcm5m3l1_cf_w_2_400_s_3_300=4.66e-11
+  mcm5m3l1_ca_w_2_400_s_9_000=5.08e-05 mcm5m3l1_cc_w_2_400_s_9_000=1.00e-13 mcm5m3l1_cf_w_2_400_s_9_000=5.19e-11
+  mcm5m3m1_ca_w_0_300_s_0_300=6.98e-05 mcm5m3m1_cc_w_0_300_s_0_300=1.12e-10 mcm5m3m1_cf_w_0_300_s_0_300=8.40e-12
+  mcm5m3m1_ca_w_0_300_s_0_360=6.98e-05 mcm5m3m1_cc_w_0_300_s_0_360=1.01e-10 mcm5m3m1_cf_w_0_300_s_0_360=1.03e-11
+  mcm5m3m1_ca_w_0_300_s_0_450=6.98e-05 mcm5m3m1_cc_w_0_300_s_0_450=8.75e-11 mcm5m3m1_cf_w_0_300_s_0_450=1.31e-11
+  mcm5m3m1_ca_w_0_300_s_0_600=6.98e-05 mcm5m3m1_cc_w_0_300_s_0_600=6.99e-11 mcm5m3m1_cf_w_0_300_s_0_600=1.75e-11
+  mcm5m3m1_ca_w_0_300_s_0_800=6.98e-05 mcm5m3m1_cc_w_0_300_s_0_800=5.33e-11 mcm5m3m1_cf_w_0_300_s_0_800=2.29e-11
+  mcm5m3m1_ca_w_0_300_s_1_000=6.98e-05 mcm5m3m1_cc_w_0_300_s_1_000=4.09e-11 mcm5m3m1_cf_w_0_300_s_1_000=2.78e-11
+  mcm5m3m1_ca_w_0_300_s_1_200=6.98e-05 mcm5m3m1_cc_w_0_300_s_1_200=3.19e-11 mcm5m3m1_cf_w_0_300_s_1_200=3.21e-11
+  mcm5m3m1_ca_w_0_300_s_2_100=6.98e-05 mcm5m3m1_cc_w_0_300_s_2_100=1.18e-11 mcm5m3m1_cf_w_0_300_s_2_100=4.54e-11
+  mcm5m3m1_ca_w_0_300_s_3_300=6.98e-05 mcm5m3m1_cc_w_0_300_s_3_300=3.44e-12 mcm5m3m1_cf_w_0_300_s_3_300=5.28e-11
+  mcm5m3m1_ca_w_0_300_s_9_000=6.98e-05 mcm5m3m1_cc_w_0_300_s_9_000=4.00e-14 mcm5m3m1_cf_w_0_300_s_9_000=5.61e-11
+  mcm5m3m1_ca_w_2_400_s_0_300=6.98e-05 mcm5m3m1_cc_w_2_400_s_0_300=1.17e-10 mcm5m3m1_cf_w_2_400_s_0_300=8.40e-12
+  mcm5m3m1_ca_w_2_400_s_0_360=6.98e-05 mcm5m3m1_cc_w_2_400_s_0_360=1.06e-10 mcm5m3m1_cf_w_2_400_s_0_360=1.03e-11
+  mcm5m3m1_ca_w_2_400_s_0_450=6.98e-05 mcm5m3m1_cc_w_2_400_s_0_450=9.13e-11 mcm5m3m1_cf_w_2_400_s_0_450=1.31e-11
+  mcm5m3m1_ca_w_2_400_s_0_600=6.98e-05 mcm5m3m1_cc_w_2_400_s_0_600=7.28e-11 mcm5m3m1_cf_w_2_400_s_0_600=1.75e-11
+  mcm5m3m1_ca_w_2_400_s_0_800=6.98e-05 mcm5m3m1_cc_w_2_400_s_0_800=5.54e-11 mcm5m3m1_cf_w_2_400_s_0_800=2.30e-11
+  mcm5m3m1_ca_w_2_400_s_1_000=6.98e-05 mcm5m3m1_cc_w_2_400_s_1_000=4.27e-11 mcm5m3m1_cf_w_2_400_s_1_000=2.80e-11
+  mcm5m3m1_ca_w_2_400_s_1_200=6.98e-05 mcm5m3m1_cc_w_2_400_s_1_200=3.33e-11 mcm5m3m1_cf_w_2_400_s_1_200=3.23e-11
+  mcm5m3m1_ca_w_2_400_s_2_100=6.98e-05 mcm5m3m1_cc_w_2_400_s_2_100=1.24e-11 mcm5m3m1_cf_w_2_400_s_2_100=4.60e-11
+  mcm5m3m1_ca_w_2_400_s_3_300=6.98e-05 mcm5m3m1_cc_w_2_400_s_3_300=3.60e-12 mcm5m3m1_cf_w_2_400_s_3_300=5.36e-11
+  mcm5m3m1_ca_w_2_400_s_9_000=6.98e-05 mcm5m3m1_cc_w_2_400_s_9_000=5.00e-14 mcm5m3m1_cf_w_2_400_s_9_000=5.71e-11
+  mcm5m3m2_ca_w_0_300_s_0_300=1.56e-04 mcm5m3m2_cc_w_0_300_s_0_300=1.01e-10 mcm5m3m2_cf_w_0_300_s_0_300=1.73e-11
+  mcm5m3m2_ca_w_0_300_s_0_360=1.56e-04 mcm5m3m2_cc_w_0_300_s_0_360=9.08e-11 mcm5m3m2_cf_w_0_300_s_0_360=2.09e-11
+  mcm5m3m2_ca_w_0_300_s_0_450=1.56e-04 mcm5m3m2_cc_w_0_300_s_0_450=7.73e-11 mcm5m3m2_cf_w_0_300_s_0_450=2.57e-11
+  mcm5m3m2_ca_w_0_300_s_0_600=1.56e-04 mcm5m3m2_cc_w_0_300_s_0_600=6.01e-11 mcm5m3m2_cf_w_0_300_s_0_600=3.28e-11
+  mcm5m3m2_ca_w_0_300_s_0_800=1.56e-04 mcm5m3m2_cc_w_0_300_s_0_800=4.39e-11 mcm5m3m2_cf_w_0_300_s_0_800=4.06e-11
+  mcm5m3m2_ca_w_0_300_s_1_000=1.56e-04 mcm5m3m2_cc_w_0_300_s_1_000=3.23e-11 mcm5m3m2_cf_w_0_300_s_1_000=4.70e-11
+  mcm5m3m2_ca_w_0_300_s_1_200=1.56e-04 mcm5m3m2_cc_w_0_300_s_1_200=2.41e-11 mcm5m3m2_cf_w_0_300_s_1_200=5.21e-11
+  mcm5m3m2_ca_w_0_300_s_2_100=1.56e-04 mcm5m3m2_cc_w_0_300_s_2_100=7.36e-12 mcm5m3m2_cf_w_0_300_s_2_100=6.53e-11
+  mcm5m3m2_ca_w_0_300_s_3_300=1.56e-04 mcm5m3m2_cc_w_0_300_s_3_300=1.66e-12 mcm5m3m2_cf_w_0_300_s_3_300=7.06e-11
+  mcm5m3m2_ca_w_0_300_s_9_000=1.56e-04 mcm5m3m2_cc_w_0_300_s_9_000=4.00e-14 mcm5m3m2_cf_w_0_300_s_9_000=7.25e-11
+  mcm5m3m2_ca_w_2_400_s_0_300=1.56e-04 mcm5m3m2_cc_w_2_400_s_0_300=1.05e-10 mcm5m3m2_cf_w_2_400_s_0_300=1.73e-11
+  mcm5m3m2_ca_w_2_400_s_0_360=1.56e-04 mcm5m3m2_cc_w_2_400_s_0_360=9.40e-11 mcm5m3m2_cf_w_2_400_s_0_360=2.08e-11
+  mcm5m3m2_ca_w_2_400_s_0_450=1.56e-04 mcm5m3m2_cc_w_2_400_s_0_450=8.03e-11 mcm5m3m2_cf_w_2_400_s_0_450=2.57e-11
+  mcm5m3m2_ca_w_2_400_s_0_600=1.56e-04 mcm5m3m2_cc_w_2_400_s_0_600=6.24e-11 mcm5m3m2_cf_w_2_400_s_0_600=3.28e-11
+  mcm5m3m2_ca_w_2_400_s_0_800=1.56e-04 mcm5m3m2_cc_w_2_400_s_0_800=4.56e-11 mcm5m3m2_cf_w_2_400_s_0_800=4.06e-11
+  mcm5m3m2_ca_w_2_400_s_1_000=1.56e-04 mcm5m3m2_cc_w_2_400_s_1_000=3.39e-11 mcm5m3m2_cf_w_2_400_s_1_000=4.72e-11
+  mcm5m3m2_ca_w_2_400_s_1_200=1.56e-04 mcm5m3m2_cc_w_2_400_s_1_200=2.53e-11 mcm5m3m2_cf_w_2_400_s_1_200=5.23e-11
+  mcm5m3m2_ca_w_2_400_s_2_100=1.56e-04 mcm5m3m2_cc_w_2_400_s_2_100=7.81e-12 mcm5m3m2_cf_w_2_400_s_2_100=6.57e-11
+  mcm5m3m2_ca_w_2_400_s_3_300=1.56e-04 mcm5m3m2_cc_w_2_400_s_3_300=1.86e-12 mcm5m3m2_cf_w_2_400_s_3_300=7.14e-11
+  mcm5m3m2_ca_w_2_400_s_9_000=1.56e-04 mcm5m3m2_cc_w_2_400_s_9_000=3.50e-14 mcm5m3m2_cf_w_2_400_s_9_000=7.34e-11
+  mcrdlm3f_ca_w_0_300_s_0_300=2.13e-05 mcrdlm3f_cc_w_0_300_s_0_300=1.22e-10 mcrdlm3f_cf_w_0_300_s_0_300=2.66e-12
+  mcrdlm3f_ca_w_0_300_s_0_360=2.13e-05 mcrdlm3f_cc_w_0_300_s_0_360=1.13e-10 mcrdlm3f_cf_w_0_300_s_0_360=3.28e-12
+  mcrdlm3f_ca_w_0_300_s_0_450=2.13e-05 mcrdlm3f_cc_w_0_300_s_0_450=1.00e-10 mcrdlm3f_cf_w_0_300_s_0_450=4.23e-12
+  mcrdlm3f_ca_w_0_300_s_0_600=2.13e-05 mcrdlm3f_cc_w_0_300_s_0_600=8.40e-11 mcrdlm3f_cf_w_0_300_s_0_600=5.77e-12
+  mcrdlm3f_ca_w_0_300_s_0_800=2.13e-05 mcrdlm3f_cc_w_0_300_s_0_800=6.90e-11 mcrdlm3f_cf_w_0_300_s_0_800=7.65e-12
+  mcrdlm3f_ca_w_0_300_s_1_000=2.13e-05 mcrdlm3f_cc_w_0_300_s_1_000=5.79e-11 mcrdlm3f_cf_w_0_300_s_1_000=9.55e-12
+  mcrdlm3f_ca_w_0_300_s_1_200=2.13e-05 mcrdlm3f_cc_w_0_300_s_1_200=4.96e-11 mcrdlm3f_cf_w_0_300_s_1_200=1.14e-11
+  mcrdlm3f_ca_w_0_300_s_2_100=2.13e-05 mcrdlm3f_cc_w_0_300_s_2_100=2.91e-11 mcrdlm3f_cf_w_0_300_s_2_100=1.88e-11
+  mcrdlm3f_ca_w_0_300_s_3_300=2.13e-05 mcrdlm3f_cc_w_0_300_s_3_300=1.71e-11 mcrdlm3f_cf_w_0_300_s_3_300=2.56e-11
+  mcrdlm3f_ca_w_0_300_s_9_000=2.13e-05 mcrdlm3f_cc_w_0_300_s_9_000=2.24e-12 mcrdlm3f_cf_w_0_300_s_9_000=3.77e-11
+  mcrdlm3f_ca_w_2_400_s_0_300=2.13e-05 mcrdlm3f_cc_w_2_400_s_0_300=1.42e-10 mcrdlm3f_cf_w_2_400_s_0_300=2.71e-12
+  mcrdlm3f_ca_w_2_400_s_0_360=2.13e-05 mcrdlm3f_cc_w_2_400_s_0_360=1.31e-10 mcrdlm3f_cf_w_2_400_s_0_360=3.33e-12
+  mcrdlm3f_ca_w_2_400_s_0_450=2.13e-05 mcrdlm3f_cc_w_2_400_s_0_450=1.17e-10 mcrdlm3f_cf_w_2_400_s_0_450=4.26e-12
+  mcrdlm3f_ca_w_2_400_s_0_600=2.13e-05 mcrdlm3f_cc_w_2_400_s_0_600=9.88e-11 mcrdlm3f_cf_w_2_400_s_0_600=5.78e-12
+  mcrdlm3f_ca_w_2_400_s_0_800=2.13e-05 mcrdlm3f_cc_w_2_400_s_0_800=8.12e-11 mcrdlm3f_cf_w_2_400_s_0_800=7.73e-12
+  mcrdlm3f_ca_w_2_400_s_1_000=2.13e-05 mcrdlm3f_cc_w_2_400_s_1_000=6.86e-11 mcrdlm3f_cf_w_2_400_s_1_000=9.65e-12
+  mcrdlm3f_ca_w_2_400_s_1_200=2.13e-05 mcrdlm3f_cc_w_2_400_s_1_200=5.90e-11 mcrdlm3f_cf_w_2_400_s_1_200=1.15e-11
+  mcrdlm3f_ca_w_2_400_s_2_100=2.13e-05 mcrdlm3f_cc_w_2_400_s_2_100=3.55e-11 mcrdlm3f_cf_w_2_400_s_2_100=1.89e-11
+  mcrdlm3f_ca_w_2_400_s_3_300=2.13e-05 mcrdlm3f_cc_w_2_400_s_3_300=2.13e-11 mcrdlm3f_cf_w_2_400_s_3_300=2.65e-11
+  mcrdlm3f_ca_w_2_400_s_9_000=2.13e-05 mcrdlm3f_cc_w_2_400_s_9_000=2.99e-12 mcrdlm3f_cf_w_2_400_s_9_000=4.09e-11
+  mcrdlm3d_ca_w_0_300_s_0_300=2.31e-05 mcrdlm3d_cc_w_0_300_s_0_300=1.22e-10 mcrdlm3d_cf_w_0_300_s_0_300=2.88e-12
+  mcrdlm3d_ca_w_0_300_s_0_360=2.31e-05 mcrdlm3d_cc_w_0_300_s_0_360=1.12e-10 mcrdlm3d_cf_w_0_300_s_0_360=3.55e-12
+  mcrdlm3d_ca_w_0_300_s_0_450=2.31e-05 mcrdlm3d_cc_w_0_300_s_0_450=9.99e-11 mcrdlm3d_cf_w_0_300_s_0_450=4.57e-12
+  mcrdlm3d_ca_w_0_300_s_0_600=2.31e-05 mcrdlm3d_cc_w_0_300_s_0_600=8.34e-11 mcrdlm3d_cf_w_0_300_s_0_600=6.22e-12
+  mcrdlm3d_ca_w_0_300_s_0_800=2.31e-05 mcrdlm3d_cc_w_0_300_s_0_800=6.83e-11 mcrdlm3d_cf_w_0_300_s_0_800=8.24e-12
+  mcrdlm3d_ca_w_0_300_s_1_000=2.31e-05 mcrdlm3d_cc_w_0_300_s_1_000=5.71e-11 mcrdlm3d_cf_w_0_300_s_1_000=1.03e-11
+  mcrdlm3d_ca_w_0_300_s_1_200=2.31e-05 mcrdlm3d_cc_w_0_300_s_1_200=4.88e-11 mcrdlm3d_cf_w_0_300_s_1_200=1.22e-11
+  mcrdlm3d_ca_w_0_300_s_2_100=2.31e-05 mcrdlm3d_cc_w_0_300_s_2_100=2.82e-11 mcrdlm3d_cf_w_0_300_s_2_100=2.00e-11
+  mcrdlm3d_ca_w_0_300_s_3_300=2.31e-05 mcrdlm3d_cc_w_0_300_s_3_300=1.63e-11 mcrdlm3d_cf_w_0_300_s_3_300=2.71e-11
+  mcrdlm3d_ca_w_0_300_s_9_000=2.31e-05 mcrdlm3d_cc_w_0_300_s_9_000=2.02e-12 mcrdlm3d_cf_w_0_300_s_9_000=3.89e-11
+  mcrdlm3d_ca_w_2_400_s_0_300=2.31e-05 mcrdlm3d_cc_w_2_400_s_0_300=1.41e-10 mcrdlm3d_cf_w_2_400_s_0_300=2.94e-12
+  mcrdlm3d_ca_w_2_400_s_0_360=2.31e-05 mcrdlm3d_cc_w_2_400_s_0_360=1.30e-10 mcrdlm3d_cf_w_2_400_s_0_360=3.61e-12
+  mcrdlm3d_ca_w_2_400_s_0_450=2.31e-05 mcrdlm3d_cc_w_2_400_s_0_450=1.16e-10 mcrdlm3d_cf_w_2_400_s_0_450=4.60e-12
+  mcrdlm3d_ca_w_2_400_s_0_600=2.31e-05 mcrdlm3d_cc_w_2_400_s_0_600=9.77e-11 mcrdlm3d_cf_w_2_400_s_0_600=6.24e-12
+  mcrdlm3d_ca_w_2_400_s_0_800=2.31e-05 mcrdlm3d_cc_w_2_400_s_0_800=8.02e-11 mcrdlm3d_cf_w_2_400_s_0_800=8.34e-12
+  mcrdlm3d_ca_w_2_400_s_1_000=2.31e-05 mcrdlm3d_cc_w_2_400_s_1_000=6.75e-11 mcrdlm3d_cf_w_2_400_s_1_000=1.04e-11
+  mcrdlm3d_ca_w_2_400_s_1_200=2.31e-05 mcrdlm3d_cc_w_2_400_s_1_200=5.79e-11 mcrdlm3d_cf_w_2_400_s_1_200=1.24e-11
+  mcrdlm3d_ca_w_2_400_s_2_100=2.31e-05 mcrdlm3d_cc_w_2_400_s_2_100=3.45e-11 mcrdlm3d_cf_w_2_400_s_2_100=2.01e-11
+  mcrdlm3d_ca_w_2_400_s_3_300=2.31e-05 mcrdlm3d_cc_w_2_400_s_3_300=2.04e-11 mcrdlm3d_cf_w_2_400_s_3_300=2.80e-11
+  mcrdlm3d_ca_w_2_400_s_9_000=2.31e-05 mcrdlm3d_cc_w_2_400_s_9_000=2.77e-12 mcrdlm3d_cf_w_2_400_s_9_000=4.21e-11
+  mcrdlm3p1_ca_w_0_300_s_0_300=2.63e-05 mcrdlm3p1_cc_w_0_300_s_0_300=1.21e-10 mcrdlm3p1_cf_w_0_300_s_0_300=3.28e-12
+  mcrdlm3p1_ca_w_0_300_s_0_360=2.63e-05 mcrdlm3p1_cc_w_0_300_s_0_360=1.12e-10 mcrdlm3p1_cf_w_0_300_s_0_360=4.04e-12
+  mcrdlm3p1_ca_w_0_300_s_0_450=2.63e-05 mcrdlm3p1_cc_w_0_300_s_0_450=9.90e-11 mcrdlm3p1_cf_w_0_300_s_0_450=5.18e-12
+  mcrdlm3p1_ca_w_0_300_s_0_600=2.63e-05 mcrdlm3p1_cc_w_0_300_s_0_600=8.24e-11 mcrdlm3p1_cf_w_0_300_s_0_600=7.04e-12
+  mcrdlm3p1_ca_w_0_300_s_0_800=2.63e-05 mcrdlm3p1_cc_w_0_300_s_0_800=6.72e-11 mcrdlm3p1_cf_w_0_300_s_0_800=9.31e-12
+  mcrdlm3p1_ca_w_0_300_s_1_000=2.63e-05 mcrdlm3p1_cc_w_0_300_s_1_000=5.59e-11 mcrdlm3p1_cf_w_0_300_s_1_000=1.16e-11
+  mcrdlm3p1_ca_w_0_300_s_1_200=2.63e-05 mcrdlm3p1_cc_w_0_300_s_1_200=4.74e-11 mcrdlm3p1_cf_w_0_300_s_1_200=1.37e-11
+  mcrdlm3p1_ca_w_0_300_s_2_100=2.63e-05 mcrdlm3p1_cc_w_0_300_s_2_100=2.68e-11 mcrdlm3p1_cf_w_0_300_s_2_100=2.21e-11
+  mcrdlm3p1_ca_w_0_300_s_3_300=2.63e-05 mcrdlm3p1_cc_w_0_300_s_3_300=1.51e-11 mcrdlm3p1_cf_w_0_300_s_3_300=2.94e-11
+  mcrdlm3p1_ca_w_0_300_s_9_000=2.63e-05 mcrdlm3p1_cc_w_0_300_s_9_000=1.73e-12 mcrdlm3p1_cf_w_0_300_s_9_000=4.08e-11
+  mcrdlm3p1_ca_w_2_400_s_0_300=2.63e-05 mcrdlm3p1_cc_w_2_400_s_0_300=1.39e-10 mcrdlm3p1_cf_w_2_400_s_0_300=3.38e-12
+  mcrdlm3p1_ca_w_2_400_s_0_360=2.63e-05 mcrdlm3p1_cc_w_2_400_s_0_360=1.28e-10 mcrdlm3p1_cf_w_2_400_s_0_360=4.12e-12
+  mcrdlm3p1_ca_w_2_400_s_0_450=2.63e-05 mcrdlm3p1_cc_w_2_400_s_0_450=1.14e-10 mcrdlm3p1_cf_w_2_400_s_0_450=5.25e-12
+  mcrdlm3p1_ca_w_2_400_s_0_600=2.63e-05 mcrdlm3p1_cc_w_2_400_s_0_600=9.58e-11 mcrdlm3p1_cf_w_2_400_s_0_600=7.09e-12
+  mcrdlm3p1_ca_w_2_400_s_0_800=2.63e-05 mcrdlm3p1_cc_w_2_400_s_0_800=7.83e-11 mcrdlm3p1_cf_w_2_400_s_0_800=9.44e-12
+  mcrdlm3p1_ca_w_2_400_s_1_000=2.63e-05 mcrdlm3p1_cc_w_2_400_s_1_000=6.57e-11 mcrdlm3p1_cf_w_2_400_s_1_000=1.17e-11
+  mcrdlm3p1_ca_w_2_400_s_1_200=2.63e-05 mcrdlm3p1_cc_w_2_400_s_1_200=5.61e-11 mcrdlm3p1_cf_w_2_400_s_1_200=1.39e-11
+  mcrdlm3p1_ca_w_2_400_s_2_100=2.63e-05 mcrdlm3p1_cc_w_2_400_s_2_100=3.29e-11 mcrdlm3p1_cf_w_2_400_s_2_100=2.23e-11
+  mcrdlm3p1_ca_w_2_400_s_3_300=2.63e-05 mcrdlm3p1_cc_w_2_400_s_3_300=1.90e-11 mcrdlm3p1_cf_w_2_400_s_3_300=3.04e-11
+  mcrdlm3p1_ca_w_2_400_s_9_000=2.63e-05 mcrdlm3p1_cc_w_2_400_s_9_000=2.41e-12 mcrdlm3p1_cf_w_2_400_s_9_000=4.41e-11
+  mcrdlm3l1_ca_w_0_300_s_0_300=3.13e-05 mcrdlm3l1_cc_w_0_300_s_0_300=1.20e-10 mcrdlm3l1_cf_w_0_300_s_0_300=3.86e-12
+  mcrdlm3l1_ca_w_0_300_s_0_360=3.13e-05 mcrdlm3l1_cc_w_0_300_s_0_360=1.11e-10 mcrdlm3l1_cf_w_0_300_s_0_360=4.75e-12
+  mcrdlm3l1_ca_w_0_300_s_0_450=3.13e-05 mcrdlm3l1_cc_w_0_300_s_0_450=9.76e-11 mcrdlm3l1_cf_w_0_300_s_0_450=6.09e-12
+  mcrdlm3l1_ca_w_0_300_s_0_600=3.13e-05 mcrdlm3l1_cc_w_0_300_s_0_600=8.09e-11 mcrdlm3l1_cf_w_0_300_s_0_600=8.24e-12
+  mcrdlm3l1_ca_w_0_300_s_0_800=3.13e-05 mcrdlm3l1_cc_w_0_300_s_0_800=6.55e-11 mcrdlm3l1_cf_w_0_300_s_0_800=1.09e-11
+  mcrdlm3l1_ca_w_0_300_s_1_000=3.13e-05 mcrdlm3l1_cc_w_0_300_s_1_000=5.41e-11 mcrdlm3l1_cf_w_0_300_s_1_000=1.35e-11
+  mcrdlm3l1_ca_w_0_300_s_1_200=3.13e-05 mcrdlm3l1_cc_w_0_300_s_1_200=4.56e-11 mcrdlm3l1_cf_w_0_300_s_1_200=1.59e-11
+  mcrdlm3l1_ca_w_0_300_s_2_100=3.13e-05 mcrdlm3l1_cc_w_0_300_s_2_100=2.51e-11 mcrdlm3l1_cf_w_0_300_s_2_100=2.51e-11
+  mcrdlm3l1_ca_w_0_300_s_3_300=3.13e-05 mcrdlm3l1_cc_w_0_300_s_3_300=1.36e-11 mcrdlm3l1_cf_w_0_300_s_3_300=3.27e-11
+  mcrdlm3l1_ca_w_0_300_s_9_000=3.13e-05 mcrdlm3l1_cc_w_0_300_s_9_000=1.45e-12 mcrdlm3l1_cf_w_0_300_s_9_000=4.33e-11
+  mcrdlm3l1_ca_w_2_400_s_0_300=3.13e-05 mcrdlm3l1_cc_w_2_400_s_0_300=1.37e-10 mcrdlm3l1_cf_w_2_400_s_0_300=3.90e-12
+  mcrdlm3l1_ca_w_2_400_s_0_360=3.13e-05 mcrdlm3l1_cc_w_2_400_s_0_360=1.26e-10 mcrdlm3l1_cf_w_2_400_s_0_360=4.79e-12
+  mcrdlm3l1_ca_w_2_400_s_0_450=3.13e-05 mcrdlm3l1_cc_w_2_400_s_0_450=1.12e-10 mcrdlm3l1_cf_w_2_400_s_0_450=6.11e-12
+  mcrdlm3l1_ca_w_2_400_s_0_600=3.13e-05 mcrdlm3l1_cc_w_2_400_s_0_600=9.35e-11 mcrdlm3l1_cf_w_2_400_s_0_600=8.25e-12
+  mcrdlm3l1_ca_w_2_400_s_0_800=3.13e-05 mcrdlm3l1_cc_w_2_400_s_0_800=7.61e-11 mcrdlm3l1_cf_w_2_400_s_0_800=1.10e-11
+  mcrdlm3l1_ca_w_2_400_s_1_000=3.13e-05 mcrdlm3l1_cc_w_2_400_s_1_000=6.34e-11 mcrdlm3l1_cf_w_2_400_s_1_000=1.36e-11
+  mcrdlm3l1_ca_w_2_400_s_1_200=3.13e-05 mcrdlm3l1_cc_w_2_400_s_1_200=5.39e-11 mcrdlm3l1_cf_w_2_400_s_1_200=1.60e-11
+  mcrdlm3l1_ca_w_2_400_s_2_100=3.13e-05 mcrdlm3l1_cc_w_2_400_s_2_100=3.08e-11 mcrdlm3l1_cf_w_2_400_s_2_100=2.52e-11
+  mcrdlm3l1_ca_w_2_400_s_3_300=3.13e-05 mcrdlm3l1_cc_w_2_400_s_3_300=1.74e-11 mcrdlm3l1_cf_w_2_400_s_3_300=3.37e-11
+  mcrdlm3l1_ca_w_2_400_s_9_000=3.13e-05 mcrdlm3l1_cc_w_2_400_s_9_000=2.03e-12 mcrdlm3l1_cf_w_2_400_s_9_000=4.67e-11
+  mcrdlm3m1_ca_w_0_300_s_0_300=5.02e-05 mcrdlm3m1_cc_w_0_300_s_0_300=1.16e-10 mcrdlm3m1_cf_w_0_300_s_0_300=6.06e-12
+  mcrdlm3m1_ca_w_0_300_s_0_360=5.02e-05 mcrdlm3m1_cc_w_0_300_s_0_360=1.06e-10 mcrdlm3m1_cf_w_0_300_s_0_360=7.43e-12
+  mcrdlm3m1_ca_w_0_300_s_0_450=5.02e-05 mcrdlm3m1_cc_w_0_300_s_0_450=9.33e-11 mcrdlm3m1_cf_w_0_300_s_0_450=9.44e-12
+  mcrdlm3m1_ca_w_0_300_s_0_600=5.02e-05 mcrdlm3m1_cc_w_0_300_s_0_600=7.63e-11 mcrdlm3m1_cf_w_0_300_s_0_600=1.26e-11
+  mcrdlm3m1_ca_w_0_300_s_0_800=5.02e-05 mcrdlm3m1_cc_w_0_300_s_0_800=6.08e-11 mcrdlm3m1_cf_w_0_300_s_0_800=1.64e-11
+  mcrdlm3m1_ca_w_0_300_s_1_000=5.02e-05 mcrdlm3m1_cc_w_0_300_s_1_000=4.93e-11 mcrdlm3m1_cf_w_0_300_s_1_000=2.00e-11
+  mcrdlm3m1_ca_w_0_300_s_1_200=5.02e-05 mcrdlm3m1_cc_w_0_300_s_1_200=4.09e-11 mcrdlm3m1_cf_w_0_300_s_1_200=2.32e-11
+  mcrdlm3m1_ca_w_0_300_s_2_100=5.02e-05 mcrdlm3m1_cc_w_0_300_s_2_100=2.07e-11 mcrdlm3m1_cf_w_0_300_s_2_100=3.43e-11
+  mcrdlm3m1_ca_w_0_300_s_3_300=5.02e-05 mcrdlm3m1_cc_w_0_300_s_3_300=1.04e-11 mcrdlm3m1_cf_w_0_300_s_3_300=4.20e-11
+  mcrdlm3m1_ca_w_0_300_s_9_000=5.02e-05 mcrdlm3m1_cc_w_0_300_s_9_000=9.15e-13 mcrdlm3m1_cf_w_0_300_s_9_000=5.07e-11
+  mcrdlm3m1_ca_w_2_400_s_0_300=5.02e-05 mcrdlm3m1_cc_w_2_400_s_0_300=1.31e-10 mcrdlm3m1_cf_w_2_400_s_0_300=6.07e-12
+  mcrdlm3m1_ca_w_2_400_s_0_360=5.02e-05 mcrdlm3m1_cc_w_2_400_s_0_360=1.20e-10 mcrdlm3m1_cf_w_2_400_s_0_360=7.44e-12
+  mcrdlm3m1_ca_w_2_400_s_0_450=5.02e-05 mcrdlm3m1_cc_w_2_400_s_0_450=1.06e-10 mcrdlm3m1_cf_w_2_400_s_0_450=9.43e-12
+  mcrdlm3m1_ca_w_2_400_s_0_600=5.02e-05 mcrdlm3m1_cc_w_2_400_s_0_600=8.76e-11 mcrdlm3m1_cf_w_2_400_s_0_600=1.26e-11
+  mcrdlm3m1_ca_w_2_400_s_0_800=5.02e-05 mcrdlm3m1_cc_w_2_400_s_0_800=7.03e-11 mcrdlm3m1_cf_w_2_400_s_0_800=1.65e-11
+  mcrdlm3m1_ca_w_2_400_s_1_000=5.02e-05 mcrdlm3m1_cc_w_2_400_s_1_000=5.79e-11 mcrdlm3m1_cf_w_2_400_s_1_000=2.01e-11
+  mcrdlm3m1_ca_w_2_400_s_1_200=5.02e-05 mcrdlm3m1_cc_w_2_400_s_1_200=4.84e-11 mcrdlm3m1_cf_w_2_400_s_1_200=2.33e-11
+  mcrdlm3m1_ca_w_2_400_s_2_100=5.02e-05 mcrdlm3m1_cc_w_2_400_s_2_100=2.64e-11 mcrdlm3m1_cf_w_2_400_s_2_100=3.44e-11
+  mcrdlm3m1_ca_w_2_400_s_3_300=5.02e-05 mcrdlm3m1_cc_w_2_400_s_3_300=1.41e-11 mcrdlm3m1_cf_w_2_400_s_3_300=4.32e-11
+  mcrdlm3m1_ca_w_2_400_s_9_000=5.02e-05 mcrdlm3m1_cc_w_2_400_s_9_000=1.45e-12 mcrdlm3m1_cf_w_2_400_s_9_000=5.46e-11
+  mcrdlm3m2_ca_w_0_300_s_0_300=1.36e-04 mcrdlm3m2_cc_w_0_300_s_0_300=1.06e-10 mcrdlm3m2_cf_w_0_300_s_0_300=1.50e-11
+  mcrdlm3m2_ca_w_0_300_s_0_360=1.36e-04 mcrdlm3m2_cc_w_0_300_s_0_360=9.60e-11 mcrdlm3m2_cf_w_0_300_s_0_360=1.80e-11
+  mcrdlm3m2_ca_w_0_300_s_0_450=1.36e-04 mcrdlm3m2_cc_w_0_300_s_0_450=8.30e-11 mcrdlm3m2_cf_w_0_300_s_0_450=2.21e-11
+  mcrdlm3m2_ca_w_0_300_s_0_600=1.36e-04 mcrdlm3m2_cc_w_0_300_s_0_600=6.66e-11 mcrdlm3m2_cf_w_0_300_s_0_600=2.79e-11
+  mcrdlm3m2_ca_w_0_300_s_0_800=1.36e-04 mcrdlm3m2_cc_w_0_300_s_0_800=5.13e-11 mcrdlm3m2_cf_w_0_300_s_0_800=3.42e-11
+  mcrdlm3m2_ca_w_0_300_s_1_000=1.36e-04 mcrdlm3m2_cc_w_0_300_s_1_000=4.06e-11 mcrdlm3m2_cf_w_0_300_s_1_000=3.95e-11
+  mcrdlm3m2_ca_w_0_300_s_1_200=1.36e-04 mcrdlm3m2_cc_w_0_300_s_1_200=3.28e-11 mcrdlm3m2_cf_w_0_300_s_1_200=4.37e-11
+  mcrdlm3m2_ca_w_0_300_s_2_100=1.36e-04 mcrdlm3m2_cc_w_0_300_s_2_100=1.49e-11 mcrdlm3m2_cf_w_0_300_s_2_100=5.62e-11
+  mcrdlm3m2_ca_w_0_300_s_3_300=1.36e-04 mcrdlm3m2_cc_w_0_300_s_3_300=6.96e-12 mcrdlm3m2_cf_w_0_300_s_3_300=6.30e-11
+  mcrdlm3m2_ca_w_0_300_s_9_000=1.36e-04 mcrdlm3m2_cc_w_0_300_s_9_000=5.60e-13 mcrdlm3m2_cf_w_0_300_s_9_000=6.92e-11
+  mcrdlm3m2_ca_w_2_400_s_0_300=1.36e-04 mcrdlm3m2_cc_w_2_400_s_0_300=1.19e-10 mcrdlm3m2_cf_w_2_400_s_0_300=1.50e-11
+  mcrdlm3m2_ca_w_2_400_s_0_360=1.36e-04 mcrdlm3m2_cc_w_2_400_s_0_360=1.08e-10 mcrdlm3m2_cf_w_2_400_s_0_360=1.80e-11
+  mcrdlm3m2_ca_w_2_400_s_0_450=1.36e-04 mcrdlm3m2_cc_w_2_400_s_0_450=9.49e-11 mcrdlm3m2_cf_w_2_400_s_0_450=2.20e-11
+  mcrdlm3m2_ca_w_2_400_s_0_600=1.36e-04 mcrdlm3m2_cc_w_2_400_s_0_600=7.72e-11 mcrdlm3m2_cf_w_2_400_s_0_600=2.79e-11
+  mcrdlm3m2_ca_w_2_400_s_0_800=1.36e-04 mcrdlm3m2_cc_w_2_400_s_0_800=6.05e-11 mcrdlm3m2_cf_w_2_400_s_0_800=3.42e-11
+  mcrdlm3m2_ca_w_2_400_s_1_000=1.36e-04 mcrdlm3m2_cc_w_2_400_s_1_000=4.89e-11 mcrdlm3m2_cf_w_2_400_s_1_000=3.95e-11
+  mcrdlm3m2_ca_w_2_400_s_1_200=1.36e-04 mcrdlm3m2_cc_w_2_400_s_1_200=4.03e-11 mcrdlm3m2_cf_w_2_400_s_1_200=4.38e-11
+  mcrdlm3m2_ca_w_2_400_s_2_100=1.36e-04 mcrdlm3m2_cc_w_2_400_s_2_100=2.07e-11 mcrdlm3m2_cf_w_2_400_s_2_100=5.65e-11
+  mcrdlm3m2_ca_w_2_400_s_3_300=1.36e-04 mcrdlm3m2_cc_w_2_400_s_3_300=1.05e-11 mcrdlm3m2_cf_w_2_400_s_3_300=6.48e-11
+  mcrdlm3m2_ca_w_2_400_s_9_000=1.36e-04 mcrdlm3m2_cc_w_2_400_s_9_000=9.10e-13 mcrdlm3m2_cf_w_2_400_s_9_000=7.37e-11
+  mcm5m4f_ca_w_0_300_s_0_300=1.26e-04 mcm5m4f_cc_w_0_300_s_0_300=1.06e-10 mcm5m4f_cf_w_0_300_s_0_300=1.31e-11
+  mcm5m4f_ca_w_0_300_s_0_360=1.26e-04 mcm5m4f_cc_w_0_300_s_0_360=9.61e-11 mcm5m4f_cf_w_0_300_s_0_360=1.58e-11
+  mcm5m4f_ca_w_0_300_s_0_450=1.26e-04 mcm5m4f_cc_w_0_300_s_0_450=8.29e-11 mcm5m4f_cf_w_0_300_s_0_450=1.96e-11
+  mcm5m4f_ca_w_0_300_s_0_600=1.26e-04 mcm5m4f_cc_w_0_300_s_0_600=6.61e-11 mcm5m4f_cf_w_0_300_s_0_600=2.52e-11
+  mcm5m4f_ca_w_0_300_s_0_800=1.26e-04 mcm5m4f_cc_w_0_300_s_0_800=5.03e-11 mcm5m4f_cf_w_0_300_s_0_800=3.14e-11
+  mcm5m4f_ca_w_0_300_s_1_000=1.26e-04 mcm5m4f_cc_w_0_300_s_1_000=3.90e-11 mcm5m4f_cf_w_0_300_s_1_000=3.68e-11
+  mcm5m4f_ca_w_0_300_s_1_200=1.26e-04 mcm5m4f_cc_w_0_300_s_1_200=3.08e-11 mcm5m4f_cf_w_0_300_s_1_200=4.11e-11
+  mcm5m4f_ca_w_0_300_s_2_100=1.26e-04 mcm5m4f_cc_w_0_300_s_2_100=1.26e-11 mcm5m4f_cf_w_0_300_s_2_100=5.38e-11
+  mcm5m4f_ca_w_0_300_s_3_300=1.26e-04 mcm5m4f_cc_w_0_300_s_3_300=4.56e-12 mcm5m4f_cf_w_0_300_s_3_300=6.06e-11
+  mcm5m4f_ca_w_0_300_s_9_000=1.26e-04 mcm5m4f_cc_w_0_300_s_9_000=1.35e-13 mcm5m4f_cf_w_0_300_s_9_000=6.50e-11
+  mcm5m4f_ca_w_2_400_s_0_300=1.26e-04 mcm5m4f_cc_w_2_400_s_0_300=1.15e-10 mcm5m4f_cf_w_2_400_s_0_300=1.31e-11
+  mcm5m4f_ca_w_2_400_s_0_360=1.26e-04 mcm5m4f_cc_w_2_400_s_0_360=1.04e-10 mcm5m4f_cf_w_2_400_s_0_360=1.58e-11
+  mcm5m4f_ca_w_2_400_s_0_450=1.26e-04 mcm5m4f_cc_w_2_400_s_0_450=9.01e-11 mcm5m4f_cf_w_2_400_s_0_450=1.95e-11
+  mcm5m4f_ca_w_2_400_s_0_600=1.26e-04 mcm5m4f_cc_w_2_400_s_0_600=7.25e-11 mcm5m4f_cf_w_2_400_s_0_600=2.51e-11
+  mcm5m4f_ca_w_2_400_s_0_800=1.26e-04 mcm5m4f_cc_w_2_400_s_0_800=5.55e-11 mcm5m4f_cf_w_2_400_s_0_800=3.14e-11
+  mcm5m4f_ca_w_2_400_s_1_000=1.26e-04 mcm5m4f_cc_w_2_400_s_1_000=4.33e-11 mcm5m4f_cf_w_2_400_s_1_000=3.68e-11
+  mcm5m4f_ca_w_2_400_s_1_200=1.26e-04 mcm5m4f_cc_w_2_400_s_1_200=3.44e-11 mcm5m4f_cf_w_2_400_s_1_200=4.12e-11
+  mcm5m4f_ca_w_2_400_s_2_100=1.26e-04 mcm5m4f_cc_w_2_400_s_2_100=1.48e-11 mcm5m4f_cf_w_2_400_s_2_100=5.42e-11
+  mcm5m4f_ca_w_2_400_s_3_300=1.26e-04 mcm5m4f_cc_w_2_400_s_3_300=5.71e-12 mcm5m4f_cf_w_2_400_s_3_300=6.20e-11
+  mcm5m4f_ca_w_2_400_s_9_000=1.26e-04 mcm5m4f_cc_w_2_400_s_9_000=1.30e-13 mcm5m4f_cf_w_2_400_s_9_000=6.74e-11
+  mcm5m4d_ca_w_0_300_s_0_300=1.26e-04 mcm5m4d_cc_w_0_300_s_0_300=1.06e-10 mcm5m4d_cf_w_0_300_s_0_300=1.32e-11
+  mcm5m4d_ca_w_0_300_s_0_360=1.26e-04 mcm5m4d_cc_w_0_300_s_0_360=9.59e-11 mcm5m4d_cf_w_0_300_s_0_360=1.59e-11
+  mcm5m4d_ca_w_0_300_s_0_450=1.26e-04 mcm5m4d_cc_w_0_300_s_0_450=8.27e-11 mcm5m4d_cf_w_0_300_s_0_450=1.97e-11
+  mcm5m4d_ca_w_0_300_s_0_600=1.26e-04 mcm5m4d_cc_w_0_300_s_0_600=6.58e-11 mcm5m4d_cf_w_0_300_s_0_600=2.54e-11
+  mcm5m4d_ca_w_0_300_s_0_800=1.26e-04 mcm5m4d_cc_w_0_300_s_0_800=5.00e-11 mcm5m4d_cf_w_0_300_s_0_800=3.17e-11
+  mcm5m4d_ca_w_0_300_s_1_000=1.26e-04 mcm5m4d_cc_w_0_300_s_1_000=3.87e-11 mcm5m4d_cf_w_0_300_s_1_000=3.71e-11
+  mcm5m4d_ca_w_0_300_s_1_200=1.26e-04 mcm5m4d_cc_w_0_300_s_1_200=3.04e-11 mcm5m4d_cf_w_0_300_s_1_200=4.14e-11
+  mcm5m4d_ca_w_0_300_s_2_100=1.26e-04 mcm5m4d_cc_w_0_300_s_2_100=1.21e-11 mcm5m4d_cf_w_0_300_s_2_100=5.41e-11
+  mcm5m4d_ca_w_0_300_s_3_300=1.26e-04 mcm5m4d_cc_w_0_300_s_3_300=4.32e-12 mcm5m4d_cf_w_0_300_s_3_300=6.10e-11
+  mcm5m4d_ca_w_0_300_s_9_000=1.26e-04 mcm5m4d_cc_w_0_300_s_9_000=1.10e-13 mcm5m4d_cf_w_0_300_s_9_000=6.52e-11
+  mcm5m4d_ca_w_2_400_s_0_300=1.26e-04 mcm5m4d_cc_w_2_400_s_0_300=1.14e-10 mcm5m4d_cf_w_2_400_s_0_300=1.32e-11
+  mcm5m4d_ca_w_2_400_s_0_360=1.26e-04 mcm5m4d_cc_w_2_400_s_0_360=1.04e-10 mcm5m4d_cf_w_2_400_s_0_360=1.59e-11
+  mcm5m4d_ca_w_2_400_s_0_450=1.26e-04 mcm5m4d_cc_w_2_400_s_0_450=8.96e-11 mcm5m4d_cf_w_2_400_s_0_450=1.97e-11
+  mcm5m4d_ca_w_2_400_s_0_600=1.26e-04 mcm5m4d_cc_w_2_400_s_0_600=7.18e-11 mcm5m4d_cf_w_2_400_s_0_600=2.53e-11
+  mcm5m4d_ca_w_2_400_s_0_800=1.26e-04 mcm5m4d_cc_w_2_400_s_0_800=5.48e-11 mcm5m4d_cf_w_2_400_s_0_800=3.17e-11
+  mcm5m4d_ca_w_2_400_s_1_000=1.26e-04 mcm5m4d_cc_w_2_400_s_1_000=4.26e-11 mcm5m4d_cf_w_2_400_s_1_000=3.71e-11
+  mcm5m4d_ca_w_2_400_s_1_200=1.26e-04 mcm5m4d_cc_w_2_400_s_1_200=3.38e-11 mcm5m4d_cf_w_2_400_s_1_200=4.16e-11
+  mcm5m4d_ca_w_2_400_s_2_100=1.26e-04 mcm5m4d_cc_w_2_400_s_2_100=1.42e-11 mcm5m4d_cf_w_2_400_s_2_100=5.46e-11
+  mcm5m4d_ca_w_2_400_s_3_300=1.26e-04 mcm5m4d_cc_w_2_400_s_3_300=5.32e-12 mcm5m4d_cf_w_2_400_s_3_300=6.24e-11
+  mcm5m4d_ca_w_2_400_s_9_000=1.26e-04 mcm5m4d_cc_w_2_400_s_9_000=8.50e-14 mcm5m4d_cf_w_2_400_s_9_000=6.74e-11
+  mcm5m4p1_ca_w_0_300_s_0_300=1.27e-04 mcm5m4p1_cc_w_0_300_s_0_300=1.06e-10 mcm5m4p1_cf_w_0_300_s_0_300=1.33e-11
+  mcm5m4p1_ca_w_0_300_s_0_360=1.27e-04 mcm5m4p1_cc_w_0_300_s_0_360=9.55e-11 mcm5m4p1_cf_w_0_300_s_0_360=1.61e-11
+  mcm5m4p1_ca_w_0_300_s_0_450=1.27e-04 mcm5m4p1_cc_w_0_300_s_0_450=8.26e-11 mcm5m4p1_cf_w_0_300_s_0_450=2.00e-11
+  mcm5m4p1_ca_w_0_300_s_0_600=1.27e-04 mcm5m4p1_cc_w_0_300_s_0_600=6.55e-11 mcm5m4p1_cf_w_0_300_s_0_600=2.57e-11
+  mcm5m4p1_ca_w_0_300_s_0_800=1.27e-04 mcm5m4p1_cc_w_0_300_s_0_800=4.95e-11 mcm5m4p1_cf_w_0_300_s_0_800=3.21e-11
+  mcm5m4p1_ca_w_0_300_s_1_000=1.27e-04 mcm5m4p1_cc_w_0_300_s_1_000=3.81e-11 mcm5m4p1_cf_w_0_300_s_1_000=3.75e-11
+  mcm5m4p1_ca_w_0_300_s_1_200=1.27e-04 mcm5m4p1_cc_w_0_300_s_1_200=2.98e-11 mcm5m4p1_cf_w_0_300_s_1_200=4.20e-11
+  mcm5m4p1_ca_w_0_300_s_2_100=1.27e-04 mcm5m4p1_cc_w_0_300_s_2_100=1.16e-11 mcm5m4p1_cf_w_0_300_s_2_100=5.48e-11
+  mcm5m4p1_ca_w_0_300_s_3_300=1.27e-04 mcm5m4p1_cc_w_0_300_s_3_300=4.02e-12 mcm5m4p1_cf_w_0_300_s_3_300=6.15e-11
+  mcm5m4p1_ca_w_0_300_s_9_000=1.27e-04 mcm5m4p1_cc_w_0_300_s_9_000=6.50e-14 mcm5m4p1_cf_w_0_300_s_9_000=6.54e-11
+  mcm5m4p1_ca_w_2_400_s_0_300=1.27e-04 mcm5m4p1_cc_w_2_400_s_0_300=1.13e-10 mcm5m4p1_cf_w_2_400_s_0_300=1.34e-11
+  mcm5m4p1_ca_w_2_400_s_0_360=1.27e-04 mcm5m4p1_cc_w_2_400_s_0_360=1.03e-10 mcm5m4p1_cf_w_2_400_s_0_360=1.61e-11
+  mcm5m4p1_ca_w_2_400_s_0_450=1.27e-04 mcm5m4p1_cc_w_2_400_s_0_450=8.86e-11 mcm5m4p1_cf_w_2_400_s_0_450=1.99e-11
+  mcm5m4p1_ca_w_2_400_s_0_600=1.27e-04 mcm5m4p1_cc_w_2_400_s_0_600=7.08e-11 mcm5m4p1_cf_w_2_400_s_0_600=2.56e-11
+  mcm5m4p1_ca_w_2_400_s_0_800=1.27e-04 mcm5m4p1_cc_w_2_400_s_0_800=5.38e-11 mcm5m4p1_cf_w_2_400_s_0_800=3.21e-11
+  mcm5m4p1_ca_w_2_400_s_1_000=1.27e-04 mcm5m4p1_cc_w_2_400_s_1_000=4.16e-11 mcm5m4p1_cf_w_2_400_s_1_000=3.77e-11
+  mcm5m4p1_ca_w_2_400_s_1_200=1.27e-04 mcm5m4p1_cc_w_2_400_s_1_200=3.29e-11 mcm5m4p1_cf_w_2_400_s_1_200=4.21e-11
+  mcm5m4p1_ca_w_2_400_s_2_100=1.27e-04 mcm5m4p1_cc_w_2_400_s_2_100=1.34e-11 mcm5m4p1_cf_w_2_400_s_2_100=5.53e-11
+  mcm5m4p1_ca_w_2_400_s_3_300=1.27e-04 mcm5m4p1_cc_w_2_400_s_3_300=4.73e-12 mcm5m4p1_cf_w_2_400_s_3_300=6.29e-11
+  mcm5m4p1_ca_w_2_400_s_9_000=1.27e-04 mcm5m4p1_cc_w_2_400_s_9_000=6.50e-14 mcm5m4p1_cf_w_2_400_s_9_000=6.74e-11
+  mcm5m4l1_ca_w_0_300_s_0_300=1.29e-04 mcm5m4l1_cc_w_0_300_s_0_300=1.06e-10 mcm5m4l1_cf_w_0_300_s_0_300=1.35e-11
+  mcm5m4l1_ca_w_0_300_s_0_360=1.29e-04 mcm5m4l1_cc_w_0_300_s_0_360=9.51e-11 mcm5m4l1_cf_w_0_300_s_0_360=1.63e-11
+  mcm5m4l1_ca_w_0_300_s_0_450=1.29e-04 mcm5m4l1_cc_w_0_300_s_0_450=8.21e-11 mcm5m4l1_cf_w_0_300_s_0_450=2.02e-11
+  mcm5m4l1_ca_w_0_300_s_0_600=1.29e-04 mcm5m4l1_cc_w_0_300_s_0_600=6.49e-11 mcm5m4l1_cf_w_0_300_s_0_600=2.61e-11
+  mcm5m4l1_ca_w_0_300_s_0_800=1.29e-04 mcm5m4l1_cc_w_0_300_s_0_800=4.89e-11 mcm5m4l1_cf_w_0_300_s_0_800=3.26e-11
+  mcm5m4l1_ca_w_0_300_s_1_000=1.29e-04 mcm5m4l1_cc_w_0_300_s_1_000=3.75e-11 mcm5m4l1_cf_w_0_300_s_1_000=3.82e-11
+  mcm5m4l1_ca_w_0_300_s_1_200=1.29e-04 mcm5m4l1_cc_w_0_300_s_1_200=2.91e-11 mcm5m4l1_cf_w_0_300_s_1_200=4.27e-11
+  mcm5m4l1_ca_w_0_300_s_2_100=1.29e-04 mcm5m4l1_cc_w_0_300_s_2_100=1.11e-11 mcm5m4l1_cf_w_0_300_s_2_100=5.55e-11
+  mcm5m4l1_ca_w_0_300_s_3_300=1.29e-04 mcm5m4l1_cc_w_0_300_s_3_300=3.57e-12 mcm5m4l1_cf_w_0_300_s_3_300=6.22e-11
+  mcm5m4l1_ca_w_0_300_s_9_000=1.29e-04 mcm5m4l1_cc_w_0_300_s_9_000=6.50e-14 mcm5m4l1_cf_w_0_300_s_9_000=6.57e-11
+  mcm5m4l1_ca_w_2_400_s_0_300=1.29e-04 mcm5m4l1_cc_w_2_400_s_0_300=1.12e-10 mcm5m4l1_cf_w_2_400_s_0_300=1.35e-11
+  mcm5m4l1_ca_w_2_400_s_0_360=1.29e-04 mcm5m4l1_cc_w_2_400_s_0_360=1.01e-10 mcm5m4l1_cf_w_2_400_s_0_360=1.63e-11
+  mcm5m4l1_ca_w_2_400_s_0_450=1.29e-04 mcm5m4l1_cc_w_2_400_s_0_450=8.76e-11 mcm5m4l1_cf_w_2_400_s_0_450=2.02e-11
+  mcm5m4l1_ca_w_2_400_s_0_600=1.29e-04 mcm5m4l1_cc_w_2_400_s_0_600=6.96e-11 mcm5m4l1_cf_w_2_400_s_0_600=2.60e-11
+  mcm5m4l1_ca_w_2_400_s_0_800=1.29e-04 mcm5m4l1_cc_w_2_400_s_0_800=5.27e-11 mcm5m4l1_cf_w_2_400_s_0_800=3.26e-11
+  mcm5m4l1_ca_w_2_400_s_1_000=1.29e-04 mcm5m4l1_cc_w_2_400_s_1_000=4.05e-11 mcm5m4l1_cf_w_2_400_s_1_000=3.83e-11
+  mcm5m4l1_ca_w_2_400_s_1_200=1.29e-04 mcm5m4l1_cc_w_2_400_s_1_200=3.18e-11 mcm5m4l1_cf_w_2_400_s_1_200=4.29e-11
+  mcm5m4l1_ca_w_2_400_s_2_100=1.29e-04 mcm5m4l1_cc_w_2_400_s_2_100=1.24e-11 mcm5m4l1_cf_w_2_400_s_2_100=5.61e-11
+  mcm5m4l1_ca_w_2_400_s_3_300=1.29e-04 mcm5m4l1_cc_w_2_400_s_3_300=4.16e-12 mcm5m4l1_cf_w_2_400_s_3_300=6.35e-11
+  mcm5m4l1_ca_w_2_400_s_9_000=1.29e-04 mcm5m4l1_cc_w_2_400_s_9_000=6.50e-14 mcm5m4l1_cf_w_2_400_s_9_000=6.75e-11
+  mcm5m4m1_ca_w_0_300_s_0_300=1.33e-04 mcm5m4m1_cc_w_0_300_s_0_300=1.04e-10 mcm5m4m1_cf_w_0_300_s_0_300=1.40e-11
+  mcm5m4m1_ca_w_0_300_s_0_360=1.33e-04 mcm5m4m1_cc_w_0_300_s_0_360=9.40e-11 mcm5m4m1_cf_w_0_300_s_0_360=1.70e-11
+  mcm5m4m1_ca_w_0_300_s_0_450=1.33e-04 mcm5m4m1_cc_w_0_300_s_0_450=8.07e-11 mcm5m4m1_cf_w_0_300_s_0_450=2.10e-11
+  mcm5m4m1_ca_w_0_300_s_0_600=1.33e-04 mcm5m4m1_cc_w_0_300_s_0_600=6.37e-11 mcm5m4m1_cf_w_0_300_s_0_600=2.71e-11
+  mcm5m4m1_ca_w_0_300_s_0_800=1.33e-04 mcm5m4m1_cc_w_0_300_s_0_800=4.73e-11 mcm5m4m1_cf_w_0_300_s_0_800=3.40e-11
+  mcm5m4m1_ca_w_0_300_s_1_000=1.33e-04 mcm5m4m1_cc_w_0_300_s_1_000=3.58e-11 mcm5m4m1_cf_w_0_300_s_1_000=3.98e-11
+  mcm5m4m1_ca_w_0_300_s_1_200=1.33e-04 mcm5m4m1_cc_w_0_300_s_1_200=2.74e-11 mcm5m4m1_cf_w_0_300_s_1_200=4.45e-11
+  mcm5m4m1_ca_w_0_300_s_2_100=1.33e-04 mcm5m4m1_cc_w_0_300_s_2_100=9.50e-12 mcm5m4m1_cf_w_0_300_s_2_100=5.75e-11
+  mcm5m4m1_ca_w_0_300_s_3_300=1.33e-04 mcm5m4m1_cc_w_0_300_s_3_300=2.66e-12 mcm5m4m1_cf_w_0_300_s_3_300=6.39e-11
+  mcm5m4m1_ca_w_0_300_s_9_000=1.33e-04 mcm5m4m1_cc_w_0_300_s_9_000=1.00e-14 mcm5m4m1_cf_w_0_300_s_9_000=6.65e-11
+  mcm5m4m1_ca_w_2_400_s_0_300=1.33e-04 mcm5m4m1_cc_w_2_400_s_0_300=1.10e-10 mcm5m4m1_cf_w_2_400_s_0_300=1.40e-11
+  mcm5m4m1_ca_w_2_400_s_0_360=1.33e-04 mcm5m4m1_cc_w_2_400_s_0_360=9.87e-11 mcm5m4m1_cf_w_2_400_s_0_360=1.69e-11
+  mcm5m4m1_ca_w_2_400_s_0_450=1.33e-04 mcm5m4m1_cc_w_2_400_s_0_450=8.49e-11 mcm5m4m1_cf_w_2_400_s_0_450=2.10e-11
+  mcm5m4m1_ca_w_2_400_s_0_600=1.33e-04 mcm5m4m1_cc_w_2_400_s_0_600=6.69e-11 mcm5m4m1_cf_w_2_400_s_0_600=2.71e-11
+  mcm5m4m1_ca_w_2_400_s_0_800=1.33e-04 mcm5m4m1_cc_w_2_400_s_0_800=5.00e-11 mcm5m4m1_cf_w_2_400_s_0_800=3.40e-11
+  mcm5m4m1_ca_w_2_400_s_1_000=1.33e-04 mcm5m4m1_cc_w_2_400_s_1_000=3.79e-11 mcm5m4m1_cf_w_2_400_s_1_000=3.99e-11
+  mcm5m4m1_ca_w_2_400_s_1_200=1.33e-04 mcm5m4m1_cc_w_2_400_s_1_200=2.92e-11 mcm5m4m1_cf_w_2_400_s_1_200=4.47e-11
+  mcm5m4m1_ca_w_2_400_s_2_100=1.33e-04 mcm5m4m1_cc_w_2_400_s_2_100=1.03e-11 mcm5m4m1_cf_w_2_400_s_2_100=5.81e-11
+  mcm5m4m1_ca_w_2_400_s_3_300=1.33e-04 mcm5m4m1_cc_w_2_400_s_3_300=2.97e-12 mcm5m4m1_cf_w_2_400_s_3_300=6.49e-11
+  mcm5m4m1_ca_w_2_400_s_9_000=1.33e-04 mcm5m4m1_cc_w_2_400_s_9_000=6.00e-14 mcm5m4m1_cf_w_2_400_s_9_000=6.78e-11
+  mcm5m4m2_ca_w_0_300_s_0_300=1.40e-04 mcm5m4m2_cc_w_0_300_s_0_300=1.03e-10 mcm5m4m2_cf_w_0_300_s_0_300=1.48e-11
+  mcm5m4m2_ca_w_0_300_s_0_360=1.40e-04 mcm5m4m2_cc_w_0_300_s_0_360=9.25e-11 mcm5m4m2_cf_w_0_300_s_0_360=1.79e-11
+  mcm5m4m2_ca_w_0_300_s_0_450=1.40e-04 mcm5m4m2_cc_w_0_300_s_0_450=7.90e-11 mcm5m4m2_cf_w_0_300_s_0_450=2.23e-11
+  mcm5m4m2_ca_w_0_300_s_0_600=1.40e-04 mcm5m4m2_cc_w_0_300_s_0_600=6.17e-11 mcm5m4m2_cf_w_0_300_s_0_600=2.87e-11
+  mcm5m4m2_ca_w_0_300_s_0_800=1.40e-04 mcm5m4m2_cc_w_0_300_s_0_800=4.51e-11 mcm5m4m2_cf_w_0_300_s_0_800=3.61e-11
+  mcm5m4m2_ca_w_0_300_s_1_000=1.40e-04 mcm5m4m2_cc_w_0_300_s_1_000=3.34e-11 mcm5m4m2_cf_w_0_300_s_1_000=4.24e-11
+  mcm5m4m2_ca_w_0_300_s_1_200=1.40e-04 mcm5m4m2_cc_w_0_300_s_1_200=2.51e-11 mcm5m4m2_cf_w_0_300_s_1_200=4.73e-11
+  mcm5m4m2_ca_w_0_300_s_2_100=1.40e-04 mcm5m4m2_cc_w_0_300_s_2_100=7.73e-12 mcm5m4m2_cf_w_0_300_s_2_100=6.05e-11
+  mcm5m4m2_ca_w_0_300_s_3_300=1.40e-04 mcm5m4m2_cc_w_0_300_s_3_300=1.81e-12 mcm5m4m2_cf_w_0_300_s_3_300=6.61e-11
+  mcm5m4m2_ca_w_0_300_s_9_000=1.40e-04 mcm5m4m2_cc_w_0_300_s_9_000=3.00e-14 mcm5m4m2_cf_w_0_300_s_9_000=6.79e-11
+  mcm5m4m2_ca_w_2_400_s_0_300=1.40e-04 mcm5m4m2_cc_w_2_400_s_0_300=1.06e-10 mcm5m4m2_cf_w_2_400_s_0_300=1.48e-11
+  mcm5m4m2_ca_w_2_400_s_0_360=1.40e-04 mcm5m4m2_cc_w_2_400_s_0_360=9.55e-11 mcm5m4m2_cf_w_2_400_s_0_360=1.79e-11
+  mcm5m4m2_ca_w_2_400_s_0_450=1.40e-04 mcm5m4m2_cc_w_2_400_s_0_450=8.17e-11 mcm5m4m2_cf_w_2_400_s_0_450=2.23e-11
+  mcm5m4m2_ca_w_2_400_s_0_600=1.40e-04 mcm5m4m2_cc_w_2_400_s_0_600=6.37e-11 mcm5m4m2_cf_w_2_400_s_0_600=2.88e-11
+  mcm5m4m2_ca_w_2_400_s_0_800=1.40e-04 mcm5m4m2_cc_w_2_400_s_0_800=4.67e-11 mcm5m4m2_cf_w_2_400_s_0_800=3.62e-11
+  mcm5m4m2_ca_w_2_400_s_1_000=1.40e-04 mcm5m4m2_cc_w_2_400_s_1_000=3.47e-11 mcm5m4m2_cf_w_2_400_s_1_000=4.25e-11
+  mcm5m4m2_ca_w_2_400_s_1_200=1.40e-04 mcm5m4m2_cc_w_2_400_s_1_200=2.60e-11 mcm5m4m2_cf_w_2_400_s_1_200=4.75e-11
+  mcm5m4m2_ca_w_2_400_s_2_100=1.40e-04 mcm5m4m2_cc_w_2_400_s_2_100=8.12e-12 mcm5m4m2_cf_w_2_400_s_2_100=6.10e-11
+  mcm5m4m2_ca_w_2_400_s_3_300=1.40e-04 mcm5m4m2_cc_w_2_400_s_3_300=1.95e-12 mcm5m4m2_cf_w_2_400_s_3_300=6.68e-11
+  mcm5m4m2_ca_w_2_400_s_9_000=1.40e-04 mcm5m4m2_cc_w_2_400_s_9_000=5.00e-14 mcm5m4m2_cf_w_2_400_s_9_000=6.87e-11
+  mcm5m4m3_ca_w_0_300_s_0_300=3.06e-04 mcm5m4m3_cc_w_0_300_s_0_300=8.45e-11 mcm5m4m3_cf_w_0_300_s_0_300=3.14e-11
+  mcm5m4m3_ca_w_0_300_s_0_360=3.06e-04 mcm5m4m3_cc_w_0_300_s_0_360=7.39e-11 mcm5m4m3_cf_w_0_300_s_0_360=3.74e-11
+  mcm5m4m3_ca_w_0_300_s_0_450=3.06e-04 mcm5m4m3_cc_w_0_300_s_0_450=6.05e-11 mcm5m4m3_cf_w_0_300_s_0_450=4.53e-11
+  mcm5m4m3_ca_w_0_300_s_0_600=3.06e-04 mcm5m4m3_cc_w_0_300_s_0_600=4.39e-11 mcm5m4m3_cf_w_0_300_s_0_600=5.64e-11
+  mcm5m4m3_ca_w_0_300_s_0_800=3.06e-04 mcm5m4m3_cc_w_0_300_s_0_800=2.85e-11 mcm5m4m3_cf_w_0_300_s_0_800=6.76e-11
+  mcm5m4m3_ca_w_0_300_s_1_000=3.06e-04 mcm5m4m3_cc_w_0_300_s_1_000=1.80e-11 mcm5m4m3_cf_w_0_300_s_1_000=7.66e-11
+  mcm5m4m3_ca_w_0_300_s_1_200=3.06e-04 mcm5m4m3_cc_w_0_300_s_1_200=1.13e-11 mcm5m4m3_cf_w_0_300_s_1_200=8.19e-11
+  mcm5m4m3_ca_w_0_300_s_2_100=3.06e-04 mcm5m4m3_cc_w_0_300_s_2_100=1.65e-12 mcm5m4m3_cf_w_0_300_s_2_100=9.09e-11
+  mcm5m4m3_ca_w_0_300_s_3_300=3.06e-04 mcm5m4m3_cc_w_0_300_s_3_300=2.50e-13 mcm5m4m3_cf_w_0_300_s_3_300=9.31e-11
+  mcm5m4m3_ca_w_0_300_s_9_000=3.06e-04 mcm5m4m3_cc_w_0_300_s_9_000=0.00e+00 mcm5m4m3_cf_w_0_300_s_9_000=9.33e-11
+  mcm5m4m3_ca_w_2_400_s_0_300=3.06e-04 mcm5m4m3_cc_w_2_400_s_0_300=8.50e-11 mcm5m4m3_cf_w_2_400_s_0_300=3.14e-11
+  mcm5m4m3_ca_w_2_400_s_0_360=3.06e-04 mcm5m4m3_cc_w_2_400_s_0_360=7.43e-11 mcm5m4m3_cf_w_2_400_s_0_360=3.73e-11
+  mcm5m4m3_ca_w_2_400_s_0_450=3.06e-04 mcm5m4m3_cc_w_2_400_s_0_450=6.08e-11 mcm5m4m3_cf_w_2_400_s_0_450=4.53e-11
+  mcm5m4m3_ca_w_2_400_s_0_600=3.06e-04 mcm5m4m3_cc_w_2_400_s_0_600=4.39e-11 mcm5m4m3_cf_w_2_400_s_0_600=5.64e-11
+  mcm5m4m3_ca_w_2_400_s_0_800=3.06e-04 mcm5m4m3_cc_w_2_400_s_0_800=2.86e-11 mcm5m4m3_cf_w_2_400_s_0_800=6.77e-11
+  mcm5m4m3_ca_w_2_400_s_1_000=3.06e-04 mcm5m4m3_cc_w_2_400_s_1_000=1.80e-11 mcm5m4m3_cf_w_2_400_s_1_000=7.63e-11
+  mcm5m4m3_ca_w_2_400_s_1_200=3.06e-04 mcm5m4m3_cc_w_2_400_s_1_200=1.13e-11 mcm5m4m3_cf_w_2_400_s_1_200=8.20e-11
+  mcm5m4m3_ca_w_2_400_s_2_100=3.06e-04 mcm5m4m3_cc_w_2_400_s_2_100=1.55e-12 mcm5m4m3_cf_w_2_400_s_2_100=9.16e-11
+  mcm5m4m3_ca_w_2_400_s_3_300=3.06e-04 mcm5m4m3_cc_w_2_400_s_3_300=2.00e-13 mcm5m4m3_cf_w_2_400_s_3_300=9.27e-11
+  mcm5m4m3_ca_w_2_400_s_9_000=3.06e-04 mcm5m4m3_cc_w_2_400_s_9_000=5.00e-14 mcm5m4m3_cf_w_2_400_s_9_000=9.32e-11
+  mcrdlm4f_ca_w_0_300_s_0_300=1.67e-05 mcrdlm4f_cc_w_0_300_s_0_300=1.25e-10 mcrdlm4f_cf_w_0_300_s_0_300=2.08e-12
+  mcrdlm4f_ca_w_0_300_s_0_360=1.67e-05 mcrdlm4f_cc_w_0_300_s_0_360=1.16e-10 mcrdlm4f_cf_w_0_300_s_0_360=2.58e-12
+  mcrdlm4f_ca_w_0_300_s_0_450=1.67e-05 mcrdlm4f_cc_w_0_300_s_0_450=1.03e-10 mcrdlm4f_cf_w_0_300_s_0_450=3.34e-12
+  mcrdlm4f_ca_w_0_300_s_0_600=1.67e-05 mcrdlm4f_cc_w_0_300_s_0_600=8.80e-11 mcrdlm4f_cf_w_0_300_s_0_600=4.59e-12
+  mcrdlm4f_ca_w_0_300_s_0_800=1.67e-05 mcrdlm4f_cc_w_0_300_s_0_800=7.32e-11 mcrdlm4f_cf_w_0_300_s_0_800=6.07e-12
+  mcrdlm4f_ca_w_0_300_s_1_000=1.67e-05 mcrdlm4f_cc_w_0_300_s_1_000=6.24e-11 mcrdlm4f_cf_w_0_300_s_1_000=7.60e-12
+  mcrdlm4f_ca_w_0_300_s_1_200=1.67e-05 mcrdlm4f_cc_w_0_300_s_1_200=5.41e-11 mcrdlm4f_cf_w_0_300_s_1_200=9.08e-12
+  mcrdlm4f_ca_w_0_300_s_2_100=1.67e-05 mcrdlm4f_cc_w_0_300_s_2_100=3.35e-11 mcrdlm4f_cf_w_0_300_s_2_100=1.54e-11
+  mcrdlm4f_ca_w_0_300_s_3_300=1.67e-05 mcrdlm4f_cc_w_0_300_s_3_300=2.07e-11 mcrdlm4f_cf_w_0_300_s_3_300=2.16e-11
+  mcrdlm4f_ca_w_0_300_s_9_000=1.67e-05 mcrdlm4f_cc_w_0_300_s_9_000=3.08e-12 mcrdlm4f_cf_w_0_300_s_9_000=3.49e-11
+  mcrdlm4f_ca_w_2_400_s_0_300=1.67e-05 mcrdlm4f_cc_w_2_400_s_0_300=1.50e-10 mcrdlm4f_cf_w_2_400_s_0_300=2.11e-12
+  mcrdlm4f_ca_w_2_400_s_0_360=1.67e-05 mcrdlm4f_cc_w_2_400_s_0_360=1.39e-10 mcrdlm4f_cf_w_2_400_s_0_360=2.60e-12
+  mcrdlm4f_ca_w_2_400_s_0_450=1.67e-05 mcrdlm4f_cc_w_2_400_s_0_450=1.25e-10 mcrdlm4f_cf_w_2_400_s_0_450=3.33e-12
+  mcrdlm4f_ca_w_2_400_s_0_600=1.67e-05 mcrdlm4f_cc_w_2_400_s_0_600=1.06e-10 mcrdlm4f_cf_w_2_400_s_0_600=4.54e-12
+  mcrdlm4f_ca_w_2_400_s_0_800=1.67e-05 mcrdlm4f_cc_w_2_400_s_0_800=8.85e-11 mcrdlm4f_cf_w_2_400_s_0_800=6.12e-12
+  mcrdlm4f_ca_w_2_400_s_1_000=1.67e-05 mcrdlm4f_cc_w_2_400_s_1_000=7.55e-11 mcrdlm4f_cf_w_2_400_s_1_000=7.67e-12
+  mcrdlm4f_ca_w_2_400_s_1_200=1.67e-05 mcrdlm4f_cc_w_2_400_s_1_200=6.57e-11 mcrdlm4f_cf_w_2_400_s_1_200=9.18e-12
+  mcrdlm4f_ca_w_2_400_s_2_100=1.67e-05 mcrdlm4f_cc_w_2_400_s_2_100=4.09e-11 mcrdlm4f_cf_w_2_400_s_2_100=1.55e-11
+  mcrdlm4f_ca_w_2_400_s_3_300=1.67e-05 mcrdlm4f_cc_w_2_400_s_3_300=2.53e-11 mcrdlm4f_cf_w_2_400_s_3_300=2.24e-11
+  mcrdlm4f_ca_w_2_400_s_9_000=1.67e-05 mcrdlm4f_cc_w_2_400_s_9_000=3.92e-12 mcrdlm4f_cf_w_2_400_s_9_000=3.80e-11
+  mcrdlm4d_ca_w_0_300_s_0_300=1.74e-05 mcrdlm4d_cc_w_0_300_s_0_300=1.25e-10 mcrdlm4d_cf_w_0_300_s_0_300=2.17e-12
+  mcrdlm4d_ca_w_0_300_s_0_360=1.74e-05 mcrdlm4d_cc_w_0_300_s_0_360=1.16e-10 mcrdlm4d_cf_w_0_300_s_0_360=2.69e-12
+  mcrdlm4d_ca_w_0_300_s_0_450=1.74e-05 mcrdlm4d_cc_w_0_300_s_0_450=1.03e-10 mcrdlm4d_cf_w_0_300_s_0_450=3.48e-12
+  mcrdlm4d_ca_w_0_300_s_0_600=1.74e-05 mcrdlm4d_cc_w_0_300_s_0_600=8.77e-11 mcrdlm4d_cf_w_0_300_s_0_600=4.78e-12
+  mcrdlm4d_ca_w_0_300_s_0_800=1.74e-05 mcrdlm4d_cc_w_0_300_s_0_800=7.29e-11 mcrdlm4d_cf_w_0_300_s_0_800=6.32e-12
+  mcrdlm4d_ca_w_0_300_s_1_000=1.74e-05 mcrdlm4d_cc_w_0_300_s_1_000=6.21e-11 mcrdlm4d_cf_w_0_300_s_1_000=7.92e-12
+  mcrdlm4d_ca_w_0_300_s_1_200=1.74e-05 mcrdlm4d_cc_w_0_300_s_1_200=5.38e-11 mcrdlm4d_cf_w_0_300_s_1_200=9.46e-12
+  mcrdlm4d_ca_w_0_300_s_2_100=1.74e-05 mcrdlm4d_cc_w_0_300_s_2_100=3.30e-11 mcrdlm4d_cf_w_0_300_s_2_100=1.59e-11
+  mcrdlm4d_ca_w_0_300_s_3_300=1.74e-05 mcrdlm4d_cc_w_0_300_s_3_300=2.02e-11 mcrdlm4d_cf_w_0_300_s_3_300=2.24e-11
+  mcrdlm4d_ca_w_0_300_s_9_000=1.74e-05 mcrdlm4d_cc_w_0_300_s_9_000=2.90e-12 mcrdlm4d_cf_w_0_300_s_9_000=3.55e-11
+  mcrdlm4d_ca_w_2_400_s_0_300=1.74e-05 mcrdlm4d_cc_w_2_400_s_0_300=1.49e-10 mcrdlm4d_cf_w_2_400_s_0_300=2.20e-12
+  mcrdlm4d_ca_w_2_400_s_0_360=1.74e-05 mcrdlm4d_cc_w_2_400_s_0_360=1.38e-10 mcrdlm4d_cf_w_2_400_s_0_360=2.71e-12
+  mcrdlm4d_ca_w_2_400_s_0_450=1.74e-05 mcrdlm4d_cc_w_2_400_s_0_450=1.24e-10 mcrdlm4d_cf_w_2_400_s_0_450=3.48e-12
+  mcrdlm4d_ca_w_2_400_s_0_600=1.74e-05 mcrdlm4d_cc_w_2_400_s_0_600=1.06e-10 mcrdlm4d_cf_w_2_400_s_0_600=4.74e-12
+  mcrdlm4d_ca_w_2_400_s_0_800=1.74e-05 mcrdlm4d_cc_w_2_400_s_0_800=8.79e-11 mcrdlm4d_cf_w_2_400_s_0_800=6.38e-12
+  mcrdlm4d_ca_w_2_400_s_1_000=1.74e-05 mcrdlm4d_cc_w_2_400_s_1_000=7.49e-11 mcrdlm4d_cf_w_2_400_s_1_000=8.00e-12
+  mcrdlm4d_ca_w_2_400_s_1_200=1.74e-05 mcrdlm4d_cc_w_2_400_s_1_200=6.50e-11 mcrdlm4d_cf_w_2_400_s_1_200=9.56e-12
+  mcrdlm4d_ca_w_2_400_s_2_100=1.74e-05 mcrdlm4d_cc_w_2_400_s_2_100=4.02e-11 mcrdlm4d_cf_w_2_400_s_2_100=1.60e-11
+  mcrdlm4d_ca_w_2_400_s_3_300=1.74e-05 mcrdlm4d_cc_w_2_400_s_3_300=2.47e-11 mcrdlm4d_cf_w_2_400_s_3_300=2.31e-11
+  mcrdlm4d_ca_w_2_400_s_9_000=1.74e-05 mcrdlm4d_cc_w_2_400_s_9_000=3.67e-12 mcrdlm4d_cf_w_2_400_s_9_000=3.87e-11
+  mcrdlm4p1_ca_w_0_300_s_0_300=1.87e-05 mcrdlm4p1_cc_w_0_300_s_0_300=1.25e-10 mcrdlm4p1_cf_w_0_300_s_0_300=2.33e-12
+  mcrdlm4p1_ca_w_0_300_s_0_360=1.87e-05 mcrdlm4p1_cc_w_0_300_s_0_360=1.15e-10 mcrdlm4p1_cf_w_0_300_s_0_360=2.88e-12
+  mcrdlm4p1_ca_w_0_300_s_0_450=1.87e-05 mcrdlm4p1_cc_w_0_300_s_0_450=1.03e-10 mcrdlm4p1_cf_w_0_300_s_0_450=3.73e-12
+  mcrdlm4p1_ca_w_0_300_s_0_600=1.87e-05 mcrdlm4p1_cc_w_0_300_s_0_600=8.72e-11 mcrdlm4p1_cf_w_0_300_s_0_600=5.11e-12
+  mcrdlm4p1_ca_w_0_300_s_0_800=1.87e-05 mcrdlm4p1_cc_w_0_300_s_0_800=7.23e-11 mcrdlm4p1_cf_w_0_300_s_0_800=6.75e-12
+  mcrdlm4p1_ca_w_0_300_s_1_000=1.87e-05 mcrdlm4p1_cc_w_0_300_s_1_000=6.13e-11 mcrdlm4p1_cf_w_0_300_s_1_000=8.45e-12
+  mcrdlm4p1_ca_w_0_300_s_1_200=1.87e-05 mcrdlm4p1_cc_w_0_300_s_1_200=5.30e-11 mcrdlm4p1_cf_w_0_300_s_1_200=1.01e-11
+  mcrdlm4p1_ca_w_0_300_s_2_100=1.87e-05 mcrdlm4p1_cc_w_0_300_s_2_100=3.23e-11 mcrdlm4p1_cf_w_0_300_s_2_100=1.69e-11
+  mcrdlm4p1_ca_w_0_300_s_3_300=1.87e-05 mcrdlm4p1_cc_w_0_300_s_3_300=1.95e-11 mcrdlm4p1_cf_w_0_300_s_3_300=2.36e-11
+  mcrdlm4p1_ca_w_0_300_s_9_000=1.87e-05 mcrdlm4p1_cc_w_0_300_s_9_000=2.61e-12 mcrdlm4p1_cf_w_0_300_s_9_000=3.66e-11
+  mcrdlm4p1_ca_w_2_400_s_0_300=1.87e-05 mcrdlm4p1_cc_w_2_400_s_0_300=1.48e-10 mcrdlm4p1_cf_w_2_400_s_0_300=2.37e-12
+  mcrdlm4p1_ca_w_2_400_s_0_360=1.87e-05 mcrdlm4p1_cc_w_2_400_s_0_360=1.37e-10 mcrdlm4p1_cf_w_2_400_s_0_360=2.92e-12
+  mcrdlm4p1_ca_w_2_400_s_0_450=1.87e-05 mcrdlm4p1_cc_w_2_400_s_0_450=1.23e-10 mcrdlm4p1_cf_w_2_400_s_0_450=3.73e-12
+  mcrdlm4p1_ca_w_2_400_s_0_600=1.87e-05 mcrdlm4p1_cc_w_2_400_s_0_600=1.04e-10 mcrdlm4p1_cf_w_2_400_s_0_600=5.08e-12
+  mcrdlm4p1_ca_w_2_400_s_0_800=1.87e-05 mcrdlm4p1_cc_w_2_400_s_0_800=8.67e-11 mcrdlm4p1_cf_w_2_400_s_0_800=6.82e-12
+  mcrdlm4p1_ca_w_2_400_s_1_000=1.87e-05 mcrdlm4p1_cc_w_2_400_s_1_000=7.39e-11 mcrdlm4p1_cf_w_2_400_s_1_000=8.54e-12
+  mcrdlm4p1_ca_w_2_400_s_1_200=1.87e-05 mcrdlm4p1_cc_w_2_400_s_1_200=6.40e-11 mcrdlm4p1_cf_w_2_400_s_1_200=1.02e-11
+  mcrdlm4p1_ca_w_2_400_s_2_100=1.87e-05 mcrdlm4p1_cc_w_2_400_s_2_100=3.92e-11 mcrdlm4p1_cf_w_2_400_s_2_100=1.70e-11
+  mcrdlm4p1_ca_w_2_400_s_3_300=1.87e-05 mcrdlm4p1_cc_w_2_400_s_3_300=2.37e-11 mcrdlm4p1_cf_w_2_400_s_3_300=2.44e-11
+  mcrdlm4p1_ca_w_2_400_s_9_000=1.87e-05 mcrdlm4p1_cc_w_2_400_s_9_000=3.30e-12 mcrdlm4p1_cf_w_2_400_s_9_000=3.98e-11
+  mcrdlm4l1_ca_w_0_300_s_0_300=2.03e-05 mcrdlm4l1_cc_w_0_300_s_0_300=1.25e-10 mcrdlm4l1_cf_w_0_300_s_0_300=2.52e-12
+  mcrdlm4l1_ca_w_0_300_s_0_360=2.03e-05 mcrdlm4l1_cc_w_0_300_s_0_360=1.15e-10 mcrdlm4l1_cf_w_0_300_s_0_360=3.12e-12
+  mcrdlm4l1_ca_w_0_300_s_0_450=2.03e-05 mcrdlm4l1_cc_w_0_300_s_0_450=1.02e-10 mcrdlm4l1_cf_w_0_300_s_0_450=4.03e-12
+  mcrdlm4l1_ca_w_0_300_s_0_600=2.03e-05 mcrdlm4l1_cc_w_0_300_s_0_600=8.67e-11 mcrdlm4l1_cf_w_0_300_s_0_600=5.51e-12
+  mcrdlm4l1_ca_w_0_300_s_0_800=2.03e-05 mcrdlm4l1_cc_w_0_300_s_0_800=7.17e-11 mcrdlm4l1_cf_w_0_300_s_0_800=7.29e-12
+  mcrdlm4l1_ca_w_0_300_s_1_000=2.03e-05 mcrdlm4l1_cc_w_0_300_s_1_000=6.06e-11 mcrdlm4l1_cf_w_0_300_s_1_000=9.12e-12
+  mcrdlm4l1_ca_w_0_300_s_1_200=2.03e-05 mcrdlm4l1_cc_w_0_300_s_1_200=5.23e-11 mcrdlm4l1_cf_w_0_300_s_1_200=1.09e-11
+  mcrdlm4l1_ca_w_0_300_s_2_100=2.03e-05 mcrdlm4l1_cc_w_0_300_s_2_100=3.14e-11 mcrdlm4l1_cf_w_0_300_s_2_100=1.80e-11
+  mcrdlm4l1_ca_w_0_300_s_3_300=2.03e-05 mcrdlm4l1_cc_w_0_300_s_3_300=1.86e-11 mcrdlm4l1_cf_w_0_300_s_3_300=2.50e-11
+  mcrdlm4l1_ca_w_0_300_s_9_000=2.03e-05 mcrdlm4l1_cc_w_0_300_s_9_000=2.31e-12 mcrdlm4l1_cf_w_0_300_s_9_000=3.79e-11
+  mcrdlm4l1_ca_w_2_400_s_0_300=2.03e-05 mcrdlm4l1_cc_w_2_400_s_0_300=1.47e-10 mcrdlm4l1_cf_w_2_400_s_0_300=2.54e-12
+  mcrdlm4l1_ca_w_2_400_s_0_360=2.03e-05 mcrdlm4l1_cc_w_2_400_s_0_360=1.36e-10 mcrdlm4l1_cf_w_2_400_s_0_360=3.13e-12
+  mcrdlm4l1_ca_w_2_400_s_0_450=2.03e-05 mcrdlm4l1_cc_w_2_400_s_0_450=1.22e-10 mcrdlm4l1_cf_w_2_400_s_0_450=4.01e-12
+  mcrdlm4l1_ca_w_2_400_s_0_600=2.03e-05 mcrdlm4l1_cc_w_2_400_s_0_600=1.04e-10 mcrdlm4l1_cf_w_2_400_s_0_600=5.45e-12
+  mcrdlm4l1_ca_w_2_400_s_0_800=2.03e-05 mcrdlm4l1_cc_w_2_400_s_0_800=8.56e-11 mcrdlm4l1_cf_w_2_400_s_0_800=7.34e-12
+  mcrdlm4l1_ca_w_2_400_s_1_000=2.03e-05 mcrdlm4l1_cc_w_2_400_s_1_000=7.27e-11 mcrdlm4l1_cf_w_2_400_s_1_000=9.19e-12
+  mcrdlm4l1_ca_w_2_400_s_1_200=2.03e-05 mcrdlm4l1_cc_w_2_400_s_1_200=6.27e-11 mcrdlm4l1_cf_w_2_400_s_1_200=1.10e-11
+  mcrdlm4l1_ca_w_2_400_s_2_100=2.03e-05 mcrdlm4l1_cc_w_2_400_s_2_100=3.81e-11 mcrdlm4l1_cf_w_2_400_s_2_100=1.82e-11
+  mcrdlm4l1_ca_w_2_400_s_3_300=2.03e-05 mcrdlm4l1_cc_w_2_400_s_3_300=2.26e-11 mcrdlm4l1_cf_w_2_400_s_3_300=2.58e-11
+  mcrdlm4l1_ca_w_2_400_s_9_000=2.03e-05 mcrdlm4l1_cc_w_2_400_s_9_000=2.94e-12 mcrdlm4l1_cf_w_2_400_s_9_000=4.10e-11
+  mcrdlm4m1_ca_w_0_300_s_0_300=2.45e-05 mcrdlm4m1_cc_w_0_300_s_0_300=1.24e-10 mcrdlm4m1_cf_w_0_300_s_0_300=3.02e-12
+  mcrdlm4m1_ca_w_0_300_s_0_360=2.45e-05 mcrdlm4m1_cc_w_0_300_s_0_360=1.14e-10 mcrdlm4m1_cf_w_0_300_s_0_360=3.74e-12
+  mcrdlm4m1_ca_w_0_300_s_0_450=2.45e-05 mcrdlm4m1_cc_w_0_300_s_0_450=1.01e-10 mcrdlm4m1_cf_w_0_300_s_0_450=4.82e-12
+  mcrdlm4m1_ca_w_0_300_s_0_600=2.45e-05 mcrdlm4m1_cc_w_0_300_s_0_600=8.53e-11 mcrdlm4m1_cf_w_0_300_s_0_600=6.57e-12
+  mcrdlm4m1_ca_w_0_300_s_0_800=2.45e-05 mcrdlm4m1_cc_w_0_300_s_0_800=7.01e-11 mcrdlm4m1_cf_w_0_300_s_0_800=8.69e-12
+  mcrdlm4m1_ca_w_0_300_s_1_000=2.45e-05 mcrdlm4m1_cc_w_0_300_s_1_000=5.89e-11 mcrdlm4m1_cf_w_0_300_s_1_000=1.08e-11
+  mcrdlm4m1_ca_w_0_300_s_1_200=2.45e-05 mcrdlm4m1_cc_w_0_300_s_1_200=5.04e-11 mcrdlm4m1_cf_w_0_300_s_1_200=1.29e-11
+  mcrdlm4m1_ca_w_0_300_s_2_100=2.45e-05 mcrdlm4m1_cc_w_0_300_s_2_100=2.94e-11 mcrdlm4m1_cf_w_0_300_s_2_100=2.10e-11
+  mcrdlm4m1_ca_w_0_300_s_3_300=2.45e-05 mcrdlm4m1_cc_w_0_300_s_3_300=1.67e-11 mcrdlm4m1_cf_w_0_300_s_3_300=2.84e-11
+  mcrdlm4m1_ca_w_0_300_s_9_000=2.45e-05 mcrdlm4m1_cc_w_0_300_s_9_000=1.78e-12 mcrdlm4m1_cf_w_0_300_s_9_000=4.07e-11
+  mcrdlm4m1_ca_w_2_400_s_0_300=2.45e-05 mcrdlm4m1_cc_w_2_400_s_0_300=1.44e-10 mcrdlm4m1_cf_w_2_400_s_0_300=3.03e-12
+  mcrdlm4m1_ca_w_2_400_s_0_360=2.45e-05 mcrdlm4m1_cc_w_2_400_s_0_360=1.34e-10 mcrdlm4m1_cf_w_2_400_s_0_360=3.74e-12
+  mcrdlm4m1_ca_w_2_400_s_0_450=2.45e-05 mcrdlm4m1_cc_w_2_400_s_0_450=1.19e-10 mcrdlm4m1_cf_w_2_400_s_0_450=4.79e-12
+  mcrdlm4m1_ca_w_2_400_s_0_600=2.45e-05 mcrdlm4m1_cc_w_2_400_s_0_600=1.01e-10 mcrdlm4m1_cf_w_2_400_s_0_600=6.51e-12
+  mcrdlm4m1_ca_w_2_400_s_0_800=2.45e-05 mcrdlm4m1_cc_w_2_400_s_0_800=8.30e-11 mcrdlm4m1_cf_w_2_400_s_0_800=8.74e-12
+  mcrdlm4m1_ca_w_2_400_s_1_000=2.45e-05 mcrdlm4m1_cc_w_2_400_s_1_000=7.00e-11 mcrdlm4m1_cf_w_2_400_s_1_000=1.09e-11
+  mcrdlm4m1_ca_w_2_400_s_1_200=2.45e-05 mcrdlm4m1_cc_w_2_400_s_1_200=6.01e-11 mcrdlm4m1_cf_w_2_400_s_1_200=1.30e-11
+  mcrdlm4m1_ca_w_2_400_s_2_100=2.45e-05 mcrdlm4m1_cc_w_2_400_s_2_100=3.55e-11 mcrdlm4m1_cf_w_2_400_s_2_100=2.12e-11
+  mcrdlm4m1_ca_w_2_400_s_3_300=2.45e-05 mcrdlm4m1_cc_w_2_400_s_3_300=2.05e-11 mcrdlm4m1_cf_w_2_400_s_3_300=2.94e-11
+  mcrdlm4m1_ca_w_2_400_s_9_000=2.45e-05 mcrdlm4m1_cc_w_2_400_s_9_000=2.33e-12 mcrdlm4m1_cf_w_2_400_s_9_000=4.40e-11
+  mcrdlm4m2_ca_w_0_300_s_0_300=3.12e-05 mcrdlm4m2_cc_w_0_300_s_0_300=1.22e-10 mcrdlm4m2_cf_w_0_300_s_0_300=3.84e-12
+  mcrdlm4m2_ca_w_0_300_s_0_360=3.12e-05 mcrdlm4m2_cc_w_0_300_s_0_360=1.12e-10 mcrdlm4m2_cf_w_0_300_s_0_360=4.73e-12
+  mcrdlm4m2_ca_w_0_300_s_0_450=3.12e-05 mcrdlm4m2_cc_w_0_300_s_0_450=9.96e-11 mcrdlm4m2_cf_w_0_300_s_0_450=6.09e-12
+  mcrdlm4m2_ca_w_0_300_s_0_600=3.12e-05 mcrdlm4m2_cc_w_0_300_s_0_600=8.32e-11 mcrdlm4m2_cf_w_0_300_s_0_600=8.24e-12
+  mcrdlm4m2_ca_w_0_300_s_0_800=3.12e-05 mcrdlm4m2_cc_w_0_300_s_0_800=6.79e-11 mcrdlm4m2_cf_w_0_300_s_0_800=1.09e-11
+  mcrdlm4m2_ca_w_0_300_s_1_000=3.12e-05 mcrdlm4m2_cc_w_0_300_s_1_000=5.65e-11 mcrdlm4m2_cf_w_0_300_s_1_000=1.35e-11
+  mcrdlm4m2_ca_w_0_300_s_1_200=3.12e-05 mcrdlm4m2_cc_w_0_300_s_1_200=4.81e-11 mcrdlm4m2_cf_w_0_300_s_1_200=1.59e-11
+  mcrdlm4m2_ca_w_0_300_s_2_100=3.12e-05 mcrdlm4m2_cc_w_0_300_s_2_100=2.68e-11 mcrdlm4m2_cf_w_0_300_s_2_100=2.52e-11
+  mcrdlm4m2_ca_w_0_300_s_3_300=3.12e-05 mcrdlm4m2_cc_w_0_300_s_3_300=1.45e-11 mcrdlm4m2_cf_w_0_300_s_3_300=3.31e-11
+  mcrdlm4m2_ca_w_0_300_s_9_000=3.12e-05 mcrdlm4m2_cc_w_0_300_s_9_000=1.29e-12 mcrdlm4m2_cf_w_0_300_s_9_000=4.45e-11
+  mcrdlm4m2_ca_w_2_400_s_0_300=3.12e-05 mcrdlm4m2_cc_w_2_400_s_0_300=1.41e-10 mcrdlm4m2_cf_w_2_400_s_0_300=3.85e-12
+  mcrdlm4m2_ca_w_2_400_s_0_360=3.12e-05 mcrdlm4m2_cc_w_2_400_s_0_360=1.30e-10 mcrdlm4m2_cf_w_2_400_s_0_360=4.74e-12
+  mcrdlm4m2_ca_w_2_400_s_0_450=3.12e-05 mcrdlm4m2_cc_w_2_400_s_0_450=1.16e-10 mcrdlm4m2_cf_w_2_400_s_0_450=6.05e-12
+  mcrdlm4m2_ca_w_2_400_s_0_600=3.12e-05 mcrdlm4m2_cc_w_2_400_s_0_600=9.74e-11 mcrdlm4m2_cf_w_2_400_s_0_600=8.19e-12
+  mcrdlm4m2_ca_w_2_400_s_0_800=3.12e-05 mcrdlm4m2_cc_w_2_400_s_0_800=7.97e-11 mcrdlm4m2_cf_w_2_400_s_0_800=1.09e-11
+  mcrdlm4m2_ca_w_2_400_s_1_000=3.12e-05 mcrdlm4m2_cc_w_2_400_s_1_000=6.67e-11 mcrdlm4m2_cf_w_2_400_s_1_000=1.36e-11
+  mcrdlm4m2_ca_w_2_400_s_1_200=3.12e-05 mcrdlm4m2_cc_w_2_400_s_1_200=5.68e-11 mcrdlm4m2_cf_w_2_400_s_1_200=1.60e-11
+  mcrdlm4m2_ca_w_2_400_s_2_100=3.12e-05 mcrdlm4m2_cc_w_2_400_s_2_100=3.25e-11 mcrdlm4m2_cf_w_2_400_s_2_100=2.54e-11
+  mcrdlm4m2_ca_w_2_400_s_3_300=3.12e-05 mcrdlm4m2_cc_w_2_400_s_3_300=1.81e-11 mcrdlm4m2_cf_w_2_400_s_3_300=3.43e-11
+  mcrdlm4m2_ca_w_2_400_s_9_000=3.12e-05 mcrdlm4m2_cc_w_2_400_s_9_000=1.71e-12 mcrdlm4m2_cf_w_2_400_s_9_000=4.79e-11
+  mcrdlm4m3_ca_w_0_300_s_0_300=1.97e-04 mcrdlm4m3_cc_w_0_300_s_0_300=1.04e-10 mcrdlm4m3_cf_w_0_300_s_0_300=2.04e-11
+  mcrdlm4m3_ca_w_0_300_s_0_360=1.97e-04 mcrdlm4m3_cc_w_0_300_s_0_360=9.37e-11 mcrdlm4m3_cf_w_0_300_s_0_360=2.41e-11
+  mcrdlm4m3_ca_w_0_300_s_0_450=1.97e-04 mcrdlm4m3_cc_w_0_300_s_0_450=8.13e-11 mcrdlm4m3_cf_w_0_300_s_0_450=2.91e-11
+  mcrdlm4m3_ca_w_0_300_s_0_600=1.97e-04 mcrdlm4m3_cc_w_0_300_s_0_600=6.53e-11 mcrdlm4m3_cf_w_0_300_s_0_600=3.59e-11
+  mcrdlm4m3_ca_w_0_300_s_0_800=1.97e-04 mcrdlm4m3_cc_w_0_300_s_0_800=5.09e-11 mcrdlm4m3_cf_w_0_300_s_0_800=4.29e-11
+  mcrdlm4m3_ca_w_0_300_s_1_000=1.97e-04 mcrdlm4m3_cc_w_0_300_s_1_000=4.01e-11 mcrdlm4m3_cf_w_0_300_s_1_000=4.85e-11
+  mcrdlm4m3_ca_w_0_300_s_1_200=1.97e-04 mcrdlm4m3_cc_w_0_300_s_1_200=3.25e-11 mcrdlm4m3_cf_w_0_300_s_1_200=5.28e-11
+  mcrdlm4m3_ca_w_0_300_s_2_100=1.97e-04 mcrdlm4m3_cc_w_0_300_s_2_100=1.51e-11 mcrdlm4m3_cf_w_0_300_s_2_100=6.54e-11
+  mcrdlm4m3_ca_w_0_300_s_3_300=1.97e-04 mcrdlm4m3_cc_w_0_300_s_3_300=6.91e-12 mcrdlm4m3_cf_w_0_300_s_3_300=7.27e-11
+  mcrdlm4m3_ca_w_0_300_s_9_000=1.97e-04 mcrdlm4m3_cc_w_0_300_s_9_000=4.20e-13 mcrdlm4m3_cf_w_0_300_s_9_000=7.89e-11
+  mcrdlm4m3_ca_w_2_400_s_0_300=1.97e-04 mcrdlm4m3_cc_w_2_400_s_0_300=1.20e-10 mcrdlm4m3_cf_w_2_400_s_0_300=2.04e-11
+  mcrdlm4m3_ca_w_2_400_s_0_360=1.97e-04 mcrdlm4m3_cc_w_2_400_s_0_360=1.09e-10 mcrdlm4m3_cf_w_2_400_s_0_360=2.41e-11
+  mcrdlm4m3_ca_w_2_400_s_0_450=1.97e-04 mcrdlm4m3_cc_w_2_400_s_0_450=9.51e-11 mcrdlm4m3_cf_w_2_400_s_0_450=2.91e-11
+  mcrdlm4m3_ca_w_2_400_s_0_600=1.97e-04 mcrdlm4m3_cc_w_2_400_s_0_600=7.79e-11 mcrdlm4m3_cf_w_2_400_s_0_600=3.58e-11
+  mcrdlm4m3_ca_w_2_400_s_0_800=1.97e-04 mcrdlm4m3_cc_w_2_400_s_0_800=6.13e-11 mcrdlm4m3_cf_w_2_400_s_0_800=4.29e-11
+  mcrdlm4m3_ca_w_2_400_s_1_000=1.97e-04 mcrdlm4m3_cc_w_2_400_s_1_000=4.95e-11 mcrdlm4m3_cf_w_2_400_s_1_000=4.86e-11
+  mcrdlm4m3_ca_w_2_400_s_1_200=1.97e-04 mcrdlm4m3_cc_w_2_400_s_1_200=4.07e-11 mcrdlm4m3_cf_w_2_400_s_1_200=5.30e-11
+  mcrdlm4m3_ca_w_2_400_s_2_100=1.97e-04 mcrdlm4m3_cc_w_2_400_s_2_100=2.07e-11 mcrdlm4m3_cf_w_2_400_s_2_100=6.62e-11
+  mcrdlm4m3_ca_w_2_400_s_3_300=1.97e-04 mcrdlm4m3_cc_w_2_400_s_3_300=1.01e-11 mcrdlm4m3_cf_w_2_400_s_3_300=7.50e-11
+  mcrdlm4m3_ca_w_2_400_s_9_000=1.97e-04 mcrdlm4m3_cc_w_2_400_s_9_000=5.80e-13 mcrdlm4m3_cf_w_2_400_s_9_000=8.40e-11
+  mcrdlm5f_ca_w_1_600_s_1_600=1.66e-05 mcrdlm5f_cc_w_1_600_s_1_600=7.83e-11 mcrdlm5f_cf_w_1_600_s_1_600=1.17e-11
+  mcrdlm5f_ca_w_1_600_s_1_700=1.66e-05 mcrdlm5f_cc_w_1_600_s_1_700=7.31e-11 mcrdlm5f_cf_w_1_600_s_1_700=1.25e-11
+  mcrdlm5f_ca_w_1_600_s_1_900=1.66e-05 mcrdlm5f_cc_w_1_600_s_1_900=6.45e-11 mcrdlm5f_cf_w_1_600_s_1_900=1.39e-11
+  mcrdlm5f_ca_w_1_600_s_2_000=1.66e-05 mcrdlm5f_cc_w_1_600_s_2_000=6.10e-11 mcrdlm5f_cf_w_1_600_s_2_000=1.46e-11
+  mcrdlm5f_ca_w_1_600_s_2_400=1.66e-05 mcrdlm5f_cc_w_1_600_s_2_400=4.95e-11 mcrdlm5f_cf_w_1_600_s_2_400=1.74e-11
+  mcrdlm5f_ca_w_1_600_s_2_800=1.66e-05 mcrdlm5f_cc_w_1_600_s_2_800=4.13e-11 mcrdlm5f_cf_w_1_600_s_2_800=1.99e-11
+  mcrdlm5f_ca_w_1_600_s_3_200=1.66e-05 mcrdlm5f_cc_w_1_600_s_3_200=3.50e-11 mcrdlm5f_cf_w_1_600_s_3_200=2.24e-11
+  mcrdlm5f_ca_w_1_600_s_4_800=1.66e-05 mcrdlm5f_cc_w_1_600_s_4_800=1.95e-11 mcrdlm5f_cf_w_1_600_s_4_800=3.04e-11
+  mcrdlm5f_ca_w_1_600_s_10_000=1.66e-05 mcrdlm5f_cc_w_1_600_s_10_000=3.62e-12 mcrdlm5f_cf_w_1_600_s_10_000=4.27e-11
+  mcrdlm5f_ca_w_1_600_s_12_000=1.66e-05 mcrdlm5f_cc_w_1_600_s_12_000=1.93e-12 mcrdlm5f_cf_w_1_600_s_12_000=4.43e-11
+  mcrdlm5f_ca_w_4_000_s_1_600=1.66e-05 mcrdlm5f_cc_w_4_000_s_1_600=8.03e-11 mcrdlm5f_cf_w_4_000_s_1_600=1.18e-11
+  mcrdlm5f_ca_w_4_000_s_1_700=1.66e-05 mcrdlm5f_cc_w_4_000_s_1_700=7.50e-11 mcrdlm5f_cf_w_4_000_s_1_700=1.25e-11
+  mcrdlm5f_ca_w_4_000_s_1_900=1.66e-05 mcrdlm5f_cc_w_4_000_s_1_900=6.63e-11 mcrdlm5f_cf_w_4_000_s_1_900=1.39e-11
+  mcrdlm5f_ca_w_4_000_s_2_000=1.66e-05 mcrdlm5f_cc_w_4_000_s_2_000=6.25e-11 mcrdlm5f_cf_w_4_000_s_2_000=1.46e-11
+  mcrdlm5f_ca_w_4_000_s_2_400=1.66e-05 mcrdlm5f_cc_w_4_000_s_2_400=5.08e-11 mcrdlm5f_cf_w_4_000_s_2_400=1.74e-11
+  mcrdlm5f_ca_w_4_000_s_2_800=1.66e-05 mcrdlm5f_cc_w_4_000_s_2_800=4.24e-11 mcrdlm5f_cf_w_4_000_s_2_800=2.00e-11
+  mcrdlm5f_ca_w_4_000_s_3_200=1.66e-05 mcrdlm5f_cc_w_4_000_s_3_200=3.60e-11 mcrdlm5f_cf_w_4_000_s_3_200=2.24e-11
+  mcrdlm5f_ca_w_4_000_s_4_800=1.66e-05 mcrdlm5f_cc_w_4_000_s_4_800=2.00e-11 mcrdlm5f_cf_w_4_000_s_4_800=3.06e-11
+  mcrdlm5f_ca_w_4_000_s_10_000=1.66e-05 mcrdlm5f_cc_w_4_000_s_10_000=3.79e-12 mcrdlm5f_cf_w_4_000_s_10_000=4.32e-11
+  mcrdlm5f_ca_w_4_000_s_12_000=1.66e-05 mcrdlm5f_cc_w_4_000_s_12_000=2.04e-12 mcrdlm5f_cf_w_4_000_s_12_000=4.48e-11
+  mcrdlm5d_ca_w_1_600_s_1_600=1.70e-05 mcrdlm5d_cc_w_1_600_s_1_600=7.79e-11 mcrdlm5d_cf_w_1_600_s_1_600=1.20e-11
+  mcrdlm5d_ca_w_1_600_s_1_700=1.70e-05 mcrdlm5d_cc_w_1_600_s_1_700=7.27e-11 mcrdlm5d_cf_w_1_600_s_1_700=1.28e-11
+  mcrdlm5d_ca_w_1_600_s_1_900=1.70e-05 mcrdlm5d_cc_w_1_600_s_1_900=6.42e-11 mcrdlm5d_cf_w_1_600_s_1_900=1.42e-11
+  mcrdlm5d_ca_w_1_600_s_2_000=1.70e-05 mcrdlm5d_cc_w_1_600_s_2_000=6.06e-11 mcrdlm5d_cf_w_1_600_s_2_000=1.49e-11
+  mcrdlm5d_ca_w_1_600_s_2_400=1.70e-05 mcrdlm5d_cc_w_1_600_s_2_400=4.90e-11 mcrdlm5d_cf_w_1_600_s_2_400=1.77e-11
+  mcrdlm5d_ca_w_1_600_s_2_800=1.70e-05 mcrdlm5d_cc_w_1_600_s_2_800=4.08e-11 mcrdlm5d_cf_w_1_600_s_2_800=2.04e-11
+  mcrdlm5d_ca_w_1_600_s_3_200=1.70e-05 mcrdlm5d_cc_w_1_600_s_3_200=3.46e-11 mcrdlm5d_cf_w_1_600_s_3_200=2.28e-11
+  mcrdlm5d_ca_w_1_600_s_4_800=1.70e-05 mcrdlm5d_cc_w_1_600_s_4_800=1.91e-11 mcrdlm5d_cf_w_1_600_s_4_800=3.10e-11
+  mcrdlm5d_ca_w_1_600_s_10_000=1.70e-05 mcrdlm5d_cc_w_1_600_s_10_000=3.48e-12 mcrdlm5d_cf_w_1_600_s_10_000=4.32e-11
+  mcrdlm5d_ca_w_1_600_s_12_000=1.70e-05 mcrdlm5d_cc_w_1_600_s_12_000=1.81e-12 mcrdlm5d_cf_w_1_600_s_12_000=4.48e-11
+  mcrdlm5d_ca_w_4_000_s_1_600=1.70e-05 mcrdlm5d_cc_w_4_000_s_1_600=7.98e-11 mcrdlm5d_cf_w_4_000_s_1_600=1.20e-11
+  mcrdlm5d_ca_w_4_000_s_1_700=1.70e-05 mcrdlm5d_cc_w_4_000_s_1_700=7.45e-11 mcrdlm5d_cf_w_4_000_s_1_700=1.28e-11
+  mcrdlm5d_ca_w_4_000_s_1_900=1.70e-05 mcrdlm5d_cc_w_4_000_s_1_900=6.58e-11 mcrdlm5d_cf_w_4_000_s_1_900=1.42e-11
+  mcrdlm5d_ca_w_4_000_s_2_000=1.70e-05 mcrdlm5d_cc_w_4_000_s_2_000=6.21e-11 mcrdlm5d_cf_w_4_000_s_2_000=1.50e-11
+  mcrdlm5d_ca_w_4_000_s_2_400=1.70e-05 mcrdlm5d_cc_w_4_000_s_2_400=5.03e-11 mcrdlm5d_cf_w_4_000_s_2_400=1.77e-11
+  mcrdlm5d_ca_w_4_000_s_2_800=1.70e-05 mcrdlm5d_cc_w_4_000_s_2_800=4.20e-11 mcrdlm5d_cf_w_4_000_s_2_800=2.04e-11
+  mcrdlm5d_ca_w_4_000_s_3_200=1.70e-05 mcrdlm5d_cc_w_4_000_s_3_200=3.55e-11 mcrdlm5d_cf_w_4_000_s_3_200=2.29e-11
+  mcrdlm5d_ca_w_4_000_s_4_800=1.70e-05 mcrdlm5d_cc_w_4_000_s_4_800=1.96e-11 mcrdlm5d_cf_w_4_000_s_4_800=3.12e-11
+  mcrdlm5d_ca_w_4_000_s_10_000=1.70e-05 mcrdlm5d_cc_w_4_000_s_10_000=3.56e-12 mcrdlm5d_cf_w_4_000_s_10_000=4.37e-11
+  mcrdlm5d_ca_w_4_000_s_12_000=1.70e-05 mcrdlm5d_cc_w_4_000_s_12_000=1.88e-12 mcrdlm5d_cf_w_4_000_s_12_000=4.53e-11
+  mcrdlm5p1_ca_w_1_600_s_1_600=1.76e-05 mcrdlm5p1_cc_w_1_600_s_1_600=7.73e-11 mcrdlm5p1_cf_w_1_600_s_1_600=1.24e-11
+  mcrdlm5p1_ca_w_1_600_s_1_700=1.76e-05 mcrdlm5p1_cc_w_1_600_s_1_700=7.21e-11 mcrdlm5p1_cf_w_1_600_s_1_700=1.32e-11
+  mcrdlm5p1_ca_w_1_600_s_1_900=1.76e-05 mcrdlm5p1_cc_w_1_600_s_1_900=6.35e-11 mcrdlm5p1_cf_w_1_600_s_1_900=1.47e-11
+  mcrdlm5p1_ca_w_1_600_s_2_000=1.76e-05 mcrdlm5p1_cc_w_1_600_s_2_000=5.99e-11 mcrdlm5p1_cf_w_1_600_s_2_000=1.54e-11
+  mcrdlm5p1_ca_w_1_600_s_2_400=1.76e-05 mcrdlm5p1_cc_w_1_600_s_2_400=4.85e-11 mcrdlm5p1_cf_w_1_600_s_2_400=1.83e-11
+  mcrdlm5p1_ca_w_1_600_s_2_800=1.76e-05 mcrdlm5p1_cc_w_1_600_s_2_800=4.03e-11 mcrdlm5p1_cf_w_1_600_s_2_800=2.11e-11
+  mcrdlm5p1_ca_w_1_600_s_3_200=1.76e-05 mcrdlm5p1_cc_w_1_600_s_3_200=3.39e-11 mcrdlm5p1_cf_w_1_600_s_3_200=2.35e-11
+  mcrdlm5p1_ca_w_1_600_s_4_800=1.76e-05 mcrdlm5p1_cc_w_1_600_s_4_800=1.85e-11 mcrdlm5p1_cf_w_1_600_s_4_800=3.18e-11
+  mcrdlm5p1_ca_w_1_600_s_10_000=1.76e-05 mcrdlm5p1_cc_w_1_600_s_10_000=3.18e-12 mcrdlm5p1_cf_w_1_600_s_10_000=4.40e-11
+  mcrdlm5p1_ca_w_1_600_s_12_000=1.76e-05 mcrdlm5p1_cc_w_1_600_s_12_000=1.62e-12 mcrdlm5p1_cf_w_1_600_s_12_000=4.55e-11
+  mcrdlm5p1_ca_w_4_000_s_1_600=1.76e-05 mcrdlm5p1_cc_w_4_000_s_1_600=7.91e-11 mcrdlm5p1_cf_w_4_000_s_1_600=1.24e-11
+  mcrdlm5p1_ca_w_4_000_s_1_700=1.76e-05 mcrdlm5p1_cc_w_4_000_s_1_700=7.38e-11 mcrdlm5p1_cf_w_4_000_s_1_700=1.32e-11
+  mcrdlm5p1_ca_w_4_000_s_1_900=1.76e-05 mcrdlm5p1_cc_w_4_000_s_1_900=6.50e-11 mcrdlm5p1_cf_w_4_000_s_1_900=1.47e-11
+  mcrdlm5p1_ca_w_4_000_s_2_000=1.76e-05 mcrdlm5p1_cc_w_4_000_s_2_000=6.13e-11 mcrdlm5p1_cf_w_4_000_s_2_000=1.55e-11
+  mcrdlm5p1_ca_w_4_000_s_2_400=1.76e-05 mcrdlm5p1_cc_w_4_000_s_2_400=4.96e-11 mcrdlm5p1_cf_w_4_000_s_2_400=1.83e-11
+  mcrdlm5p1_ca_w_4_000_s_2_800=1.76e-05 mcrdlm5p1_cc_w_4_000_s_2_800=4.12e-11 mcrdlm5p1_cf_w_4_000_s_2_800=2.11e-11
+  mcrdlm5p1_ca_w_4_000_s_3_200=1.76e-05 mcrdlm5p1_cc_w_4_000_s_3_200=3.48e-11 mcrdlm5p1_cf_w_4_000_s_3_200=2.36e-11
+  mcrdlm5p1_ca_w_4_000_s_4_800=1.76e-05 mcrdlm5p1_cc_w_4_000_s_4_800=1.90e-11 mcrdlm5p1_cf_w_4_000_s_4_800=3.20e-11
+  mcrdlm5p1_ca_w_4_000_s_10_000=1.76e-05 mcrdlm5p1_cc_w_4_000_s_10_000=3.30e-12 mcrdlm5p1_cf_w_4_000_s_10_000=4.44e-11
+  mcrdlm5p1_ca_w_4_000_s_12_000=1.76e-05 mcrdlm5p1_cc_w_4_000_s_12_000=1.69e-12 mcrdlm5p1_cf_w_4_000_s_12_000=4.59e-11
+  mcrdlm5l1_ca_w_1_600_s_1_600=1.83e-05 mcrdlm5l1_cc_w_1_600_s_1_600=7.66e-11 mcrdlm5l1_cf_w_1_600_s_1_600=1.29e-11
+  mcrdlm5l1_ca_w_1_600_s_1_700=1.83e-05 mcrdlm5l1_cc_w_1_600_s_1_700=7.14e-11 mcrdlm5l1_cf_w_1_600_s_1_700=1.37e-11
+  mcrdlm5l1_ca_w_1_600_s_1_900=1.83e-05 mcrdlm5l1_cc_w_1_600_s_1_900=6.28e-11 mcrdlm5l1_cf_w_1_600_s_1_900=1.53e-11
+  mcrdlm5l1_ca_w_1_600_s_2_000=1.83e-05 mcrdlm5l1_cc_w_1_600_s_2_000=5.92e-11 mcrdlm5l1_cf_w_1_600_s_2_000=1.60e-11
+  mcrdlm5l1_ca_w_1_600_s_2_400=1.83e-05 mcrdlm5l1_cc_w_1_600_s_2_400=4.78e-11 mcrdlm5l1_cf_w_1_600_s_2_400=1.90e-11
+  mcrdlm5l1_ca_w_1_600_s_2_800=1.83e-05 mcrdlm5l1_cc_w_1_600_s_2_800=3.95e-11 mcrdlm5l1_cf_w_1_600_s_2_800=2.18e-11
+  mcrdlm5l1_ca_w_1_600_s_3_200=1.83e-05 mcrdlm5l1_cc_w_1_600_s_3_200=3.32e-11 mcrdlm5l1_cf_w_1_600_s_3_200=2.44e-11
+  mcrdlm5l1_ca_w_1_600_s_4_800=1.83e-05 mcrdlm5l1_cc_w_1_600_s_4_800=1.78e-11 mcrdlm5l1_cf_w_1_600_s_4_800=3.29e-11
+  mcrdlm5l1_ca_w_1_600_s_10_000=1.83e-05 mcrdlm5l1_cc_w_1_600_s_10_000=2.89e-12 mcrdlm5l1_cf_w_1_600_s_10_000=4.49e-11
+  mcrdlm5l1_ca_w_1_600_s_12_000=1.83e-05 mcrdlm5l1_cc_w_1_600_s_12_000=1.46e-12 mcrdlm5l1_cf_w_1_600_s_12_000=4.62e-11
+  mcrdlm5l1_ca_w_4_000_s_1_600=1.83e-05 mcrdlm5l1_cc_w_4_000_s_1_600=7.83e-11 mcrdlm5l1_cf_w_4_000_s_1_600=1.29e-11
+  mcrdlm5l1_ca_w_4_000_s_1_700=1.83e-05 mcrdlm5l1_cc_w_4_000_s_1_700=7.30e-11 mcrdlm5l1_cf_w_4_000_s_1_700=1.37e-11
+  mcrdlm5l1_ca_w_4_000_s_1_900=1.83e-05 mcrdlm5l1_cc_w_4_000_s_1_900=6.42e-11 mcrdlm5l1_cf_w_4_000_s_1_900=1.53e-11
+  mcrdlm5l1_ca_w_4_000_s_2_000=1.83e-05 mcrdlm5l1_cc_w_4_000_s_2_000=6.05e-11 mcrdlm5l1_cf_w_4_000_s_2_000=1.61e-11
+  mcrdlm5l1_ca_w_4_000_s_2_400=1.83e-05 mcrdlm5l1_cc_w_4_000_s_2_400=4.87e-11 mcrdlm5l1_cf_w_4_000_s_2_400=1.90e-11
+  mcrdlm5l1_ca_w_4_000_s_2_800=1.83e-05 mcrdlm5l1_cc_w_4_000_s_2_800=4.04e-11 mcrdlm5l1_cf_w_4_000_s_2_800=2.19e-11
+  mcrdlm5l1_ca_w_4_000_s_3_200=1.83e-05 mcrdlm5l1_cc_w_4_000_s_3_200=3.39e-11 mcrdlm5l1_cf_w_4_000_s_3_200=2.45e-11
+  mcrdlm5l1_ca_w_4_000_s_4_800=1.83e-05 mcrdlm5l1_cc_w_4_000_s_4_800=1.83e-11 mcrdlm5l1_cf_w_4_000_s_4_800=3.30e-11
+  mcrdlm5l1_ca_w_4_000_s_10_000=1.83e-05 mcrdlm5l1_cc_w_4_000_s_10_000=2.98e-12 mcrdlm5l1_cf_w_4_000_s_10_000=4.53e-11
+  mcrdlm5l1_ca_w_4_000_s_12_000=1.83e-05 mcrdlm5l1_cc_w_4_000_s_12_000=1.51e-12 mcrdlm5l1_cf_w_4_000_s_12_000=4.67e-11
+  mcrdlm5m1_ca_w_1_600_s_1_600=2.00e-05 mcrdlm5m1_cc_w_1_600_s_1_600=7.52e-11 mcrdlm5m1_cf_w_1_600_s_1_600=1.40e-11
+  mcrdlm5m1_ca_w_1_600_s_1_700=2.00e-05 mcrdlm5m1_cc_w_1_600_s_1_700=6.99e-11 mcrdlm5m1_cf_w_1_600_s_1_700=1.49e-11
+  mcrdlm5m1_ca_w_1_600_s_1_900=2.00e-05 mcrdlm5m1_cc_w_1_600_s_1_900=6.13e-11 mcrdlm5m1_cf_w_1_600_s_1_900=1.66e-11
+  mcrdlm5m1_ca_w_1_600_s_2_000=2.00e-05 mcrdlm5m1_cc_w_1_600_s_2_000=5.77e-11 mcrdlm5m1_cf_w_1_600_s_2_000=1.74e-11
+  mcrdlm5m1_ca_w_1_600_s_2_400=2.00e-05 mcrdlm5m1_cc_w_1_600_s_2_400=4.63e-11 mcrdlm5m1_cf_w_1_600_s_2_400=2.06e-11
+  mcrdlm5m1_ca_w_1_600_s_2_800=2.00e-05 mcrdlm5m1_cc_w_1_600_s_2_800=3.80e-11 mcrdlm5m1_cf_w_1_600_s_2_800=2.36e-11
+  mcrdlm5m1_ca_w_1_600_s_3_200=2.00e-05 mcrdlm5m1_cc_w_1_600_s_3_200=3.17e-11 mcrdlm5m1_cf_w_1_600_s_3_200=2.63e-11
+  mcrdlm5m1_ca_w_1_600_s_4_800=2.00e-05 mcrdlm5m1_cc_w_1_600_s_4_800=1.64e-11 mcrdlm5m1_cf_w_1_600_s_4_800=3.51e-11
+  mcrdlm5m1_ca_w_1_600_s_10_000=2.00e-05 mcrdlm5m1_cc_w_1_600_s_10_000=2.40e-12 mcrdlm5m1_cf_w_1_600_s_10_000=4.68e-11
+  mcrdlm5m1_ca_w_1_600_s_12_000=2.00e-05 mcrdlm5m1_cc_w_1_600_s_12_000=1.13e-12 mcrdlm5m1_cf_w_1_600_s_12_000=4.79e-11
+  mcrdlm5m1_ca_w_4_000_s_1_600=2.00e-05 mcrdlm5m1_cc_w_4_000_s_1_600=7.66e-11 mcrdlm5m1_cf_w_4_000_s_1_600=1.40e-11
+  mcrdlm5m1_ca_w_4_000_s_1_700=2.00e-05 mcrdlm5m1_cc_w_4_000_s_1_700=7.10e-11 mcrdlm5m1_cf_w_4_000_s_1_700=1.49e-11
+  mcrdlm5m1_ca_w_4_000_s_1_900=2.00e-05 mcrdlm5m1_cc_w_4_000_s_1_900=6.25e-11 mcrdlm5m1_cf_w_4_000_s_1_900=1.66e-11
+  mcrdlm5m1_ca_w_4_000_s_2_000=2.00e-05 mcrdlm5m1_cc_w_4_000_s_2_000=5.88e-11 mcrdlm5m1_cf_w_4_000_s_2_000=1.74e-11
+  mcrdlm5m1_ca_w_4_000_s_2_400=2.00e-05 mcrdlm5m1_cc_w_4_000_s_2_400=4.71e-11 mcrdlm5m1_cf_w_4_000_s_2_400=2.06e-11
+  mcrdlm5m1_ca_w_4_000_s_2_800=2.00e-05 mcrdlm5m1_cc_w_4_000_s_2_800=3.87e-11 mcrdlm5m1_cf_w_4_000_s_2_800=2.37e-11
+  mcrdlm5m1_ca_w_4_000_s_3_200=2.00e-05 mcrdlm5m1_cc_w_4_000_s_3_200=3.23e-11 mcrdlm5m1_cf_w_4_000_s_3_200=2.64e-11
+  mcrdlm5m1_ca_w_4_000_s_4_800=2.00e-05 mcrdlm5m1_cc_w_4_000_s_4_800=1.68e-11 mcrdlm5m1_cf_w_4_000_s_4_800=3.53e-11
+  mcrdlm5m1_ca_w_4_000_s_10_000=2.00e-05 mcrdlm5m1_cc_w_4_000_s_10_000=2.43e-12 mcrdlm5m1_cf_w_4_000_s_10_000=4.71e-11
+  mcrdlm5m1_ca_w_4_000_s_12_000=2.00e-05 mcrdlm5m1_cc_w_4_000_s_12_000=1.16e-12 mcrdlm5m1_cf_w_4_000_s_12_000=4.84e-11
+  mcrdlm5m2_ca_w_1_600_s_1_600=2.21e-05 mcrdlm5m2_cc_w_1_600_s_1_600=7.35e-11 mcrdlm5m2_cf_w_1_600_s_1_600=1.54e-11
+  mcrdlm5m2_ca_w_1_600_s_1_700=2.21e-05 mcrdlm5m2_cc_w_1_600_s_1_700=6.82e-11 mcrdlm5m2_cf_w_1_600_s_1_700=1.64e-11
+  mcrdlm5m2_ca_w_1_600_s_1_900=2.21e-05 mcrdlm5m2_cc_w_1_600_s_1_900=5.96e-11 mcrdlm5m2_cf_w_1_600_s_1_900=1.82e-11
+  mcrdlm5m2_ca_w_1_600_s_2_000=2.21e-05 mcrdlm5m2_cc_w_1_600_s_2_000=5.60e-11 mcrdlm5m2_cf_w_1_600_s_2_000=1.91e-11
+  mcrdlm5m2_ca_w_1_600_s_2_400=2.21e-05 mcrdlm5m2_cc_w_1_600_s_2_400=4.45e-11 mcrdlm5m2_cf_w_1_600_s_2_400=2.26e-11
+  mcrdlm5m2_ca_w_1_600_s_2_800=2.21e-05 mcrdlm5m2_cc_w_1_600_s_2_800=3.63e-11 mcrdlm5m2_cf_w_1_600_s_2_800=2.58e-11
+  mcrdlm5m2_ca_w_1_600_s_3_200=2.21e-05 mcrdlm5m2_cc_w_1_600_s_3_200=3.00e-11 mcrdlm5m2_cf_w_1_600_s_3_200=2.87e-11
+  mcrdlm5m2_ca_w_1_600_s_4_800=2.21e-05 mcrdlm5m2_cc_w_1_600_s_4_800=1.50e-11 mcrdlm5m2_cf_w_1_600_s_4_800=3.79e-11
+  mcrdlm5m2_ca_w_1_600_s_10_000=2.21e-05 mcrdlm5m2_cc_w_1_600_s_10_000=1.92e-12 mcrdlm5m2_cf_w_1_600_s_10_000=4.89e-11
+  mcrdlm5m2_ca_w_1_600_s_12_000=2.21e-05 mcrdlm5m2_cc_w_1_600_s_12_000=8.45e-13 mcrdlm5m2_cf_w_1_600_s_12_000=5.00e-11
+  mcrdlm5m2_ca_w_4_000_s_1_600=2.21e-05 mcrdlm5m2_cc_w_4_000_s_1_600=7.47e-11 mcrdlm5m2_cf_w_4_000_s_1_600=1.55e-11
+  mcrdlm5m2_ca_w_4_000_s_1_700=2.21e-05 mcrdlm5m2_cc_w_4_000_s_1_700=6.93e-11 mcrdlm5m2_cf_w_4_000_s_1_700=1.64e-11
+  mcrdlm5m2_ca_w_4_000_s_1_900=2.21e-05 mcrdlm5m2_cc_w_4_000_s_1_900=6.05e-11 mcrdlm5m2_cf_w_4_000_s_1_900=1.82e-11
+  mcrdlm5m2_ca_w_4_000_s_2_000=2.21e-05 mcrdlm5m2_cc_w_4_000_s_2_000=5.70e-11 mcrdlm5m2_cf_w_4_000_s_2_000=1.91e-11
+  mcrdlm5m2_ca_w_4_000_s_2_400=2.21e-05 mcrdlm5m2_cc_w_4_000_s_2_400=4.53e-11 mcrdlm5m2_cf_w_4_000_s_2_400=2.26e-11
+  mcrdlm5m2_ca_w_4_000_s_2_800=2.21e-05 mcrdlm5m2_cc_w_4_000_s_2_800=3.69e-11 mcrdlm5m2_cf_w_4_000_s_2_800=2.58e-11
+  mcrdlm5m2_ca_w_4_000_s_3_200=2.21e-05 mcrdlm5m2_cc_w_4_000_s_3_200=3.05e-11 mcrdlm5m2_cf_w_4_000_s_3_200=2.88e-11
+  mcrdlm5m2_ca_w_4_000_s_4_800=2.21e-05 mcrdlm5m2_cc_w_4_000_s_4_800=1.53e-11 mcrdlm5m2_cf_w_4_000_s_4_800=3.80e-11
+  mcrdlm5m2_ca_w_4_000_s_10_000=2.21e-05 mcrdlm5m2_cc_w_4_000_s_10_000=1.96e-12 mcrdlm5m2_cf_w_4_000_s_10_000=4.93e-11
+  mcrdlm5m2_ca_w_4_000_s_12_000=2.21e-05 mcrdlm5m2_cc_w_4_000_s_12_000=8.90e-13 mcrdlm5m2_cf_w_4_000_s_12_000=5.03e-11
+  mcrdlm5m3_ca_w_1_600_s_1_600=3.34e-05 mcrdlm5m3_cc_w_1_600_s_1_600=6.72e-11 mcrdlm5m3_cf_w_1_600_s_1_600=2.23e-11
+  mcrdlm5m3_ca_w_1_600_s_1_700=3.34e-05 mcrdlm5m3_cc_w_1_600_s_1_700=6.20e-11 mcrdlm5m3_cf_w_1_600_s_1_700=2.36e-11
+  mcrdlm5m3_ca_w_1_600_s_1_900=3.34e-05 mcrdlm5m3_cc_w_1_600_s_1_900=5.33e-11 mcrdlm5m3_cf_w_1_600_s_1_900=2.61e-11
+  mcrdlm5m3_ca_w_1_600_s_2_000=3.34e-05 mcrdlm5m3_cc_w_1_600_s_2_000=4.96e-11 mcrdlm5m3_cf_w_1_600_s_2_000=2.73e-11
+  mcrdlm5m3_ca_w_1_600_s_2_400=3.34e-05 mcrdlm5m3_cc_w_1_600_s_2_400=3.82e-11 mcrdlm5m3_cf_w_1_600_s_2_400=3.19e-11
+  mcrdlm5m3_ca_w_1_600_s_2_800=3.34e-05 mcrdlm5m3_cc_w_1_600_s_2_800=3.02e-11 mcrdlm5m3_cf_w_1_600_s_2_800=3.58e-11
+  mcrdlm5m3_ca_w_1_600_s_3_200=3.34e-05 mcrdlm5m3_cc_w_1_600_s_3_200=2.41e-11 mcrdlm5m3_cf_w_1_600_s_3_200=3.94e-11
+  mcrdlm5m3_ca_w_1_600_s_4_800=3.34e-05 mcrdlm5m3_cc_w_1_600_s_4_800=1.05e-11 mcrdlm5m3_cf_w_1_600_s_4_800=4.92e-11
+  mcrdlm5m3_ca_w_1_600_s_10_000=3.34e-05 mcrdlm5m3_cc_w_1_600_s_10_000=8.80e-13 mcrdlm5m3_cf_w_1_600_s_10_000=5.79e-11
+  mcrdlm5m3_ca_w_1_600_s_12_000=3.34e-05 mcrdlm5m3_cc_w_1_600_s_12_000=3.15e-13 mcrdlm5m3_cf_w_1_600_s_12_000=5.85e-11
+  mcrdlm5m3_ca_w_4_000_s_1_600=3.34e-05 mcrdlm5m3_cc_w_4_000_s_1_600=6.81e-11 mcrdlm5m3_cf_w_4_000_s_1_600=2.23e-11
+  mcrdlm5m3_ca_w_4_000_s_1_700=3.34e-05 mcrdlm5m3_cc_w_4_000_s_1_700=6.28e-11 mcrdlm5m3_cf_w_4_000_s_1_700=2.36e-11
+  mcrdlm5m3_ca_w_4_000_s_1_900=3.34e-05 mcrdlm5m3_cc_w_4_000_s_1_900=5.42e-11 mcrdlm5m3_cf_w_4_000_s_1_900=2.61e-11
+  mcrdlm5m3_ca_w_4_000_s_2_000=3.34e-05 mcrdlm5m3_cc_w_4_000_s_2_000=5.04e-11 mcrdlm5m3_cf_w_4_000_s_2_000=2.74e-11
+  mcrdlm5m3_ca_w_4_000_s_2_400=3.34e-05 mcrdlm5m3_cc_w_4_000_s_2_400=3.89e-11 mcrdlm5m3_cf_w_4_000_s_2_400=3.19e-11
+  mcrdlm5m3_ca_w_4_000_s_2_800=3.34e-05 mcrdlm5m3_cc_w_4_000_s_2_800=3.07e-11 mcrdlm5m3_cf_w_4_000_s_2_800=3.59e-11
+  mcrdlm5m3_ca_w_4_000_s_3_200=3.34e-05 mcrdlm5m3_cc_w_4_000_s_3_200=2.45e-11 mcrdlm5m3_cf_w_4_000_s_3_200=3.95e-11
+  mcrdlm5m3_ca_w_4_000_s_4_800=3.34e-05 mcrdlm5m3_cc_w_4_000_s_4_800=1.08e-11 mcrdlm5m3_cf_w_4_000_s_4_800=4.93e-11
+  mcrdlm5m3_ca_w_4_000_s_10_000=3.34e-05 mcrdlm5m3_cc_w_4_000_s_10_000=8.85e-13 mcrdlm5m3_cf_w_4_000_s_10_000=5.83e-11
+  mcrdlm5m3_ca_w_4_000_s_12_000=3.34e-05 mcrdlm5m3_cc_w_4_000_s_12_000=3.55e-13 mcrdlm5m3_cf_w_4_000_s_12_000=5.89e-11
+  mcrdlm5m4_ca_w_1_600_s_1_600=1.24e-04 mcrdlm5m4_cc_w_1_600_s_1_600=5.14e-11 mcrdlm5m4_cf_w_1_600_s_1_600=5.78e-11
+  mcrdlm5m4_ca_w_1_600_s_1_700=1.24e-04 mcrdlm5m4_cc_w_1_600_s_1_700=4.64e-11 mcrdlm5m4_cf_w_1_600_s_1_700=6.00e-11
+  mcrdlm5m4_ca_w_1_600_s_1_900=1.24e-04 mcrdlm5m4_cc_w_1_600_s_1_900=3.83e-11 mcrdlm5m4_cf_w_1_600_s_1_900=6.41e-11
+  mcrdlm5m4_ca_w_1_600_s_2_000=1.24e-04 mcrdlm5m4_cc_w_1_600_s_2_000=3.49e-11 mcrdlm5m4_cf_w_1_600_s_2_000=6.61e-11
+  mcrdlm5m4_ca_w_1_600_s_2_400=1.24e-04 mcrdlm5m4_cc_w_1_600_s_2_400=2.49e-11 mcrdlm5m4_cf_w_1_600_s_2_400=7.24e-11
+  mcrdlm5m4_ca_w_1_600_s_2_800=1.24e-04 mcrdlm5m4_cc_w_1_600_s_2_800=1.83e-11 mcrdlm5m4_cf_w_1_600_s_2_800=7.72e-11
+  mcrdlm5m4_ca_w_1_600_s_3_200=1.24e-04 mcrdlm5m4_cc_w_1_600_s_3_200=1.36e-11 mcrdlm5m4_cf_w_1_600_s_3_200=8.09e-11
+  mcrdlm5m4_ca_w_1_600_s_4_800=1.24e-04 mcrdlm5m4_cc_w_1_600_s_4_800=4.57e-12 mcrdlm5m4_cf_w_1_600_s_4_800=8.89e-11
+  mcrdlm5m4_ca_w_1_600_s_10_000=1.24e-04 mcrdlm5m4_cc_w_1_600_s_10_000=2.10e-13 mcrdlm5m4_cf_w_1_600_s_10_000=9.34e-11
+  mcrdlm5m4_ca_w_1_600_s_12_000=1.24e-04 mcrdlm5m4_cc_w_1_600_s_12_000=7.50e-14 mcrdlm5m4_cf_w_1_600_s_12_000=9.36e-11
+  mcrdlm5m4_ca_w_4_000_s_1_600=1.24e-04 mcrdlm5m4_cc_w_4_000_s_1_600=5.23e-11 mcrdlm5m4_cf_w_4_000_s_1_600=5.77e-11
+  mcrdlm5m4_ca_w_4_000_s_1_700=1.24e-04 mcrdlm5m4_cc_w_4_000_s_1_700=4.73e-11 mcrdlm5m4_cf_w_4_000_s_1_700=6.01e-11
+  mcrdlm5m4_ca_w_4_000_s_1_900=1.24e-04 mcrdlm5m4_cc_w_4_000_s_1_900=3.90e-11 mcrdlm5m4_cf_w_4_000_s_1_900=6.42e-11
+  mcrdlm5m4_ca_w_4_000_s_2_000=1.24e-04 mcrdlm5m4_cc_w_4_000_s_2_000=3.58e-11 mcrdlm5m4_cf_w_4_000_s_2_000=6.61e-11
+  mcrdlm5m4_ca_w_4_000_s_2_400=1.24e-04 mcrdlm5m4_cc_w_4_000_s_2_400=2.55e-11 mcrdlm5m4_cf_w_4_000_s_2_400=7.24e-11
+  mcrdlm5m4_ca_w_4_000_s_2_800=1.24e-04 mcrdlm5m4_cc_w_4_000_s_2_800=1.88e-11 mcrdlm5m4_cf_w_4_000_s_2_800=7.73e-11
+  mcrdlm5m4_ca_w_4_000_s_3_200=1.24e-04 mcrdlm5m4_cc_w_4_000_s_3_200=1.40e-11 mcrdlm5m4_cf_w_4_000_s_3_200=8.10e-11
+  mcrdlm5m4_ca_w_4_000_s_4_800=1.24e-04 mcrdlm5m4_cc_w_4_000_s_4_800=4.81e-12 mcrdlm5m4_cf_w_4_000_s_4_800=8.92e-11
+  mcrdlm5m4_ca_w_4_000_s_10_000=1.24e-04 mcrdlm5m4_cc_w_4_000_s_10_000=2.30e-13 mcrdlm5m4_cf_w_4_000_s_10_000=9.39e-11
+  mcrdlm5m4_ca_w_4_000_s_12_000=1.24e-04 mcrdlm5m4_cc_w_4_000_s_12_000=9.50e-14 mcrdlm5m4_cf_w_4_000_s_12_000=9.41e-11
+  cp1f=1.55e-04 cp1fsw=1.02e-10
+  cl1f=4.97e-05 cl1fsw=1.04e-10
+  cl1d=7.09e-05 cl1dsw=1.03e-10
+  cl1p1=1.74e-04 cl1p1sw=1.02e-10
+  cm1f=3.57e-05 cm1fsw=1.32e-10
+  cm1d=4.54e-05 cm1dsw=1.31e-10
+  cm1p1=7.32e-05 cm1p1sw=1.30e-10
+  cm1l1=2.15e-04 cm1l1sw=1.26e-10
+  cm2f=2.35e-05 cm2fsw=1.33e-10
+  cm2d=2.74e-05 cm2dsw=1.32e-10
+  cm2p1=3.55e-05 cm2p1sw=1.32e-10
+  cm2l1=5.23e-05 cm2l1sw=1.31e-10
+  cm2m1=3.13e-04 cm2m1sw=1.26e-10
+  cm3f=1.63e-05 cm3fsw=1.26e-10
+  cm3d=1.81e-05 cm3dsw=1.26e-10
+  cm3p1=2.13e-05 cm3p1sw=1.25e-10
+  cm3l1=2.63e-05 cm3l1sw=1.25e-10
+  cm3m1=4.52e-05 cm3m1sw=1.23e-10
+  cm3m2=1.31e-04 cm3m2sw=1.22e-10
+  cm4f=1.07e-05 cm4fsw=1.29e-10
+  cm4d=1.14e-05 cm4dsw=1.28e-10
+  cm4p1=1.26e-05 cm4p1sw=1.28e-10
+  cm4l1=1.43e-05 cm4l1sw=1.28e-10
+  cm4m1=1.85e-05 cm4m1sw=1.27e-10
+  cm4m2=2.52e-05 cm4m2sw=1.27e-10
+  cm4m3=1.91e-04 cm4m3sw=1.25e-10
+  cm5f=7.76e-06 cm5fsw=9.43e-11
+  cm5d=8.14e-06 cm5dsw=9.41e-11
+  cm5p1=8.74e-06 cm5p1sw=9.39e-11
+  cm5l1=9.48e-06 cm5l1sw=9.37e-11
+  cm5m1=1.12e-05 cm5m1sw=9.32e-11
+  cm5m2=1.33e-05 cm5m2sw=9.29e-11
+  cm5m3=2.46e-05 cm5m3sw=9.33e-11
+  cm5m4=1.15e-04 cm5m4sw=1.13e-10
+  crdlf=3.49e-06 crdlfsw=7.63e-11
+  crdld=3.57e-06 crdldsw=7.61e-11
+  crdlp1=3.67e-06 crdlp1sw=7.60e-11
+  crdll1=3.80e-06 crdll1sw=7.59e-11
+  crdlm1=4.04e-06 crdlm1sw=7.57e-11
+  crdlm2=4.29e-06 crdlm2sw=7.54e-11
+  crdlm3=5.04e-06 crdlm3sw=7.51e-11
+  crdlm4=6.01e-06 crdlm4sw=7.48e-11
+  crdlm5=8.81e-06 crdlm5sw=7.52e-11
+  cl1p1f=3.29e-04 cl1p1fsw=9.71e-11
+  cm1p1f=2.29e-04 cm1p1fsw=9.88e-11
+  cm2p1f=1.91e-04 cm2p1fsw=1.01e-10
+  cm3p1f=1.76e-04 cm3p1fsw=1.01e-10
+  cm4p1f=1.67e-04 cm4p1fsw=1.02e-10
+  cm5p1f=1.64e-04 cm5p1fsw=1.02e-10
+  crdlp1f=1.58e-04 crdlp1fsw=1.02e-10
+  cm1l1f=2.66e-04 cm1l1fsw=9.75e-11
+  cm1l1d=2.87e-04 cm1l1dsw=9.64e-11
+  cm1l1p1=3.91e-04 cm1l1p1sw=9.52e-11
+  cm2l1f=1.02e-04 cm2l1fsw=1.01e-10
+  cm2l1d=1.23e-04 cm2l1dsw=9.99e-11
+  cm2l1p1=2.27e-04 cm2l1p1sw=9.88e-11
+  cm3l1f=7.60e-05 cm3l1fsw=1.03e-10
+  cm3l1d=9.72e-05 cm3l1dsw=1.02e-10
+  cm3l1p1=2.01e-04 cm3l1p1sw=1.01e-10
+  cm4l1f=6.40e-05 cm4l1fsw=1.03e-10
+  cm4l1d=8.52e-05 cm4l1dsw=1.02e-10
+  cm4l1p1=1.88e-04 cm4l1p1sw=1.01e-10
+  cm5l1f=5.92e-05 cm5l1fsw=1.04e-10
+  cm5l1d=8.04e-05 cm5l1dsw=1.03e-10
+  cm5l1p1=1.84e-04 cm5l1p1sw=1.02e-10
+  crdll1f=5.35e-05 crdll1fsw=1.04e-10
+  crdll1d=7.47e-05 crdll1dsw=1.03e-10
+  crdll1p1=1.78e-04 crdll1p1sw=1.02e-10
+  cm2m1f=3.49e-04 cm2m1fsw=1.24e-10
+  cm2m1d=3.58e-04 cm2m1dsw=1.23e-10
+  cm2m1p1=3.86e-04 cm2m1p1sw=1.21e-10
+  cm2m1l1=5.28e-04 cm2m1l1sw=1.18e-10
+  cm3m1f=8.09e-05 cm3m1fsw=1.29e-10
+  cm3m1d=9.07e-05 cm3m1dsw=1.29e-10
+  cm3m1p1=1.18e-04 cm3m1p1sw=1.25e-10
+  cm3m1l1=2.60e-04 cm3m1l1sw=1.22e-10
+  cm4m1f=5.42e-05 cm4m1fsw=1.31e-10
+  cm4m1d=6.39e-05 cm4m1dsw=1.30e-10
+  cm4m1p1=9.17e-05 cm4m1p1sw=1.27e-10
+  cm4m1l1=2.34e-04 cm4m1l1sw=1.24e-10
+  cm5m1f=4.68e-05 cm5m1fsw=1.32e-10
+  cm5m1d=5.66e-05 cm5m1dsw=1.31e-10
+  cm5m1p1=8.43e-05 cm5m1p1sw=1.28e-10
+  cm5m1l1=2.26e-04 cm5m1l1sw=1.25e-10
+  crdlm1f=3.97e-05 crdlm1fsw=1.33e-10
+  crdlm1d=4.95e-05 crdlm1dsw=1.32e-10
+  crdlm1p1=7.72e-05 crdlm1p1sw=1.28e-10
+  crdlm1l1=2.19e-04 crdlm1l1sw=1.25e-10
+  cm3m2f=1.55e-04 cm3m2fsw=1.26e-10
+  cm3m2d=1.59e-04 cm3m2dsw=1.26e-10
+  cm3m2p1=1.67e-04 cm3m2p1sw=1.25e-10
+  cm3m2l1=1.83e-04 cm3m2l1sw=1.23e-10
+  cm3m2m1=4.44e-04 cm3m2m1sw=1.20e-10
+  cm4m2f=4.88e-05 cm4m2fsw=1.31e-10
+  cm4m2d=5.26e-05 cm4m2dsw=1.30e-10
+  cm4m2p1=6.08e-05 cm4m2p1sw=1.32e-10
+  cm4m2l1=7.75e-05 cm4m2l1sw=1.28e-10
+  cm4m2m1=3.38e-04 cm4m2m1sw=1.23e-10
+  cm5m2f=3.68e-05 cm5m2fsw=1.32e-10
+  cm5m2d=4.07e-05 cm5m2dsw=1.31e-10
+  cm5m2p1=4.89e-05 cm5m2p1sw=1.32e-10
+  cm5m2l1=6.56e-05 cm5m2l1sw=1.29e-10
+  cm5m2m1=3.26e-04 cm5m2m1sw=1.24e-10
+  crdlm2f=2.78e-05 crdlm2fsw=1.33e-10
+  crdlm2d=3.17e-05 crdlm2dsw=1.33e-10
+  crdlm2p1=3.98e-05 crdlm2p1sw=1.33e-10
+  crdlm2l1=5.66e-05 crdlm2l1sw=1.29e-10
+  crdlm2m1=3.17e-04 crdlm2m1sw=1.25e-10
+  cm4m3f=2.08e-04 cm4m3fsw=1.19e-10
+  cm4m3d=2.09e-04 cm4m3dsw=1.19e-10
+  cm4m3p1=2.13e-04 cm4m3p1sw=1.19e-10
+  cm4m3l1=2.18e-04 cm4m3l1sw=1.18e-10
+  cm4m3m1=2.37e-04 cm4m3m1sw=1.16e-10
+  cm4m3m2=3.22e-04 cm4m3m2sw=1.15e-10
+  cm5m3f=4.08e-05 cm5m3fsw=1.23e-10
+  cm5m3d=4.26e-05 cm5m3dsw=1.23e-10
+  cm5m3p1=4.58e-05 cm5m3p1sw=1.22e-10
+  cm5m3l1=5.08e-05 cm5m3l1sw=1.21e-10
+  cm5m3m1=6.98e-05 cm5m3m1sw=1.20e-10
+  cm5m3m2=1.56e-04 cm5m3m2sw=1.18e-10
+  crdlm3f=2.13e-05 crdlm3fsw=1.25e-10
+  crdlm3d=2.31e-05 crdlm3dsw=1.25e-10
+  crdlm3p1=2.63e-05 crdlm3p1sw=1.25e-10
+  crdlm3l1=3.13e-05 crdlm3l1sw=1.24e-10
+  crdlm3m1=5.02e-05 crdlm3m1sw=1.22e-10
+  crdlm3m2=1.36e-04 crdlm3m2sw=1.21e-10
+  cm5m4f=1.26e-04 cm5m4fsw=1.20e-10
+  cm5m4d=1.26e-04 cm5m4dsw=1.19e-10
+  cm5m4p1=1.27e-04 cm5m4p1sw=1.19e-10
+  cm5m4l1=1.29e-04 cm5m4l1sw=1.19e-10
+  cm5m4m1=1.33e-04 cm5m4m1sw=1.19e-10
+  cm5m4m2=1.40e-04 cm5m4m2sw=1.18e-10
+  cm5m4m3=3.06e-04 cm5m4m3sw=1.16e-10
+  crdlm4f=1.67e-05 crdlm4fsw=1.28e-10
+  crdlm4d=1.74e-05 crdlm4dsw=1.27e-10
+  crdlm4p1=1.87e-05 crdlm4p1sw=1.27e-10
+  crdlm4l1=2.03e-05 crdlm4l1sw=1.27e-10
+  crdlm4m1=2.45e-05 crdlm4m1sw=1.27e-10
+  crdlm4m2=3.12e-05 crdlm4m2sw=1.26e-10
+  crdlm4m3=1.97e-04 crdlm4m3sw=1.24e-10
+  crdlm5f=1.66e-05 crdlm5fsw=9.01e-11
+  crdlm5d=1.70e-05 crdlm5dsw=8.99e-11
+  crdlm5p1=1.76e-05 crdlm5p1sw=8.98e-11
+  crdlm5l1=1.83e-05 crdlm5l1sw=8.95e-11
+  crdlm5m1=2.00e-05 crdlm5m1sw=8.92e-11
+  crdlm5m2=2.21e-05 crdlm5m2sw=8.89e-11
+  crdlm5m3=3.34e-05 crdlm5m3sw=8.95e-11
+  crdlm5m4=1.24e-04 crdlm5m4sw=1.09e-10
