* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 49
.param
+  sky130_fd_pr__pfet_g5v0d10v5__toxe_mult=0.94
+  sky130_fd_pr__pfet_g5v0d10v5__rshp_mult=1.0
+  sky130_fd_pr__pfet_g5v0d10v5__overlap_mult=0.70
+  sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult=9.3222e-1
+  sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult=9.4436e-1
+  sky130_fd_pr__pfet_g5v0d10v5__lint_diff=1.7325e-8
+  sky130_fd_pr__pfet_g5v0d10v5__wint_diff=-3.2175e-8
+  sky130_fd_pr__pfet_g5v0d10v5__dlc_diff=1.7325e-8
+  sky130_fd_pr__pfet_g5v0d10v5__dwc_diff=-3.2175e-8
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 000, W = 10.0, L = 0.5
* -------------------------------
+  sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_0=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_0=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ub_diff_0=-8.1068e-19
+  sky130_fd_pr__pfet_g5v0d10v5__ua_diff_0=-5.8946e-13
+  sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_0=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__keta_diff_0=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_0=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_0=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_0=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__a0_diff_0=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_0=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b0_diff_0=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__k2_diff_0=0.019265
+  sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_0=0.92279
+  sky130_fd_pr__pfet_g5v0d10v5__u0_diff_0=-0.0024588
+  sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_0=0.029881
+  sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_0=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_0=-3965.1
+  sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_0=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__voff_diff_0=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b1_diff_0=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ags_diff_0=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_0=0.0
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 001, W = 15.0, L = 1.0
* -------------------------------
+  sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_1=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_1=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_1=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ub_diff_1=-1.0086e-19
+  sky130_fd_pr__pfet_g5v0d10v5__ua_diff_1=1.3345e-12
+  sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_1=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__keta_diff_1=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_1=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_1=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_1=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__a0_diff_1=-0.021649
+  sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_1=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b0_diff_1=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__k2_diff_1=0.0080331
+  sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_1=0.35569
+  sky130_fd_pr__pfet_g5v0d10v5__u0_diff_1=-0.00091756
+  sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_1=0.024505
+  sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_1=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_1=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_1=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__voff_diff_1=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b1_diff_1=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ags_diff_1=-0.034924
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 002, W = 15.0, L = 0.5
* -------------------------------
+  sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_2=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__voff_diff_2=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b1_diff_2=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ags_diff_2=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_2=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_2=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_2=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_2=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ub_diff_2=-6.4117e-19
+  sky130_fd_pr__pfet_g5v0d10v5__ua_diff_2=2.5554e-13
+  sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_2=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__keta_diff_2=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_2=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_2=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_2=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__a0_diff_2=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_2=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b0_diff_2=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__k2_diff_2=0.020797
+  sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_2=0.44022
+  sky130_fd_pr__pfet_g5v0d10v5__u0_diff_2=-0.0021939
+  sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_2=0.041746
+  sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_2=-3087.7
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 003, W = 1.5, L = 1.0
* ------------------------------
+  sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_3=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_3=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__voff_diff_3=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b1_diff_3=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ags_diff_3=-0.069521
+  sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_3=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_3=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_3=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_3=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ub_diff_3=-3.3536e-19
+  sky130_fd_pr__pfet_g5v0d10v5__ua_diff_3=2.7072e-13
+  sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_3=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__keta_diff_3=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_3=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_3=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_3=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__a0_diff_3=0.026441
+  sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_3=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b0_diff_3=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__k2_diff_3=0.0032184
+  sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_3=0.51928
+  sky130_fd_pr__pfet_g5v0d10v5__u0_diff_3=-0.0012151
+  sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_3=0.049005
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 004, W = 1.5, L = 2.0
* ------------------------------
+  sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_4=0.53933
+  sky130_fd_pr__pfet_g5v0d10v5__u0_diff_4=-0.00096391
+  sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_4=0.033612
+  sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_4=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_4=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__voff_diff_4=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b1_diff_4=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ags_diff_4=-0.031072
+  sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_4=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_4=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_4=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_4=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ub_diff_4=-3.0365e-19
+  sky130_fd_pr__pfet_g5v0d10v5__ua_diff_4=-1.9852e-13
+  sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_4=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__keta_diff_4=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_4=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_4=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_4=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__a0_diff_4=0.0069066
+  sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_4=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b0_diff_4=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__k2_diff_4=0.0026716
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 005, W = 1.5, L = 4.0
* ------------------------------
+  sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_5=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b0_diff_5=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__k2_diff_5=0.0047086
+  sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_5=0.62963
+  sky130_fd_pr__pfet_g5v0d10v5__u0_diff_5=-0.0018767
+  sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_5=0.035092
+  sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_5=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_5=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b1_diff_5=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ags_diff_5=0.00016238
+  sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_5=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_5=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__voff_diff_5=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_5=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_5=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ub_diff_5=-5.045e-19
+  sky130_fd_pr__pfet_g5v0d10v5__ua_diff_5=1.2416e-13
+  sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_5=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__keta_diff_5=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_5=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_5=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_5=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__a0_diff_5=-0.0002908
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 006, W = 1.5, L = 0.5
* ------------------------------
+  sky130_fd_pr__pfet_g5v0d10v5__a0_diff_6=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_6=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b0_diff_6=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__k2_diff_6=0.019041
+  sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_6=0.62826
+  sky130_fd_pr__pfet_g5v0d10v5__u0_diff_6=-0.0034483
+  sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_6=0.069383
+  sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_6=-9946.4
+  sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_6=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b1_diff_6=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ags_diff_6=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_6=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_6=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__voff_diff_6=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_6=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_6=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ub_diff_6=-1.1687e-18
+  sky130_fd_pr__pfet_g5v0d10v5__ua_diff_6=-2.1854e-12
+  sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_6=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__keta_diff_6=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_6=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_6=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_6=0.0
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 007, W = 1.0, L = 1.0
* ------------------------------
+  sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_7=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_7=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__a0_diff_7=-0.023831
+  sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_7=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b0_diff_7=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__k2_diff_7=0.0084689
+  sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_7=0.049563
+  sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_7=0.52602
+  sky130_fd_pr__pfet_g5v0d10v5__u0_diff_7=-0.0013725
+  sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_7=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_7=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b1_diff_7=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ags_diff_7=-0.047184
+  sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_7=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_7=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__voff_diff_7=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_7=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_7=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ub_diff_7=-4.2337e-19
+  sky130_fd_pr__pfet_g5v0d10v5__ua_diff_7=-3.5098e-13
+  sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_7=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__keta_diff_7=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_7=0.0
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 008, W = 1.0, L = 2.0
* ------------------------------
+  sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_8=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_8=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_8=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__a0_diff_8=-0.032394
+  sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_8=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b0_diff_8=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__k2_diff_8=0.0067604
+  sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_8=0.048453
+  sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_8=0.52597
+  sky130_fd_pr__pfet_g5v0d10v5__u0_diff_8=-0.0014593
+  sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_8=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_8=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b1_diff_8=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ags_diff_8=-0.053538
+  sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_8=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_8=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__voff_diff_8=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_8=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_8=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ub_diff_8=-5.0813e-19
+  sky130_fd_pr__pfet_g5v0d10v5__ua_diff_8=-5.8602e-13
+  sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_8=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__keta_diff_8=0.0
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 009, W = 1.0, L = 4.0
* ------------------------------
+  sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_9=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__keta_diff_9=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_9=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_9=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_9=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__a0_diff_9=0.0047331
+  sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_9=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b0_diff_9=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__k2_diff_9=0.0025401
+  sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_9=0.031854
+  sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_9=0.78025
+  sky130_fd_pr__pfet_g5v0d10v5__u0_diff_9=-0.0010746
+  sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_9=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_9=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b1_diff_9=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ags_diff_9=-0.025322
+  sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_9=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_9=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__voff_diff_9=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_9=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_9=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ub_diff_9=-2.6015e-19
+  sky130_fd_pr__pfet_g5v0d10v5__ua_diff_9=-2.9672e-14
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 010, W = 1.0, L = 8.0
* ------------------------------
+  sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_10=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_10=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__voff_diff_10=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b0_diff_10=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b1_diff_10=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_10=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_10=0.76718
+  sky130_fd_pr__pfet_g5v0d10v5__u0_diff_10=-0.0010652
+  sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_10=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_10=0.037456
+  sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_10=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ags_diff_10=-0.015852
+  sky130_fd_pr__pfet_g5v0d10v5__keta_diff_10=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_10=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__k2_diff_10=0.0033082
+  sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_10=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ua_diff_10=3.7574e-13
+  sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_10=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ub_diff_10=-1.9776e-19
+  sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_10=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_10=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_10=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__a0_diff_10=0.0022763
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 011, W = 1.0, L = 0.5
* ------------------------------
+  sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_11=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_11=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__a0_diff_11=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_11=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_11=-20938.0
+  sky130_fd_pr__pfet_g5v0d10v5__voff_diff_11=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b0_diff_11=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b1_diff_11=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_11=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_11=0.81024
+  sky130_fd_pr__pfet_g5v0d10v5__u0_diff_11=-0.0019065
+  sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_11=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_11=0.031367
+  sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_11=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ags_diff_11=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__keta_diff_11=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_11=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__k2_diff_11=0.019312
+  sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_11=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ua_diff_11=8.5779e-13
+  sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_11=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ub_diff_11=-4.1882e-19
+  sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_11=0.0
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 012, W = 1.0, L = 0.6
* ------------------------------
+  sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_12=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_12=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_12=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__a0_diff_12=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_12=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_12=-9517.3
+  sky130_fd_pr__pfet_g5v0d10v5__voff_diff_12=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b0_diff_12=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b1_diff_12=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_12=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_12=0.42675
+  sky130_fd_pr__pfet_g5v0d10v5__u0_diff_12=-0.0031096
+  sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_12=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_12=0.06505
+  sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_12=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ags_diff_12=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__keta_diff_12=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_12=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__k2_diff_12=0.011937
+  sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_12=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ua_diff_12=-8.4463e-13
+  sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_12=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ub_diff_12=-8.4748e-19
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 013, W = 1.0, L = 0.8
* ------------------------------
+  sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_13=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ub_diff_13=-6.9753e-19
+  sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_13=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_13=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_13=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__a0_diff_13=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_13=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_13=-4426.9
+  sky130_fd_pr__pfet_g5v0d10v5__voff_diff_13=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b0_diff_13=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b1_diff_13=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_13=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_13=0.34957
+  sky130_fd_pr__pfet_g5v0d10v5__u0_diff_13=-0.002059
+  sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_13=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_13=0.042239
+  sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_13=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ags_diff_13=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__keta_diff_13=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_13=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__k2_diff_13=0.012626
+  sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_13=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ua_diff_13=-1.3471e-12
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 014, W = 20.0, L = 1.0
* -------------------------------
+  sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_14=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ua_diff_14=6.5821e-13
+  sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_14=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ub_diff_14=-4.0194e-19
+  sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_14=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_14=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_14=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__a0_diff_14=-0.016665
+  sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_14=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_14=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__voff_diff_14=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b0_diff_14=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b1_diff_14=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_14=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_14=0.29074
+  sky130_fd_pr__pfet_g5v0d10v5__u0_diff_14=-0.0015647
+  sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_14=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_14=0.024415
+  sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_14=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ags_diff_14=-0.026998
+  sky130_fd_pr__pfet_g5v0d10v5__keta_diff_14=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_14=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__k2_diff_14=0.008511
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 015, W = 20.0, L = 0.5
* -------------------------------
+  sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_15=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ags_diff_15=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__keta_diff_15=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_15=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__k2_diff_15=0.018378
+  sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_15=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ua_diff_15=3.9683e-13
+  sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_15=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ub_diff_15=-7.8901e-19
+  sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_15=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_15=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_15=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__a0_diff_15=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_15=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_15=-3884.3
+  sky130_fd_pr__pfet_g5v0d10v5__voff_diff_15=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b0_diff_15=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b1_diff_15=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_15=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_15=0.85294
+  sky130_fd_pr__pfet_g5v0d10v5__u0_diff_15=-0.0027952
+  sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_15=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_15=0.026385
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 016, W = 3.0, L = 1.0
* ------------------------------
+  sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_16=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_16=0.040793
+  sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_16=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ags_diff_16=-0.030763
+  sky130_fd_pr__pfet_g5v0d10v5__keta_diff_16=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_16=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__k2_diff_16=0.008808
+  sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_16=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ua_diff_16=4.6538e-13
+  sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_16=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ub_diff_16=-6.6411e-19
+  sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_16=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_16=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_16=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__a0_diff_16=-0.016503
+  sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_16=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_16=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__voff_diff_16=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b0_diff_16=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b1_diff_16=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_16=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_16=0.49653
+  sky130_fd_pr__pfet_g5v0d10v5__u0_diff_16=-0.0025485
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 017, W = 3.0, L = 2.0
* ------------------------------
+  sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_17=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_17=0.15271
+  sky130_fd_pr__pfet_g5v0d10v5__u0_diff_17=-0.00068848
+  sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_17=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_17=0.022874
+  sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_17=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ags_diff_17=-0.013211
+  sky130_fd_pr__pfet_g5v0d10v5__keta_diff_17=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_17=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__k2_diff_17=0.0016068
+  sky130_fd_pr__pfet_g5v0d10v5__ua_diff_17=1.4383e-12
+  sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_17=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_17=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ub_diff_17=1.57e-20
+  sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_17=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_17=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_17=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__a0_diff_17=0.0015256
+  sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_17=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_17=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__voff_diff_17=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b0_diff_17=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b1_diff_17=0.0
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 018, W = 3.0, L = 4.0
* ------------------------------
+  sky130_fd_pr__pfet_g5v0d10v5__b1_diff_18=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_18=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_18=1.023
+  sky130_fd_pr__pfet_g5v0d10v5__u0_diff_18=-0.0021335
+  sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_18=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_18=0.041838
+  sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_18=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ags_diff_18=-0.0095856
+  sky130_fd_pr__pfet_g5v0d10v5__keta_diff_18=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_18=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__k2_diff_18=0.0029978
+  sky130_fd_pr__pfet_g5v0d10v5__ua_diff_18=4.4933e-13
+  sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_18=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_18=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ub_diff_18=-5.6175e-19
+  sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_18=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_18=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_18=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__a0_diff_18=0.0018439
+  sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_18=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_18=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__voff_diff_18=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b0_diff_18=0.0
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 019, W = 3.0, L = 8.0
* ------------------------------
+  sky130_fd_pr__pfet_g5v0d10v5__voff_diff_19=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b0_diff_19=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b1_diff_19=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_19=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_19=0.72939
+  sky130_fd_pr__pfet_g5v0d10v5__u0_diff_19=-0.0014519
+  sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_19=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_19=0.035431
+  sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_19=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ags_diff_19=-0.0050121
+  sky130_fd_pr__pfet_g5v0d10v5__keta_diff_19=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_19=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__k2_diff_19=0.00066506
+  sky130_fd_pr__pfet_g5v0d10v5__ua_diff_19=6.1444e-13
+  sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_19=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_19=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ub_diff_19=-3.157e-19
+  sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_19=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_19=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_19=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__a0_diff_19=0.00066294
+  sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_19=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_19=0.0
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 020, W = 3.0, L = 0.5
* ------------------------------
+  sky130_fd_pr__pfet_g5v0d10v5__voff_diff_20=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b0_diff_20=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b1_diff_20=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_20=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_20=0.92468
+  sky130_fd_pr__pfet_g5v0d10v5__u0_diff_20=-0.0021126
+  sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_20=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_20=0.024595
+  sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_20=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ags_diff_20=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__keta_diff_20=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_20=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__k2_diff_20=0.020516
+  sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_20=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ua_diff_20=1.4571e-12
+  sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_20=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ub_diff_20=-4.573e-19
+  sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_20=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_20=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_20=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__a0_diff_20=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_20=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_20=-23962.0
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 021, W = 3.0, L = 0.6
* ------------------------------
+  sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_21=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_21=-7800.3
+  sky130_fd_pr__pfet_g5v0d10v5__voff_diff_21=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b0_diff_21=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b1_diff_21=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_21=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_21=0.53151
+  sky130_fd_pr__pfet_g5v0d10v5__u0_diff_21=-0.0032065
+  sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_21=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_21=0.057297
+  sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_21=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ags_diff_21=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__keta_diff_21=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_21=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__k2_diff_21=0.015471
+  sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_21=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ua_diff_21=-5.568e-13
+  sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_21=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ub_diff_21=-8.928e-19
+  sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_21=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_21=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_21=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__a0_diff_21=0.0
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 022, W = 5.0, L = 1.0
* ------------------------------
+  sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_22=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_22=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__a0_diff_22=-0.010622
+  sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_22=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_22=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__voff_diff_22=-0.030587
+  sky130_fd_pr__pfet_g5v0d10v5__b0_diff_22=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b1_diff_22=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_22=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_22=0.25335
+  sky130_fd_pr__pfet_g5v0d10v5__u0_diff_22=-0.00011051
+  sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_22=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_22=0.0024631
+  sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_22=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ags_diff_22=-0.017178
+  sky130_fd_pr__pfet_g5v0d10v5__keta_diff_22=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_22=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__k2_diff_22=0.0040145
+  sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_22=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ua_diff_22=2.3221e-12
+  sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_22=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ub_diff_22=2.4278e-19
+  sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_22=0.0
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 023, W = 5.0, L = 2.0
* ------------------------------
+  sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_23=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_23=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_23=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__a0_diff_23=0.00021003
+  sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_23=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_23=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__voff_diff_23=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b0_diff_23=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b1_diff_23=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_23=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_23=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__u0_diff_23=-0.0011579
+  sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_23=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_23=0.018254
+  sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_23=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ags_diff_23=-0.0037978
+  sky130_fd_pr__pfet_g5v0d10v5__keta_diff_23=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_23=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__k2_diff_23=0.00031172
+  sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_23=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ua_diff_23=1.2987e-12
+  sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_23=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ub_diff_23=-2.3608e-19
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 024, W = 5.0, L = 4.0
* ------------------------------
+  sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_24=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ub_diff_24=-6.3305e-19
+  sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_24=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_24=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_24=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__a0_diff_24=0.0010943
+  sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_24=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_24=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__voff_diff_24=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b0_diff_24=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b1_diff_24=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_24=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_24=1.0538
+  sky130_fd_pr__pfet_g5v0d10v5__u0_diff_24=-0.0025093
+  sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_24=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_24=0.037325
+  sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_24=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ags_diff_24=-0.0034495
+  sky130_fd_pr__pfet_g5v0d10v5__keta_diff_24=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_24=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__k2_diff_24=0.0035991
+  sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_24=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ua_diff_24=8.8967e-13
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 025, W = 5.0, L = 8.0
* ------------------------------
+  sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_25=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ua_diff_25=8.0711e-13
+  sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_25=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ub_diff_25=-5.0441e-19
+  sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_25=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_25=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_25=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__a0_diff_25=-0.00085579
+  sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_25=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_25=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__voff_diff_25=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b0_diff_25=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b1_diff_25=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_25=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_25=0.72536
+  sky130_fd_pr__pfet_g5v0d10v5__u0_diff_25=-0.002061
+  sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_25=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_25=0.034248
+  sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_25=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ags_diff_25=0.0042769
+  sky130_fd_pr__pfet_g5v0d10v5__keta_diff_25=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_25=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__k2_diff_25=0.00052637
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 026, W = 5.0, L = 0.5
* ------------------------------
+  sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_26=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ags_diff_26=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__keta_diff_26=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_26=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__k2_diff_26=0.015878
+  sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_26=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ua_diff_26=2.7094e-12
+  sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_26=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ub_diff_26=-3.8525e-19
+  sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_26=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_26=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_26=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__a0_diff_26=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_26=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_26=-4782.4
+  sky130_fd_pr__pfet_g5v0d10v5__voff_diff_26=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b0_diff_26=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b1_diff_26=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_26=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_26=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__u0_diff_26=-0.0022969
+  sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_26=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_26=0.020333
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 027, W = 5.0, L = 0.6
* ------------------------------
+  sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_27=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_27=0.027956
+  sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_27=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ags_diff_27=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__keta_diff_27=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_27=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__k2_diff_27=0.015383
+  sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_27=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ua_diff_27=1.2388e-12
+  sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_27=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ub_diff_27=-1.4023e-18
+  sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_27=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_27=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_27=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__a0_diff_27=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_27=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_27=-2900.8
+  sky130_fd_pr__pfet_g5v0d10v5__voff_diff_27=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b0_diff_27=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b1_diff_27=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_27=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_27=0.51167
+  sky130_fd_pr__pfet_g5v0d10v5__u0_diff_27=-0.0047977
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 028, W = 5.0, L = 0.8
* ------------------------------
+  sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_28=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_28=0.32322
+  sky130_fd_pr__pfet_g5v0d10v5__u0_diff_28=-0.003291
+  sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_28=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_28=0.024803
+  sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_28=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ags_diff_28=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__keta_diff_28=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_28=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__k2_diff_28=0.0074048
+  sky130_fd_pr__pfet_g5v0d10v5__ua_diff_28=-5.0866e-13
+  sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_28=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_28=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ub_diff_28=-1.027e-18
+  sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_28=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_28=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_28=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__a0_diff_28=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_28=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_28=-3132.1
+  sky130_fd_pr__pfet_g5v0d10v5__voff_diff_28=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b0_diff_28=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b1_diff_28=0.0
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 029, W = 7.0, L = 1.0
* ------------------------------
+  sky130_fd_pr__pfet_g5v0d10v5__b1_diff_29=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_29=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_29=0.46918
+  sky130_fd_pr__pfet_g5v0d10v5__u0_diff_29=-0.0019752
+  sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_29=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_29=0.035895
+  sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_29=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ags_diff_29=-0.049364
+  sky130_fd_pr__pfet_g5v0d10v5__keta_diff_29=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_29=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__k2_diff_29=0.008623
+  sky130_fd_pr__pfet_g5v0d10v5__ua_diff_29=1.0863e-12
+  sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_29=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_29=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ub_diff_29=-4.4728e-19
+  sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_29=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_29=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_29=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__a0_diff_29=-0.030186
+  sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_29=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_29=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__voff_diff_29=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b0_diff_29=0.0
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 030, W = 7.0, L = 2.0
* ------------------------------
+  sky130_fd_pr__pfet_g5v0d10v5__voff_diff_30=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b0_diff_30=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b1_diff_30=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_30=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_30=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_30=0.12821
+  sky130_fd_pr__pfet_g5v0d10v5__u0_diff_30=-0.0011218
+  sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_30=0.016042
+  sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_30=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ags_diff_30=0.0034884
+  sky130_fd_pr__pfet_g5v0d10v5__keta_diff_30=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_30=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__k2_diff_30=0.00077199
+  sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_30=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ua_diff_30=1.0547e-12
+  sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_30=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ub_diff_30=-2.2772e-19
+  sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_30=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_30=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_30=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__a0_diff_30=-0.00085806
+  sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_30=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_30=0.0
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 031, W = 7.0, L = 4.0
* ------------------------------
+  sky130_fd_pr__pfet_g5v0d10v5__voff_diff_31=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b0_diff_31=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b1_diff_31=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_31=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_31=0.99463
+  sky130_fd_pr__pfet_g5v0d10v5__u0_diff_31=-0.002448
+  sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_31=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_31=0.036665
+  sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_31=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ags_diff_31=0.0079843
+  sky130_fd_pr__pfet_g5v0d10v5__keta_diff_31=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_31=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__k2_diff_31=0.0029578
+  sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_31=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ua_diff_31=1.463e-12
+  sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_31=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ub_diff_31=-5.4101e-19
+  sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_31=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_31=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_31=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__a0_diff_31=-0.0010532
+  sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_31=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_31=0.0
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 032, W = 7.0, L = 8.0
* ------------------------------
+  sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_32=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_32=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__voff_diff_32=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b0_diff_32=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b1_diff_32=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_32=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_32=0.71444
+  sky130_fd_pr__pfet_g5v0d10v5__u0_diff_32=-0.0019471
+  sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_32=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_32=0.035445
+  sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_32=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ags_diff_32=0.0068898
+  sky130_fd_pr__pfet_g5v0d10v5__keta_diff_32=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_32=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__k2_diff_32=0.00046848
+  sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_32=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ua_diff_32=1.0384e-12
+  sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_32=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ub_diff_32=-4.4536e-19
+  sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_32=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_32=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_32=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__a0_diff_32=-0.0013947
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 033, W = 7.0, L = 0.5
* ------------------------------
+  sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_33=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_33=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__a0_diff_33=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_33=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_33=-4311.0
+  sky130_fd_pr__pfet_g5v0d10v5__voff_diff_33=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b0_diff_33=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b1_diff_33=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_33=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_33=0.87408
+  sky130_fd_pr__pfet_g5v0d10v5__u0_diff_33=-0.0030453
+  sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_33=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_33=0.021812
+  sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_33=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ags_diff_33=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__keta_diff_33=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_33=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__k2_diff_33=0.019486
+  sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_33=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ua_diff_33=2.8817e-13
+  sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_33=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ub_diff_33=-8.2061e-19
+  sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_33=0.0
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 034, W = 7.0, L = 0.8
* ------------------------------
+  sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_34=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_34=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_34=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__a0_diff_34=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_34=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_34=-2734.0
+  sky130_fd_pr__pfet_g5v0d10v5__voff_diff_34=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b0_diff_34=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b1_diff_34=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_34=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_34=0.36517
+  sky130_fd_pr__pfet_g5v0d10v5__u0_diff_34=-0.003633
+  sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_34=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_34=0.032387
+  sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_34=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ags_diff_34=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__keta_diff_34=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_34=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__k2_diff_34=0.0080238
+  sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_34=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ua_diff_34=3.887e-13
+  sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_34=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ub_diff_34=-1.0184e-18
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 035, W = 0.42, L = 1.0
* -------------------------------
+  sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_35=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ub_diff_35=2.5095e-19
+  sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_35=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_35=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_35=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__a0_diff_35=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_35=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_35=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__voff_diff_35=-0.032724
+  sky130_fd_pr__pfet_g5v0d10v5__b0_diff_35=6.1346e-8
+  sky130_fd_pr__pfet_g5v0d10v5__b1_diff_35=1.2231e-9
+  sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_35=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_35=0.24131
+  sky130_fd_pr__pfet_g5v0d10v5__u0_diff_35=0.00083875
+  sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_35=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_35=0.028205
+  sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_35=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ags_diff_35=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__keta_diff_35=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_35=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__k2_diff_35=0.0035595
+  sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_35=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ua_diff_35=5.9894e-13
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 036, W = 0.42, L = 20.0
* --------------------------------
+  sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_36=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ua_diff_36=4.7238e-13
+  sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_36=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ub_diff_36=8.7499e-20
+  sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_36=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_36=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_36=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__a0_diff_36=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_36=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_36=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__voff_diff_36=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b0_diff_36=2.3627e-8
+  sky130_fd_pr__pfet_g5v0d10v5__b1_diff_36=1.0455e-9
+  sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_36=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_36=1.0069
+  sky130_fd_pr__pfet_g5v0d10v5__u0_diff_36=-5.5268e-5
+  sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_36=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_36=0.021615
+  sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_36=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ags_diff_36=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__keta_diff_36=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_36=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__k2_diff_36=-0.00025779
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 037, W = 0.42, L = 2.0
* -------------------------------
+  sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_37=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ags_diff_37=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__keta_diff_37=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_37=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__k2_diff_37=-0.0013459
+  sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_37=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ua_diff_37=-1.2717e-13
+  sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_37=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ub_diff_37=2.4827e-19
+  sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_37=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_37=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_37=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__a0_diff_37=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_37=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_37=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__voff_diff_37=-0.044516
+  sky130_fd_pr__pfet_g5v0d10v5__b0_diff_37=6.7541e-8
+  sky130_fd_pr__pfet_g5v0d10v5__b1_diff_37=6.4156e-8
+  sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_37=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_37=0.29283
+  sky130_fd_pr__pfet_g5v0d10v5__u0_diff_37=0.0009913
+  sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_37=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_37=0.036907
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 038, W = 0.42, L = 4.0
* -------------------------------
+  sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_38=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_38=0.031128
+  sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_38=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ags_diff_38=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__keta_diff_38=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_38=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__k2_diff_38=2.4551e-5
+  sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_38=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ua_diff_38=3.9386e-13
+  sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_38=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ub_diff_38=2.2142e-19
+  sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_38=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_38=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_38=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__a0_diff_38=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_38=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_38=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__voff_diff_38=-0.040882
+  sky130_fd_pr__pfet_g5v0d10v5__b0_diff_38=6.659e-8
+  sky130_fd_pr__pfet_g5v0d10v5__b1_diff_38=6.8754e-9
+  sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_38=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_38=0.24051
+  sky130_fd_pr__pfet_g5v0d10v5__u0_diff_38=0.00066016
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 039, W = 0.42, L = 8.0
* -------------------------------
+  sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_39=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_39=0.63931
+  sky130_fd_pr__pfet_g5v0d10v5__u0_diff_39=-0.00040288
+  sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_39=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_39=0.042789
+  sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_39=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ags_diff_39=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__keta_diff_39=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_39=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__k2_diff_39=0.0017461
+  sky130_fd_pr__pfet_g5v0d10v5__ua_diff_39=2.2233e-13
+  sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_39=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_39=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ub_diff_39=-6.3117e-20
+  sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_39=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_39=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_39=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__a0_diff_39=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_39=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_39=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__voff_diff_39=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b0_diff_39=6.3852e-8
+  sky130_fd_pr__pfet_g5v0d10v5__b1_diff_39=7.4391e-8
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 040, W = 0.42, L = 0.5
* -------------------------------
+  sky130_fd_pr__pfet_g5v0d10v5__b1_diff_40=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_40=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_40=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_40=0.71606
+  sky130_fd_pr__pfet_g5v0d10v5__u0_diff_40=-0.0042826
+  sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_40=0.14266
+  sky130_fd_pr__pfet_g5v0d10v5__keta_diff_40=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__k2_diff_40=0.031311
+  sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_40=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ags_diff_40=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_40=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_40=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ua_diff_40=-5.0918e-12
+  sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_40=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ub_diff_40=-1.8296e-18
+  sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_40=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_40=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_40=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__a0_diff_40=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_40=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_40=-18056.0
+  sky130_fd_pr__pfet_g5v0d10v5__voff_diff_40=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b0_diff_40=0.0
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 041, W = 0.42, L = 0.6
* -------------------------------
+  sky130_fd_pr__pfet_g5v0d10v5__voff_diff_41=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b0_diff_41=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b1_diff_41=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_41=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_41=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_41=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__u0_diff_41=0.00015782
+  sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_41=0.061213
+  sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_41=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ags_diff_41=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__keta_diff_41=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_41=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__k2_diff_41=0.013589
+  sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_41=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ua_diff_41=-2.67e-13
+  sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_41=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ub_diff_41=-8.3946e-20
+  sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_41=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_41=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_41=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__a0_diff_41=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_41=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_41=-11763.0
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 042, W = 0.42, L = 0.8
* -------------------------------
+  sky130_fd_pr__pfet_g5v0d10v5__voff_diff_42=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b0_diff_42=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b1_diff_42=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_42=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_42=0.83075
+  sky130_fd_pr__pfet_g5v0d10v5__u0_diff_42=-0.0014079
+  sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_42=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_42=0.090452
+  sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_42=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ags_diff_42=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__keta_diff_42=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_42=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__k2_diff_42=0.013318
+  sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_42=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ua_diff_42=2.5227e-12
+  sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_42=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ub_diff_42=-1.1626e-19
+  sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_42=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_42=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_42=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__a0_diff_42=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_42=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_42=-8835.0
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 043, W = 0.75, L = 1.0
* -------------------------------
+  sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_43=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_43=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__voff_diff_43=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b0_diff_43=2.3794e-7
+  sky130_fd_pr__pfet_g5v0d10v5__b1_diff_43=2.867e-10
+  sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_43=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_43=0.4302
+  sky130_fd_pr__pfet_g5v0d10v5__u0_diff_43=-0.0020643
+  sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_43=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_43=0.051387
+  sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_43=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ags_diff_43=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__keta_diff_43=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_43=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__k2_diff_43=0.0079272
+  sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_43=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ua_diff_43=-2.503e-12
+  sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_43=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ub_diff_43=-8.6763e-19
+  sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_43=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_43=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_43=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__a0_diff_43=0.0
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 044, W = 0.75, L = 2.0
* -------------------------------
+  sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_44=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_44=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__a0_diff_44=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_44=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_44=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__voff_diff_44=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b0_diff_44=1.5134e-7
+  sky130_fd_pr__pfet_g5v0d10v5__b1_diff_44=3.504e-10
+  sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_44=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_44=0.46436
+  sky130_fd_pr__pfet_g5v0d10v5__u0_diff_44=-0.0024078
+  sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_44=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_44=0.041458
+  sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_44=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ags_diff_44=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__keta_diff_44=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_44=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__k2_diff_44=0.0089111
+  sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_44=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ua_diff_44=-2.2688e-12
+  sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_44=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ub_diff_44=-9.51e-19
+  sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_44=0.0
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 045, W = 0.75, L = 4.0
* -------------------------------
+  sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_45=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_45=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_45=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__a0_diff_45=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_45=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_45=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__voff_diff_45=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b0_diff_45=9.3768e-8
+  sky130_fd_pr__pfet_g5v0d10v5__b1_diff_45=3.0925e-10
+  sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_45=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_45=0.77641
+  sky130_fd_pr__pfet_g5v0d10v5__u0_diff_45=-0.0012711
+  sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_45=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_45=0.041834
+  sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_45=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ags_diff_45=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__keta_diff_45=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_45=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__k2_diff_45=0.0053491
+  sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_45=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ua_diff_45=-8.113e-14
+  sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_45=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ub_diff_45=-3.3415e-19
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 046, W = 0.75, L = 0.5
* -------------------------------
+  sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_46=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ub_diff_46=-1.3254e-18
+  sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_46=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_46=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_46=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__a0_diff_46=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_46=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_46=-10829.0
+  sky130_fd_pr__pfet_g5v0d10v5__voff_diff_46=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b0_diff_46=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b1_diff_46=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_46=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_46=0.65931
+  sky130_fd_pr__pfet_g5v0d10v5__u0_diff_46=-0.0034037
+  sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_46=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_46=0.092606
+  sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_46=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ags_diff_46=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__keta_diff_46=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_46=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__k2_diff_46=0.023517
+  sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_46=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ua_diff_46=-3.6609e-12
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 047, W = 0.75, L = 0.8
* -------------------------------
+  sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_47=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ua_diff_47=-1.7538e-12
+  sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_47=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ub_diff_47=-1.0172e-18
+  sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_47=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_47=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_47=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__a0_diff_47=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_47=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_47=-11219.0
+  sky130_fd_pr__pfet_g5v0d10v5__voff_diff_47=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b0_diff_47=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b1_diff_47=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_47=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_47=0.44652
+  sky130_fd_pr__pfet_g5v0d10v5__u0_diff_47=-0.0030917
+  sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_47=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_47=0.05111
+  sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_47=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ags_diff_47=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__keta_diff_47=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_47=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__k2_diff_47=0.011414
*
* sky130_fd_pr__pfet_g5v0d10v5, Bin 048, W = 0.7, L = 0.6
* ------------------------------
+  sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_48=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ags_diff_48=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__keta_diff_48=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_48=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__k2_diff_48=0.011228
+  sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_48=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ua_diff_48=-2.9549e-14
+  sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_48=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__ub_diff_48=-1.2932e-19
+  sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_48=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_48=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_48=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__a0_diff_48=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_48=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_48=-8790.2
+  sky130_fd_pr__pfet_g5v0d10v5__voff_diff_48=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b0_diff_48=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__b1_diff_48=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_48=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_48=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__u0_diff_48=-0.00040428
+  sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_48=0.0
+  sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_48=0.033461
.include "sky130_fd_pr__pfet_g5v0d10v5.pm3.spice"
