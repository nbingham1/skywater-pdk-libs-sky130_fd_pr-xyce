* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 8
.param
+  sky130_fd_pr__rf_nfet_g5v0d10v5_b__toxe_mult=1.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_b__rbpb_mult=1.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult=0.89805
+  sky130_fd_pr__rf_nfet_g5v0d10v5_b__ajunction_mult=0.99505
+  sky130_fd_pr__rf_nfet_g5v0d10v5_b__pjunction_mult=1.0144
+  sky130_fd_pr__rf_nfet_g5v0d10v5_b__lint_diff=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_b__wint_diff=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_b__rshg_diff=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_b__xgw_diff=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_b__dlc_diff=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_b__dwc_diff=0.0
*
* sky130_fd_pr__rf_nfet_g5v0d10v5_bM02, Bin 000, W = 3.01, L = 0.5
* --------------------------------------------
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__voff_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__ub_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__vth0_diff_0=-0.015262
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__nfactor_diff_0=-0.36148
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__ua_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__vsat_diff_0=-3503.4
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__a0_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__rdsw_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__b0_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__ags_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__k2_diff_0=0.0013127
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__kt1_diff_0=-0.26612
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__pclm_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__u0_diff_0=-0.0029685
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__b1_diff_0=0.0
*
* sky130_fd_pr__rf_nfet_g5v0d10v5_bM02, Bin 001, W = 5.05, L = 0.5
* --------------------------------------------
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__b1_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__voff_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__ub_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__vth0_diff_1=-0.0025365
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__nfactor_diff_1=-0.53521
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__ua_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__vsat_diff_1=323.35
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__a0_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__rdsw_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__b0_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__ags_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__k2_diff_1=-0.00053421
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__kt1_diff_1=-0.25074
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__pclm_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__u0_diff_1=-0.0010115
*
* sky130_fd_pr__rf_nfet_g5v0d10v5_bM04, Bin 000, W = 3.01, L = 0.5
* --------------------------------------------
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__nfactor_diff_0=-0.39264
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__vsat_diff_0=-3946.4
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__vth0_diff_0=-0.024526
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__a0_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__b0_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__k2_diff_0=0.0010173
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__u0_diff_0=-0.0031271
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__b1_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__ags_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__kt1_diff_0=-0.21392
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__voff_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__pclm_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__ub_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__ua_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__rdsw_diff_0=0.0
*
* sky130_fd_pr__rf_nfet_g5v0d10v5_bM04, Bin 001, W = 5.05, L = 0.5
* --------------------------------------------
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__nfactor_diff_1=-0.41153
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__vsat_diff_1=-1841.7
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__vth0_diff_1=-0.0099998
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__a0_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__b0_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__k2_diff_1=-0.00057848
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__u0_diff_1=-0.0013993
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__b1_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__ags_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__kt1_diff_1=-0.19547
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__voff_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__pclm_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__ub_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__ua_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__rdsw_diff_1=0.0
*
* sky130_fd_pr__rf_nfet_g5v0d10v5_bM04, Bin 002, W = 7.09, L = 0.5
* --------------------------------------------
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__rdsw_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__nfactor_diff_2=-0.52459
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__vsat_diff_2=-2994.9
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__vth0_diff_2=-0.0082165
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__a0_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__b0_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__k2_diff_2=-0.0015137
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__u0_diff_2=-0.003002
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__b1_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__ags_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__kt1_diff_2=-0.18326
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__voff_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__pclm_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__ub_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__ua_diff_2=0.0
*
* sky130_fd_pr__rf_nfet_g5v0d10v5_bM10, Bin 000, W = 3.01, L = 0.5
* ---------------------------------------------
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__ags_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__ua_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__rdsw_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__k2_diff_0=0.00059498
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__kt1_diff_0=-0.11421
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__pclm_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__u0_diff_0=-0.0016449
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__b1_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__voff_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__nfactor_diff_0=-0.54235
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__ub_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__vth0_diff_0=-0.015075
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__vsat_diff_0=1100.9
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__a0_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__b0_diff_0=0.0
*
* sky130_fd_pr__rf_nfet_g5v0d10v5_bM10, Bin 001, W = 5.05, L = 0.5
* ---------------------------------------------
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__b0_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__ags_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__ua_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__rdsw_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__k2_diff_1=-0.0068059
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__kt1_diff_1=-0.12465
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__pclm_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__u0_diff_1=-0.002939
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__b1_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__voff_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__nfactor_diff_1=-0.60297
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__ub_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__vth0_diff_1=-0.012671
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__vsat_diff_1=-3862.9
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__a0_diff_1=0.0
*
* sky130_fd_pr__rf_nfet_g5v0d10v5_bM10, Bin 002, W = 7.09, L = 0.5
* ---------------------------------------------
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__a0_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__b0_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__ua_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__ags_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__rdsw_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__k2_diff_2=-0.0017173
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__kt1_diff_2=-0.14457
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__pclm_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__u0_diff_2=-0.0041054
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__b1_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__voff_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__nfactor_diff_2=-0.5182
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__ub_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__vth0_diff_2=-0.022123
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__vsat_diff_2=-5556.8
.include "sky130_fd_pr__rf_nfet_g5v0d10v5_b.pm3.spice"
