* Diode Vth

* Include SkyWater sky130 device models
.include "../../pfet_g5v0d10v5/sky130_fd_pr__pfet_g5v0d10v5__tt.corner.spice"
.include "../../../models/sky130_fd_pr__model__diode_pd2nw_11v0.model.spice"

X1 3 0 sky130_fd_pr__esd_rf_diode_pd2nw_11v0_300 area=1.0 M=1
Rd 3 4 100

* DC source for current measure
Vid 4 5
Vdd 5 0 DC 0V

.control
* Sweep Vdd from 0 to 2.0V
dc Vdd 0 2.0 0.05
* NOTE:  Internally accessed names MUST be in lowercase
wrdata sky130_fd_pr__esd_rf_diode_pd2nw_11v0_300__iv.data -Vid#branch V ( 3 )
* Find threshold
let ih=-Vid#branch[38]
let il=-Vid#branch[28]
let vh=V(3)[38]
let vl=V(3)[28]
let vth=((vl - vh ) / ( ih - il ) ) * ih vh
echo threshold voltage
print vth
quit
.endc
.end
