* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 18
.param
+  sky130_fd_pr__rf_nfet_01v8_b__toxe_mult=0.948
+  sky130_fd_pr__rf_nfet_01v8_b__rbpb_mult=0.8
+  sky130_fd_pr__rf_nfet_01v8_b__overlap_mult=0.94816
+  sky130_fd_pr__rf_nfet_01v8_b__ajunction_mult=0.7739
+  sky130_fd_pr__rf_nfet_01v8_b__pjunction_mult=0.79336
+  sky130_fd_pr__rf_nfet_01v8_b__lint_diff=1.7325e-8
+  sky130_fd_pr__rf_nfet_01v8_b__wint_diff=-3.2175e-8
+  sky130_fd_pr__rf_nfet_01v8_b__rshg_diff=-7.0
+  sky130_fd_pr__rf_nfet_01v8_b__xgw_diff=-6.425e-8
+  sky130_fd_pr__rf_nfet_01v8_b__dlc_diff=12.773e-9
+  sky130_fd_pr__rf_nfet_01v8_b__dwc_diff=0.0
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 000, W = 1.65, L = 0.15
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_bM02__ags_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__vth0_diff_0=-0.075991
+  sky130_fd_pr__rf_nfet_01v8_bM02__vsat_diff_0=-22417.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__a0_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__b0_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__k2_diff_0=0.010085
+  sky130_fd_pr__rf_nfet_01v8_bM02__nfactor_diff_0=0.27569
+  sky130_fd_pr__rf_nfet_01v8_bM02__u0_diff_0=0.00074749
+  sky130_fd_pr__rf_nfet_01v8_bM02__rdsw_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__ua_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__voff_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__b1_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__kt1_diff_0=-0.049406
+  sky130_fd_pr__rf_nfet_01v8_bM02__ub_diff_0=0.0
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 001, W = 1.65, L = 0.18
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_bM02__ags_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__vth0_diff_1=-0.039487
+  sky130_fd_pr__rf_nfet_01v8_bM02__vsat_diff_1=-19233.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__a0_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__b0_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__k2_diff_1=0.020683
+  sky130_fd_pr__rf_nfet_01v8_bM02__nfactor_diff_1=2.6612
+  sky130_fd_pr__rf_nfet_01v8_bM02__u0_diff_1=0.0011292
+  sky130_fd_pr__rf_nfet_01v8_bM02__rdsw_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__ua_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__voff_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__b1_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__kt1_diff_1=-0.15593
+  sky130_fd_pr__rf_nfet_01v8_bM02__ub_diff_1=0.0
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 002, W = 1.65, L = 0.25
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_bM02__kt1_diff_2=-0.21378
+  sky130_fd_pr__rf_nfet_01v8_bM02__ub_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__ags_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__vth0_diff_2=-0.043022
+  sky130_fd_pr__rf_nfet_01v8_bM02__vsat_diff_2=-16781.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__a0_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__b0_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__k2_diff_2=0.038033
+  sky130_fd_pr__rf_nfet_01v8_bM02__nfactor_diff_2=2.8985
+  sky130_fd_pr__rf_nfet_01v8_bM02__u0_diff_2=0.0006468
+  sky130_fd_pr__rf_nfet_01v8_bM02__rdsw_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__ua_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__voff_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__b1_diff_2=0.0
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 003, W = 3.01, L = 0.15
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_bM02__kt1_diff_3=-0.015285
+  sky130_fd_pr__rf_nfet_01v8_bM02__ub_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__ags_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__vth0_diff_3=-0.035105
+  sky130_fd_pr__rf_nfet_01v8_bM02__vsat_diff_3=-28463.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__a0_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__b0_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__k2_diff_3=0.010626
+  sky130_fd_pr__rf_nfet_01v8_bM02__nfactor_diff_3=-0.45239
+  sky130_fd_pr__rf_nfet_01v8_bM02__u0_diff_3=-0.0036794
+  sky130_fd_pr__rf_nfet_01v8_bM02__rdsw_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__ua_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__voff_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__b1_diff_3=0.0
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 004, W = 3.01, L = 0.18
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_bM02__voff_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__b1_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__rdsw_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__kt1_diff_4=-0.10619
+  sky130_fd_pr__rf_nfet_01v8_bM02__ub_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__ags_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__vth0_diff_4=-0.05182
+  sky130_fd_pr__rf_nfet_01v8_bM02__vsat_diff_4=-25171.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__a0_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__b0_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__k2_diff_4=0.030375
+  sky130_fd_pr__rf_nfet_01v8_bM02__nfactor_diff_4=1.8023
+  sky130_fd_pr__rf_nfet_01v8_bM02__u0_diff_4=-0.0033229
+  sky130_fd_pr__rf_nfet_01v8_bM02__ua_diff_4=0.0
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 005, W = 3.01, L = 0.25
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_bM02__nfactor_diff_5=2.2537
+  sky130_fd_pr__rf_nfet_01v8_bM02__ua_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__voff_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__b1_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__rdsw_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__kt1_diff_5=-0.15849
+  sky130_fd_pr__rf_nfet_01v8_bM02__ub_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__ags_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__vth0_diff_5=-0.032322
+  sky130_fd_pr__rf_nfet_01v8_bM02__vsat_diff_5=-20257.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__a0_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__b0_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__k2_diff_5=0.042979
+  sky130_fd_pr__rf_nfet_01v8_bM02__u0_diff_5=0.0011015
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 006, W = 5.05, L = 0.15
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_bM02__u0_diff_6=-0.0033456
+  sky130_fd_pr__rf_nfet_01v8_bM02__nfactor_diff_6=-0.5594
+  sky130_fd_pr__rf_nfet_01v8_bM02__ua_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__voff_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__b1_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__rdsw_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__kt1_diff_6=0.01851
+  sky130_fd_pr__rf_nfet_01v8_bM02__ub_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__ags_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__vth0_diff_6=-0.041439
+  sky130_fd_pr__rf_nfet_01v8_bM02__vsat_diff_6=-28660.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__a0_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__b0_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__k2_diff_6=0.0064952
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 007, W = 5.05, L = 0.18
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_bM02__b0_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__k2_diff_7=0.02645
+  sky130_fd_pr__rf_nfet_01v8_bM02__u0_diff_7=-0.0036669
+  sky130_fd_pr__rf_nfet_01v8_bM02__nfactor_diff_7=1.5456
+  sky130_fd_pr__rf_nfet_01v8_bM02__ua_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__b1_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__rdsw_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__voff_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__kt1_diff_7=-0.057816
+  sky130_fd_pr__rf_nfet_01v8_bM02__ub_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__ags_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__vth0_diff_7=-0.045761
+  sky130_fd_pr__rf_nfet_01v8_bM02__vsat_diff_7=-23039.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__a0_diff_7=0.0
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 008, W = 5.05, L = 0.25
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_bM02__a0_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__b0_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__k2_diff_8=0.04175
+  sky130_fd_pr__rf_nfet_01v8_bM02__u0_diff_8=-0.0010573
+  sky130_fd_pr__rf_nfet_01v8_bM02__nfactor_diff_8=1.379
+  sky130_fd_pr__rf_nfet_01v8_bM02__ua_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__b1_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__rdsw_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__voff_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__kt1_diff_8=-0.10787
+  sky130_fd_pr__rf_nfet_01v8_bM02__ub_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__ags_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM02__vth0_diff_8=-0.032973
+  sky130_fd_pr__rf_nfet_01v8_bM02__vsat_diff_8=-16043.0
*
* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 000, W = 1.65, L = 0.15
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_bM04__rdsw_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__ua_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__k2_diff_0=0.0091842
+  sky130_fd_pr__rf_nfet_01v8_bM04__u0_diff_0=-0.00070926
+  sky130_fd_pr__rf_nfet_01v8_bM04__vth0_diff_0=-0.051501
+  sky130_fd_pr__rf_nfet_01v8_bM04__voff_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__b1_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__kt1_diff_0=-0.022227
+  sky130_fd_pr__rf_nfet_01v8_bM04__nfactor_diff_0=0.0033312
+  sky130_fd_pr__rf_nfet_01v8_bM04__ub_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__vsat_diff_0=-31984.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__ags_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__a0_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__b0_diff_0=0.0
*
* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 001, W = 1.65, L = 0.18
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_bM04__b0_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__rdsw_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__ua_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__k2_diff_1=0.028977
+  sky130_fd_pr__rf_nfet_01v8_bM04__u0_diff_1=-0.0013648
+  sky130_fd_pr__rf_nfet_01v8_bM04__vth0_diff_1=-0.058125
+  sky130_fd_pr__rf_nfet_01v8_bM04__voff_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__b1_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__kt1_diff_1=-0.10064
+  sky130_fd_pr__rf_nfet_01v8_bM04__nfactor_diff_1=1.9273
+  sky130_fd_pr__rf_nfet_01v8_bM04__ub_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__vsat_diff_1=-23564.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__ags_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__a0_diff_1=0.0
*
* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 002, W = 1.65, L = 0.25
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_bM04__ags_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__a0_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__b0_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__ua_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__rdsw_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__k2_diff_2=0.042169
+  sky130_fd_pr__rf_nfet_01v8_bM04__u0_diff_2=-0.00035031
+  sky130_fd_pr__rf_nfet_01v8_bM04__vth0_diff_2=-0.046633
+  sky130_fd_pr__rf_nfet_01v8_bM04__voff_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__b1_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__kt1_diff_2=-0.15022
+  sky130_fd_pr__rf_nfet_01v8_bM04__nfactor_diff_2=1.7231
+  sky130_fd_pr__rf_nfet_01v8_bM04__ub_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__vsat_diff_2=-19030.0
*
* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 003, W = 3.01, L = 0.15
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_bM04__vsat_diff_3=-30928.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__ags_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__a0_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__b0_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__ua_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__rdsw_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__k2_diff_3=0.013856
+  sky130_fd_pr__rf_nfet_01v8_bM04__u0_diff_3=-0.0048131
+  sky130_fd_pr__rf_nfet_01v8_bM04__vth0_diff_3=-0.046817
+  sky130_fd_pr__rf_nfet_01v8_bM04__voff_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__b1_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__kt1_diff_3=-0.091215
+  sky130_fd_pr__rf_nfet_01v8_bM04__nfactor_diff_3=0.17482
+  sky130_fd_pr__rf_nfet_01v8_bM04__ub_diff_3=0.0
*
* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 004, W = 3.01, L = 0.18
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_bM04__kt1_diff_4=-0.1562
+  sky130_fd_pr__rf_nfet_01v8_bM04__nfactor_diff_4=1.7824
+  sky130_fd_pr__rf_nfet_01v8_bM04__ub_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__vsat_diff_4=-24921.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__ags_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__a0_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__b0_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__ua_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__rdsw_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__k2_diff_4=0.034977
+  sky130_fd_pr__rf_nfet_01v8_bM04__u0_diff_4=-0.0071423
+  sky130_fd_pr__rf_nfet_01v8_bM04__vth0_diff_4=-0.061148
+  sky130_fd_pr__rf_nfet_01v8_bM04__voff_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__b1_diff_4=0.0
*
* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 005, W = 3.01, L = 0.25
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_bM04__voff_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__kt1_diff_5=-0.19439
+  sky130_fd_pr__rf_nfet_01v8_bM04__nfactor_diff_5=1.8393
+  sky130_fd_pr__rf_nfet_01v8_bM04__ub_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__vsat_diff_5=-8528.2
+  sky130_fd_pr__rf_nfet_01v8_bM04__ags_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__a0_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__b0_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__ua_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__rdsw_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__k2_diff_5=0.045401
+  sky130_fd_pr__rf_nfet_01v8_bM04__u0_diff_5=-0.0043436
+  sky130_fd_pr__rf_nfet_01v8_bM04__vth0_diff_5=-0.04118
+  sky130_fd_pr__rf_nfet_01v8_bM04__b1_diff_5=0.0
*
* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 006, W = 5.05, L = 0.15
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_bM04__b1_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__voff_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__kt1_diff_6=-0.073142
+  sky130_fd_pr__rf_nfet_01v8_bM04__nfactor_diff_6=0.42429
+  sky130_fd_pr__rf_nfet_01v8_bM04__ub_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__vsat_diff_6=-29958.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__ags_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__a0_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__b0_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__ua_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__rdsw_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__k2_diff_6=0.009601
+  sky130_fd_pr__rf_nfet_01v8_bM04__u0_diff_6=-0.0033405
+  sky130_fd_pr__rf_nfet_01v8_bM04__vth0_diff_6=-0.04502
*
* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 007, W = 5.05, L = 0.18
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_bM04__u0_diff_7=-0.0060347
+  sky130_fd_pr__rf_nfet_01v8_bM04__b1_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__voff_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__kt1_diff_7=-0.11011
+  sky130_fd_pr__rf_nfet_01v8_bM04__ub_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__nfactor_diff_7=1.2003
+  sky130_fd_pr__rf_nfet_01v8_bM04__vsat_diff_7=-26996.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__ags_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__a0_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__b0_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__ua_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__rdsw_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__k2_diff_7=0.031931
+  sky130_fd_pr__rf_nfet_01v8_bM04__vth0_diff_7=-0.060436
*
* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 008, W = 5.05, L = 0.25
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_bM04__vth0_diff_8=-0.0389
+  sky130_fd_pr__rf_nfet_01v8_bM04__u0_diff_8=-0.0030982
+  sky130_fd_pr__rf_nfet_01v8_bM04__b1_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__voff_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__kt1_diff_8=-0.15194
+  sky130_fd_pr__rf_nfet_01v8_bM04__ub_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__nfactor_diff_8=1.4418
+  sky130_fd_pr__rf_nfet_01v8_bM04__vsat_diff_8=-11896.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__ags_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__a0_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__b0_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__ua_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__rdsw_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_bM04__k2_diff_8=0.044114
.include "sky130_fd_pr__rf_nfet_01v8_b.pm3.spice"
