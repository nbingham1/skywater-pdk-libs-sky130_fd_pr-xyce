* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 8
.param
+  sky130_fd_pr__rf_nfet_g5v0d10v5_b__toxe_mult=0.94
+  sky130_fd_pr__rf_nfet_g5v0d10v5_b__rbpb_mult=0.8
+  sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult=0.76246
+  sky130_fd_pr__rf_nfet_g5v0d10v5_b__ajunction_mult=0.81753
+  sky130_fd_pr__rf_nfet_g5v0d10v5_b__pjunction_mult=0.77786
+  sky130_fd_pr__rf_nfet_g5v0d10v5_b__lint_diff=1.7325e-8
+  sky130_fd_pr__rf_nfet_g5v0d10v5_b__wint_diff=-3.2175e-8
+  sky130_fd_pr__rf_nfet_g5v0d10v5_b__rshg_diff=-7.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_b__xgw_diff=-6.425e-8
+  sky130_fd_pr__rf_nfet_g5v0d10v5_b__dlc_diff=1.7325e-8
+  sky130_fd_pr__rf_nfet_g5v0d10v5_b__dwc_diff=0.0
*
* sky130_fd_pr__rf_nfet_g5v0d10v5_bM02, Bin 000, W = 3.01, L = 0.5
* --------------------------------------------
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__voff_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__ub_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__vth0_diff_0=-0.096862
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__nfactor_diff_0=-0.33307
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__ua_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__vsat_diff_0=-12674.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__a0_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__rdsw_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__b0_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__ags_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__k2_diff_0=-0.0035704
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__kt1_diff_0=-0.32676
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__pclm_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__u0_diff_0=-0.0051274
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__b1_diff_0=0.0
*
* sky130_fd_pr__rf_nfet_g5v0d10v5_bM02, Bin 001, W = 5.05, L = 0.5
* --------------------------------------------
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__b1_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__voff_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__ub_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__vth0_diff_1=-0.073057
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__nfactor_diff_1=-0.50082
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__ua_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__vsat_diff_1=-6173.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__a0_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__rdsw_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__b0_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__ags_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__k2_diff_1=-0.011741
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__kt1_diff_1=-0.32836
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__pclm_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__u0_diff_1=-0.0039209
*
* sky130_fd_pr__rf_nfet_g5v0d10v5_bM04, Bin 000, W = 3.01, L = 0.5
* --------------------------------------------
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__nfactor_diff_0=-0.37193
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__vsat_diff_0=-12970.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__vth0_diff_0=-0.10565
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__a0_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__b0_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__k2_diff_0=-0.0039729
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__u0_diff_0=-0.0051626
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__b1_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__ags_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__kt1_diff_0=-0.28517
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__voff_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__pclm_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__ub_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__ua_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__rdsw_diff_0=0.0
*
* sky130_fd_pr__rf_nfet_g5v0d10v5_bM04, Bin 001, W = 5.05, L = 0.5
* --------------------------------------------
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__nfactor_diff_1=-0.38675
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__vsat_diff_1=-8042.9
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__vth0_diff_1=-0.080494
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__a0_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__b0_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__k2_diff_1=-0.011251
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__u0_diff_1=-0.0041751
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__b1_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__ags_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__kt1_diff_1=-0.28285
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__voff_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__pclm_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__ub_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__ua_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__rdsw_diff_1=0.0
*
* sky130_fd_pr__rf_nfet_g5v0d10v5_bM04, Bin 002, W = 7.09, L = 0.5
* --------------------------------------------
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__rdsw_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__nfactor_diff_2=-0.509
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__vsat_diff_2=-9472.9
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__vth0_diff_2=-0.082655
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__a0_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__b0_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__k2_diff_2=-0.0094809
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__u0_diff_2=-0.0051933
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__b1_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__ags_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__kt1_diff_2=-0.28355
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__voff_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__pclm_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__ub_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__ua_diff_2=0.0
*
* sky130_fd_pr__rf_nfet_g5v0d10v5_bM10, Bin 000, W = 3.01, L = 0.5
* ---------------------------------------------
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__ags_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__ua_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__rdsw_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__k2_diff_0=-0.0041159
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__kt1_diff_0=-0.22789
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__pclm_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__u0_diff_0=-0.0035707
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__b1_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__voff_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__nfactor_diff_0=-0.53245
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__ub_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__vth0_diff_0=-0.096572
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__vsat_diff_0=-10255.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__a0_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__b0_diff_0=0.0
*
* sky130_fd_pr__rf_nfet_g5v0d10v5_bM10, Bin 001, W = 5.05, L = 0.5
* ---------------------------------------------
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__b0_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__ags_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__ua_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__rdsw_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__k2_diff_1=-0.016447
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__kt1_diff_1=-0.25497
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__pclm_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__u0_diff_1=-0.0053074
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__b1_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__voff_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__nfactor_diff_1=-0.58953
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__ub_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__vth0_diff_1=-0.083034
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__vsat_diff_1=-10453.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__a0_diff_1=0.0
*
* sky130_fd_pr__rf_nfet_g5v0d10v5_bM10, Bin 002, W = 7.09, L = 0.5
* ---------------------------------------------
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__a0_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__b0_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__ua_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__ags_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__rdsw_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__k2_diff_2=-0.0084536
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__kt1_diff_2=-0.24814
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__pclm_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__u0_diff_2=-0.0025043
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__b1_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__voff_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__nfactor_diff_2=-0.51293
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__ub_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__vth0_diff_2=-0.095613
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__vsat_diff_2=-15629.0
.include "sky130_fd_pr__rf_nfet_g5v0d10v5_b.pm3.spice"
