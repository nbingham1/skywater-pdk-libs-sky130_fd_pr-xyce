* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 52
.param
+  sky130_fd_pr__pfet_01v8__toxe_mult=1.052
+  sky130_fd_pr__pfet_01v8__rshp_mult=1.0
+  sky130_fd_pr__pfet_01v8__overlap_mult=1.1934
+  sky130_fd_pr__pfet_01v8__ajunction_mult=1.0909
+  sky130_fd_pr__pfet_01v8__pjunction_mult=1.096
+  sky130_fd_pr__pfet_01v8__lint_diff=-1.7325e-8
+  sky130_fd_pr__pfet_01v8__wint_diff=3.2175e-8
+  sky130_fd_pr__pfet_01v8__dlc_diff=-1.7325e-8
+  sky130_fd_pr__pfet_01v8__dwc_diff=3.2175e-8
*
* sky130_fd_pr__pfet_01v8, Bin 000, W = 1.26, L = 0.15
* -----------------------------------
+  sky130_fd_pr__pfet_01v8__agidl_diff_0=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_0=-0.15387
+  sky130_fd_pr__pfet_01v8__vsat_diff_0=12312.0
+  sky130_fd_pr__pfet_01v8__a0_diff_0=0.0
+  sky130_fd_pr__pfet_01v8__pdits_diff_0=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_0=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_0=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_0=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_0=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_0=2.6386e-11
+  sky130_fd_pr__pfet_01v8__keta_diff_0=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_0=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_0=-0.020902
+  sky130_fd_pr__pfet_01v8__vth0_diff_0=0.060085
+  sky130_fd_pr__pfet_01v8__pditsd_diff_0=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_0=7.6365e-5
+  sky130_fd_pr__pfet_01v8__b1_diff_0=0.0
+  sky130_fd_pr__pfet_01v8__cgidl_diff_0=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_0=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_0=0.061939
+  sky130_fd_pr__pfet_01v8__ags_diff_0=0.0
+  sky130_fd_pr__pfet_01v8__bgidl_diff_0=0.0
+  sky130_fd_pr__pfet_01v8__ub_diff_0=5.2476e-20
*
* sky130_fd_pr__pfet_01v8, Bin 001, W = 1.68, L = 0.15
* -----------------------------------
+  sky130_fd_pr__pfet_01v8__bgidl_diff_1=0.0
+  sky130_fd_pr__pfet_01v8__ub_diff_1=7.4573e-20
+  sky130_fd_pr__pfet_01v8__agidl_diff_1=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_1=-0.2062
+  sky130_fd_pr__pfet_01v8__vsat_diff_1=-2828.9
+  sky130_fd_pr__pfet_01v8__a0_diff_1=0.0
+  sky130_fd_pr__pfet_01v8__pdits_diff_1=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_1=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_1=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_1=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_1=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_1=3.1342e-11
+  sky130_fd_pr__pfet_01v8__keta_diff_1=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_1=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_1=-0.025224
+  sky130_fd_pr__pfet_01v8__vth0_diff_1=0.022784
+  sky130_fd_pr__pfet_01v8__pditsd_diff_1=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_1=0.00039046
+  sky130_fd_pr__pfet_01v8__b1_diff_1=0.0
+  sky130_fd_pr__pfet_01v8__cgidl_diff_1=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_1=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_1=0.054627
+  sky130_fd_pr__pfet_01v8__ags_diff_1=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 002, W = 1.0, L = 1.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__cgidl_diff_2=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_2=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_2=-0.021888
+  sky130_fd_pr__pfet_01v8__ags_diff_2=-0.067356
+  sky130_fd_pr__pfet_01v8__bgidl_diff_2=0.0
+  sky130_fd_pr__pfet_01v8__ub_diff_2=-6.194e-20
+  sky130_fd_pr__pfet_01v8__agidl_diff_2=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_2=0.050635
+  sky130_fd_pr__pfet_01v8__vsat_diff_2=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_2=0.072953
+  sky130_fd_pr__pfet_01v8__pdits_diff_2=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_2=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_2=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_2=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_2=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_2=1.6609e-11
+  sky130_fd_pr__pfet_01v8__keta_diff_2=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_2=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_2=-0.0099625
+  sky130_fd_pr__pfet_01v8__vth0_diff_2=-0.018831
+  sky130_fd_pr__pfet_01v8__pditsd_diff_2=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_2=0.00017033
+  sky130_fd_pr__pfet_01v8__b1_diff_2=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 003, W = 1.0, L = 2.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__b1_diff_3=0.0
+  sky130_fd_pr__pfet_01v8__cgidl_diff_3=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_3=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_3=-0.0075694
+  sky130_fd_pr__pfet_01v8__ags_diff_3=-0.0010758
+  sky130_fd_pr__pfet_01v8__bgidl_diff_3=0.0
+  sky130_fd_pr__pfet_01v8__ub_diff_3=-3.3431e-20
+  sky130_fd_pr__pfet_01v8__nfactor_diff_3=0.0086468
+  sky130_fd_pr__pfet_01v8__vsat_diff_3=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_3=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_3=0.0012821
+  sky130_fd_pr__pfet_01v8__pdits_diff_3=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_3=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_3=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_3=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_3=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_3=-9.0993e-14
+  sky130_fd_pr__pfet_01v8__keta_diff_3=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_3=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_3=-0.0048481
+  sky130_fd_pr__pfet_01v8__vth0_diff_3='0.0029452-0.015'
+  sky130_fd_pr__pfet_01v8__pditsd_diff_3=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_3=-0.00021812
*
* sky130_fd_pr__pfet_01v8, Bin 004, W = 1.0, L = 4.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__pditsd_diff_4=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_4=2.0928e-4
+  sky130_fd_pr__pfet_01v8__vth0_diff_4=-1.4100e-2
+  sky130_fd_pr__pfet_01v8__b1_diff_4=0.0
+  sky130_fd_pr__pfet_01v8__cgidl_diff_4=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_4=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_4=-0.0023693
+  sky130_fd_pr__pfet_01v8__ags_diff_4=-0.036839
+  sky130_fd_pr__pfet_01v8__ub_diff_4=-4.5792e-20
+  sky130_fd_pr__pfet_01v8__bgidl_diff_4=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_4=6.8951e-1
+  sky130_fd_pr__pfet_01v8__vsat_diff_4=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_4=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_4=0.040186
+  sky130_fd_pr__pfet_01v8__pdits_diff_4=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_4=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_4=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_4=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_4=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_4=6.1033e-11
+  sky130_fd_pr__pfet_01v8__keta_diff_4=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_4=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_4=-8.9077e-3
*
* sky130_fd_pr__pfet_01v8, Bin 005, W = 1.0, L = 8.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__keta_diff_5=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_5=-0.002402
+  sky130_fd_pr__pfet_01v8__pditsd_diff_5=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_5=6.7503e-5
+  sky130_fd_pr__pfet_01v8__vth0_diff_5=-0.006956
+  sky130_fd_pr__pfet_01v8__b1_diff_5=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_5=0.0032535
+  sky130_fd_pr__pfet_01v8__cgidl_diff_5=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_5=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_5=0.014051
+  sky130_fd_pr__pfet_01v8__ub_diff_5=1.8544e-20
+  sky130_fd_pr__pfet_01v8__bgidl_diff_5=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_5=-0.010861
+  sky130_fd_pr__pfet_01v8__vsat_diff_5=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_5=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_5=-0.013944
+  sky130_fd_pr__pfet_01v8__pdits_diff_5=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_5=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_5=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_5=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_5=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_5=-6.8402e-13
+  sky130_fd_pr__pfet_01v8__rdsw_diff_5=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 006, W = 1.0, L = 0.15
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__rdsw_diff_6=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_6=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_6=-0.030031
+  sky130_fd_pr__pfet_01v8__pditsd_diff_6=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_6=0.00019683
+  sky130_fd_pr__pfet_01v8__vth0_diff_6=-0.0046281
+  sky130_fd_pr__pfet_01v8__b1_diff_6=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_6=0.072202
+  sky130_fd_pr__pfet_01v8__cgidl_diff_6=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_6=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_6=0.0
+  sky130_fd_pr__pfet_01v8__ub_diff_6=4.351e-20
+  sky130_fd_pr__pfet_01v8__bgidl_diff_6=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_6=-0.39035
+  sky130_fd_pr__pfet_01v8__vsat_diff_6=22908.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_6=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_6=0.0
+  sky130_fd_pr__pfet_01v8__pdits_diff_6=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_6=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_6=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_6=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_6=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_6=1.88e-11
*
* sky130_fd_pr__pfet_01v8, Bin 007, W = 1.0, L = 0.18
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__kt1_diff_7=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_7=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_7=-1.7731e-10
+  sky130_fd_pr__pfet_01v8__rdsw_diff_7=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_7=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_7=-0.016624
+  sky130_fd_pr__pfet_01v8__pditsd_diff_7=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_7=-0.00057746
+  sky130_fd_pr__pfet_01v8__vth0_diff_7=-0.0043154
+  sky130_fd_pr__pfet_01v8__b1_diff_7=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_7=0.028739
+  sky130_fd_pr__pfet_01v8__cgidl_diff_7=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_7=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_7=0.0
+  sky130_fd_pr__pfet_01v8__ub_diff_7=1.5991e-19
+  sky130_fd_pr__pfet_01v8__bgidl_diff_7=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_7=-1.2
+  sky130_fd_pr__pfet_01v8__vsat_diff_7=100000.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_7=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_7=0.0
+  sky130_fd_pr__pfet_01v8__pdits_diff_7=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_7=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_7=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 008, W = 1.0, L = 0.25
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__pclm_diff_8=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_8=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_8=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_8=7.3685e-13
+  sky130_fd_pr__pfet_01v8__rdsw_diff_8=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_8=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_8=-0.012695
+  sky130_fd_pr__pfet_01v8__pditsd_diff_8=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_8=-0.0011527
+  sky130_fd_pr__pfet_01v8__vth0_diff_8=-0.00029106
+  sky130_fd_pr__pfet_01v8__b1_diff_8=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_8=0.039188
+  sky130_fd_pr__pfet_01v8__cgidl_diff_8=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_8=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_8=0.0
+  sky130_fd_pr__pfet_01v8__ub_diff_8=-1.754e-20
+  sky130_fd_pr__pfet_01v8__bgidl_diff_8=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_8=-0.063136
+  sky130_fd_pr__pfet_01v8__vsat_diff_8=20056.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_8=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_8=0.0
+  sky130_fd_pr__pfet_01v8__pdits_diff_8=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_8=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 009, W = 1.0, L = 0.5
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__pdits_diff_9=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_9=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_9=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_9=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_9=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_9=-2.2486e-12
+  sky130_fd_pr__pfet_01v8__rdsw_diff_9=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_9=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_9=-0.011013
+  sky130_fd_pr__pfet_01v8__pditsd_diff_9=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_9=6.5249e-5
+  sky130_fd_pr__pfet_01v8__vth0_diff_9=0.00064906
+  sky130_fd_pr__pfet_01v8__b1_diff_9=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_9=-0.0014484
+  sky130_fd_pr__pfet_01v8__cgidl_diff_9=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_9=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_9=0.0
+  sky130_fd_pr__pfet_01v8__ub_diff_9=-3.9528e-20
+  sky130_fd_pr__pfet_01v8__bgidl_diff_9=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_9=0.00087378
+  sky130_fd_pr__pfet_01v8__vsat_diff_9=1476.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_9=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_9=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 010, W = 2.0, L = 0.15
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__pditsd_diff_10=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_10=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_10=100000.0
+  sky130_fd_pr__pfet_01v8__u0_diff_10=0.00084428
+  sky130_fd_pr__pfet_01v8__vth0_diff_10=-0.0081773
+  sky130_fd_pr__pfet_01v8__cgidl_diff_10=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_10=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_10=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_10=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_10=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_10=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_10=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_10=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_10=-2.3682e-10
+  sky130_fd_pr__pfet_01v8__bgidl_diff_10=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_10=-0.31789
+  sky130_fd_pr__pfet_01v8__ub_diff_10=8.0286e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_10=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_10=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_10=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_10=-0.027023
+  sky130_fd_pr__pfet_01v8__voff_diff_10=-0.04329
+  sky130_fd_pr__pfet_01v8__a0_diff_10=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 011, W = 3.0, L = 1.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__voff_diff_11=-0.0081755
+  sky130_fd_pr__pfet_01v8__a0_diff_11=0.0058522
+  sky130_fd_pr__pfet_01v8__pditsd_diff_11=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_11=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_11=19709.0
+  sky130_fd_pr__pfet_01v8__u0_diff_11=0.00081366
+  sky130_fd_pr__pfet_01v8__vth0_diff_11=-0.028283
+  sky130_fd_pr__pfet_01v8__cgidl_diff_11=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_11=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_11=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_11=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_11=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_11=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_11=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_11=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_11=-1.8009e-11
+  sky130_fd_pr__pfet_01v8__bgidl_diff_11=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_11=-0.0078229
+  sky130_fd_pr__pfet_01v8__ub_diff_11=1.9411e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_11=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_11=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_11=-0.0033389
+  sky130_fd_pr__pfet_01v8__k2_diff_11=-0.014914
*
* sky130_fd_pr__pfet_01v8, Bin 012, W = 3.0, L = 2.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__pdits_diff_12=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_12=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_12=0.00021421
+  sky130_fd_pr__pfet_01v8__k2_diff_12=-0.011993
+  sky130_fd_pr__pfet_01v8__voff_diff_12=-0.0086635
+  sky130_fd_pr__pfet_01v8__a0_diff_12=0.00082978
+  sky130_fd_pr__pfet_01v8__pditsd_diff_12=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_12=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_12=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_12=0.0010777
+  sky130_fd_pr__pfet_01v8__vth0_diff_12=-0.021747
+  sky130_fd_pr__pfet_01v8__cgidl_diff_12=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_12=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_12=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_12=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_12=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_12=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_12=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_12=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_12=-1.7159e-13
+  sky130_fd_pr__pfet_01v8__bgidl_diff_12=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_12=0.0013748
+  sky130_fd_pr__pfet_01v8__ub_diff_12=2.2018e-19
*
* sky130_fd_pr__pfet_01v8, Bin 013, W = 3.0, L = 4.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__bgidl_diff_13=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_13=0.011813
+  sky130_fd_pr__pfet_01v8__ub_diff_13=1.6685e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_13=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_13=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_13=0.006201
+  sky130_fd_pr__pfet_01v8__k2_diff_13=-0.010269
+  sky130_fd_pr__pfet_01v8__voff_diff_13=-0.011641
+  sky130_fd_pr__pfet_01v8__a0_diff_13=-0.007114
+  sky130_fd_pr__pfet_01v8__eta0_diff_13=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_13=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_13=0.00087385
+  sky130_fd_pr__pfet_01v8__vsat_diff_13=0.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_13=-0.011971
+  sky130_fd_pr__pfet_01v8__cgidl_diff_13=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_13=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_13=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_13=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_13=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_13=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_13=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_13=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_13=-1.5741e-12
*
* sky130_fd_pr__pfet_01v8, Bin 014, W = 3.0, L = 8.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__agidl_diff_14=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_14=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_14=9.0904e-14
+  sky130_fd_pr__pfet_01v8__bgidl_diff_14=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_14=-0.0029708
+  sky130_fd_pr__pfet_01v8__ub_diff_14=8.057e-20
+  sky130_fd_pr__pfet_01v8__pdits_diff_14=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_14=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_14=-0.019832
+  sky130_fd_pr__pfet_01v8__k2_diff_14=-0.0088747
+  sky130_fd_pr__pfet_01v8__voff_diff_14=0.0026403
+  sky130_fd_pr__pfet_01v8__eta0_diff_14=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_14=0.027053
+  sky130_fd_pr__pfet_01v8__pditsd_diff_14=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_14=0.00053856
+  sky130_fd_pr__pfet_01v8__vsat_diff_14=0.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_14=-0.0067419
+  sky130_fd_pr__pfet_01v8__cgidl_diff_14=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_14=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_14=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_14=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_14=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_14=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 015, W = 3.0, L = 0.15
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__b0_diff_15=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_15=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_15=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_15=3.0205e-11
+  sky130_fd_pr__pfet_01v8__bgidl_diff_15=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_15=-0.33753
+  sky130_fd_pr__pfet_01v8__ub_diff_15=1.5966e-19
+  sky130_fd_pr__pfet_01v8__tvoff_diff_15=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_15=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_15=-0.020627
+  sky130_fd_pr__pfet_01v8__pdits_diff_15=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_15=0.042365
+  sky130_fd_pr__pfet_01v8__eta0_diff_15=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_15=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_15=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_15=0.0006404
+  sky130_fd_pr__pfet_01v8__vsat_diff_15=-7189.6
+  sky130_fd_pr__pfet_01v8__vth0_diff_15=0.029889
+  sky130_fd_pr__pfet_01v8__cgidl_diff_15=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_15=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_15=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_15=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_15=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 016, W = 3.0, L = 0.18
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__pclm_diff_16=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_16=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_16=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_16=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_16=7.9914e-12
+  sky130_fd_pr__pfet_01v8__bgidl_diff_16=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_16=-0.0046728
+  sky130_fd_pr__pfet_01v8__tvoff_diff_16=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_16=0.0
+  sky130_fd_pr__pfet_01v8__ub_diff_16=1.929e-19
+  sky130_fd_pr__pfet_01v8__k2_diff_16=-0.021859
+  sky130_fd_pr__pfet_01v8__pdits_diff_16=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_16=0.0072438
+  sky130_fd_pr__pfet_01v8__eta0_diff_16=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_16=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_16=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_16=0.00065136
+  sky130_fd_pr__pfet_01v8__vsat_diff_16=12923.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_16=0.029819
+  sky130_fd_pr__pfet_01v8__cgidl_diff_16=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_16=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_16=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_16=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 017, W = 3.0, L = 0.25
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__kt1_diff_17=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_17=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_17=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_17=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_17=0.0
+  sky130_fd_pr__pfet_01v8__bgidl_diff_17=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_17=0.049985
+  sky130_fd_pr__pfet_01v8__ua_diff_17=1.3799e-11
+  sky130_fd_pr__pfet_01v8__tvoff_diff_17=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_17=0.0
+  sky130_fd_pr__pfet_01v8__ub_diff_17=2.4784e-19
+  sky130_fd_pr__pfet_01v8__k2_diff_17=-0.013872
+  sky130_fd_pr__pfet_01v8__pdits_diff_17=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_17=0.0058902
+  sky130_fd_pr__pfet_01v8__eta0_diff_17=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_17=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_17=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_17=0.0004052
+  sky130_fd_pr__pfet_01v8__vsat_diff_17=8345.2
+  sky130_fd_pr__pfet_01v8__vth0_diff_17=-0.017331
+  sky130_fd_pr__pfet_01v8__cgidl_diff_17=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_17=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_17=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 018, W = 3.0, L = 0.5
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__rdsw_diff_18=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_18=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_18=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_18=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_18=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_18=0.0
+  sky130_fd_pr__pfet_01v8__bgidl_diff_18=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_18=0.11924
+  sky130_fd_pr__pfet_01v8__ua_diff_18=1.5351e-11
+  sky130_fd_pr__pfet_01v8__tvoff_diff_18=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_18=0.0
+  sky130_fd_pr__pfet_01v8__ub_diff_18=4.5605e-20
+  sky130_fd_pr__pfet_01v8__k2_diff_18=-0.0179
+  sky130_fd_pr__pfet_01v8__pdits_diff_18=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_18=0.0020774
+  sky130_fd_pr__pfet_01v8__eta0_diff_18=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_18=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_18=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_18=0.00039988
+  sky130_fd_pr__pfet_01v8__vsat_diff_18=-15442.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_18=-0.0143
+  sky130_fd_pr__pfet_01v8__cgidl_diff_18=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_18=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 019, W = 5.0, L = 1.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__cgidl_diff_19=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_19=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_19=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_19=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_19=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_19=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_19=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_19=0.0
+  sky130_fd_pr__pfet_01v8__bgidl_diff_19=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_19=0.0068817
+  sky130_fd_pr__pfet_01v8__ua_diff_19=9.7659e-13
+  sky130_fd_pr__pfet_01v8__tvoff_diff_19=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_19=-0.0033056
+  sky130_fd_pr__pfet_01v8__ub_diff_19=1.867e-19
+  sky130_fd_pr__pfet_01v8__k2_diff_19=-0.010736
+  sky130_fd_pr__pfet_01v8__pdits_diff_19=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_19=-0.0030155
+  sky130_fd_pr__pfet_01v8__eta0_diff_19=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_19=0.0045486
+  sky130_fd_pr__pfet_01v8__pditsd_diff_19=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_19=0.00083392
+  sky130_fd_pr__pfet_01v8__vsat_diff_19=0.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_19=-0.010897
*
* sky130_fd_pr__pfet_01v8, Bin 020, W = 5.0, L = 2.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__u0_diff_20=0.00081534
+  sky130_fd_pr__pfet_01v8__vth0_diff_20=-0.012957
+  sky130_fd_pr__pfet_01v8__cgidl_diff_20=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_20=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_20=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_20=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_20=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_20=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_20=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_20=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_20=-2.324e-12
+  sky130_fd_pr__pfet_01v8__bgidl_diff_20=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_20=0.0025067
+  sky130_fd_pr__pfet_01v8__ub_diff_20=1.7952e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_20=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_20=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_20=0.011887
+  sky130_fd_pr__pfet_01v8__k2_diff_20=-0.014239
+  sky130_fd_pr__pfet_01v8__voff_diff_20=-0.0086647
+  sky130_fd_pr__pfet_01v8__a0_diff_20=-0.014029
+  sky130_fd_pr__pfet_01v8__pditsd_diff_20=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_20=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_20=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 021, W = 5.0, L = 4.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__pditsd_diff_21=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_21=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_21=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_21=0.00084715
+  sky130_fd_pr__pfet_01v8__vth0_diff_21=-0.0084659
+  sky130_fd_pr__pfet_01v8__cgidl_diff_21=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_21=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_21=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_21=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_21=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_21=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_21=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_21=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_21=-6.6031e-13
+  sky130_fd_pr__pfet_01v8__bgidl_diff_21=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_21=0.029962
+  sky130_fd_pr__pfet_01v8__ub_diff_21=1.3354e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_21=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_21=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_21=-0.027829
+  sky130_fd_pr__pfet_01v8__k2_diff_21=-0.013535
+  sky130_fd_pr__pfet_01v8__voff_diff_21=-0.011017
+  sky130_fd_pr__pfet_01v8__a0_diff_21=0.034702
*
* sky130_fd_pr__pfet_01v8, Bin 022, W = 5.0, L = 8.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__voff_diff_22=-0.0065224
+  sky130_fd_pr__pfet_01v8__a0_diff_22=0.03716
+  sky130_fd_pr__pfet_01v8__pditsd_diff_22=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_22=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_22=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_22=0.00096429
+  sky130_fd_pr__pfet_01v8__vth0_diff_22=-0.0098069
+  sky130_fd_pr__pfet_01v8__cgidl_diff_22=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_22=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_22=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_22=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_22=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_22=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_22=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_22=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_22=1.3577e-12
+  sky130_fd_pr__pfet_01v8__bgidl_diff_22=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_22=0.019253
+  sky130_fd_pr__pfet_01v8__ub_diff_22=1.6138e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_22=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_22=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_22=-0.029663
+  sky130_fd_pr__pfet_01v8__k2_diff_22=-0.013737
*
* sky130_fd_pr__pfet_01v8, Bin 023, W = 5.0, L = 0.15
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__pdits_diff_23=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_23=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_23=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_23=-0.015836
+  sky130_fd_pr__pfet_01v8__voff_diff_23=0.031231
+  sky130_fd_pr__pfet_01v8__a0_diff_23=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_23=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_23=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_23=-1927.7
+  sky130_fd_pr__pfet_01v8__u0_diff_23=0.00075287
+  sky130_fd_pr__pfet_01v8__vth0_diff_23=0.045642
+  sky130_fd_pr__pfet_01v8__cgidl_diff_23=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_23=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_23=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_23=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_23=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_23=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_23=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_23=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_23=2.4652e-11
+  sky130_fd_pr__pfet_01v8__bgidl_diff_23=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_23=-0.12369
+  sky130_fd_pr__pfet_01v8__ub_diff_23=2.248e-19
*
* sky130_fd_pr__pfet_01v8, Bin 024, W = 5.0, L = 0.18
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__bgidl_diff_24=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_24=-0.025825
+  sky130_fd_pr__pfet_01v8__ub_diff_24=2.1321e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_24=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_24=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_24=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_24=-0.016314
+  sky130_fd_pr__pfet_01v8__voff_diff_24=0.025017
+  sky130_fd_pr__pfet_01v8__a0_diff_24=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_24=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_24=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_24=0.00061006
+  sky130_fd_pr__pfet_01v8__vsat_diff_24=7672.5
+  sky130_fd_pr__pfet_01v8__vth0_diff_24=0.021064
+  sky130_fd_pr__pfet_01v8__cgidl_diff_24=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_24=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_24=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_24=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_24=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_24=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_24=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_24=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_24=1.4456e-11
*
* sky130_fd_pr__pfet_01v8, Bin 025, W = 5.0, L = 0.25
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__agidl_diff_25=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_25=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_25=2.1966e-11
+  sky130_fd_pr__pfet_01v8__bgidl_diff_25=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_25=0.11918
+  sky130_fd_pr__pfet_01v8__ub_diff_25=3.1716e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_25=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_25=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_25=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_25=-0.012834
+  sky130_fd_pr__pfet_01v8__voff_diff_25=0.0035883
+  sky130_fd_pr__pfet_01v8__eta0_diff_25=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_25=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_25=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_25=0.00084025
+  sky130_fd_pr__pfet_01v8__vsat_diff_25=-17913.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_25=-0.016258
+  sky130_fd_pr__pfet_01v8__cgidl_diff_25=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_25=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_25=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_25=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_25=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_25=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 026, W = 5.0, L = 0.5
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__b0_diff_26=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_26=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_26=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_26=1.5671e-11
+  sky130_fd_pr__pfet_01v8__bgidl_diff_26=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_26=0.11768
+  sky130_fd_pr__pfet_01v8__ub_diff_26=2.1565e-19
+  sky130_fd_pr__pfet_01v8__tvoff_diff_26=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_26=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_26=-0.018335
+  sky130_fd_pr__pfet_01v8__pdits_diff_26=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_26=0.0034029
+  sky130_fd_pr__pfet_01v8__eta0_diff_26=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_26=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_26=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_26=0.00098147
+  sky130_fd_pr__pfet_01v8__vsat_diff_26=4431.7
+  sky130_fd_pr__pfet_01v8__vth0_diff_26=-0.018479
+  sky130_fd_pr__pfet_01v8__cgidl_diff_26=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_26=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_26=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_26=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_26=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 027, W = 7.0, L = 1.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__pclm_diff_27=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_27=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_27=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_27=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_27=-4.6987e-12
+  sky130_fd_pr__pfet_01v8__bgidl_diff_27=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_27=-0.039309
+  sky130_fd_pr__pfet_01v8__tvoff_diff_27=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_27=0.040827
+  sky130_fd_pr__pfet_01v8__ub_diff_27=1.5882e-19
+  sky130_fd_pr__pfet_01v8__k2_diff_27=-0.011414
+  sky130_fd_pr__pfet_01v8__pdits_diff_27=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_27=0.0055857
+  sky130_fd_pr__pfet_01v8__eta0_diff_27=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_27=-0.063252
+  sky130_fd_pr__pfet_01v8__pditsd_diff_27=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_27=0.00068323
+  sky130_fd_pr__pfet_01v8__vsat_diff_27=0.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_27=-0.011313
+  sky130_fd_pr__pfet_01v8__cgidl_diff_27=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_27=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_27=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_27=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 028, W = 7.0, L = 2.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__kt1_diff_28=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_28=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_28=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_28=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_28=0.0
+  sky130_fd_pr__pfet_01v8__bgidl_diff_28=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_28=-0.012968
+  sky130_fd_pr__pfet_01v8__ua_diff_28=-3.1066e-12
+  sky130_fd_pr__pfet_01v8__tvoff_diff_28=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_28=0.0090376
+  sky130_fd_pr__pfet_01v8__ub_diff_28=1.7884e-19
+  sky130_fd_pr__pfet_01v8__k2_diff_28=-0.014487
+  sky130_fd_pr__pfet_01v8__pdits_diff_28=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_28=-0.012762
+  sky130_fd_pr__pfet_01v8__eta0_diff_28=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_28=-0.010764
+  sky130_fd_pr__pfet_01v8__pditsd_diff_28=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_28=0.00093257
+  sky130_fd_pr__pfet_01v8__vsat_diff_28=0.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_28=-0.0097323
+  sky130_fd_pr__pfet_01v8__cgidl_diff_28=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_28=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_28=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 029, W = 7.0, L = 4.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__rdsw_diff_29=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_29=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_29=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_29=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_29=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_29=0.0
+  sky130_fd_pr__pfet_01v8__bgidl_diff_29=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_29=0.028777
+  sky130_fd_pr__pfet_01v8__ua_diff_29=7.4104e-13
+  sky130_fd_pr__pfet_01v8__tvoff_diff_29=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_29=-0.023155
+  sky130_fd_pr__pfet_01v8__ub_diff_29=1.8618e-19
+  sky130_fd_pr__pfet_01v8__k2_diff_29=-0.013893
+  sky130_fd_pr__pfet_01v8__pdits_diff_29=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_29=-0.013585
+  sky130_fd_pr__pfet_01v8__eta0_diff_29=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_29=0.03048
+  sky130_fd_pr__pfet_01v8__pditsd_diff_29=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_29=0.0011116
+  sky130_fd_pr__pfet_01v8__vsat_diff_29=0.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_29=-0.010286
+  sky130_fd_pr__pfet_01v8__cgidl_diff_29=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_29=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 030, W = 7.0, L = 8.0
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__cgidl_diff_30=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_30=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_30=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_30=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_30=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_30=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_30=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_30=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_30=-3.8115e-13
+  sky130_fd_pr__pfet_01v8__bgidl_diff_30=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_30=0.043698
+  sky130_fd_pr__pfet_01v8__ub_diff_30=2.3432e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_30=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_30=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_30=-0.092915
+  sky130_fd_pr__pfet_01v8__k2_diff_30=-0.014979
+  sky130_fd_pr__pfet_01v8__voff_diff_30=-0.015304
+  sky130_fd_pr__pfet_01v8__a0_diff_30=0.11379
+  sky130_fd_pr__pfet_01v8__pditsd_diff_30=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_30=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_30=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_30=0.0013354
+  sky130_fd_pr__pfet_01v8__vth0_diff_30=-0.010082
*
* sky130_fd_pr__pfet_01v8, Bin 031, W = 7.0, L = 0.15
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__u0_diff_31=0.00078003
+  sky130_fd_pr__pfet_01v8__vth0_diff_31=0.034559
+  sky130_fd_pr__pfet_01v8__cgidl_diff_31=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_31=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_31=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_31=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_31=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_31=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_31=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_31=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_31=1.8602e-11
+  sky130_fd_pr__pfet_01v8__bgidl_diff_31=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_31=-0.10955
+  sky130_fd_pr__pfet_01v8__ub_diff_31=2.5095e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_31=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_31=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_31=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_31=-0.016429
+  sky130_fd_pr__pfet_01v8__voff_diff_31=-0.0044396
+  sky130_fd_pr__pfet_01v8__a0_diff_31=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_31=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_31=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_31=-7491.4
*
* sky130_fd_pr__pfet_01v8, Bin 032, W = 7.0, L = 0.18
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__pditsd_diff_32=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_32=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_32=3750.8
+  sky130_fd_pr__pfet_01v8__u0_diff_32=0.00094023
+  sky130_fd_pr__pfet_01v8__vth0_diff_32=0.026491
+  sky130_fd_pr__pfet_01v8__cgidl_diff_32=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_32=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_32=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_32=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_32=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_32=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_32=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_32=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_32=1.7893e-11
+  sky130_fd_pr__pfet_01v8__bgidl_diff_32=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_32=-0.11453
+  sky130_fd_pr__pfet_01v8__ub_diff_32=3.1706e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_32=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_32=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_32=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_32=-0.018725
+  sky130_fd_pr__pfet_01v8__voff_diff_32=0.035851
+  sky130_fd_pr__pfet_01v8__a0_diff_32=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 033, W = 7.0, L = 0.25
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__voff_diff_33=0.017453
+  sky130_fd_pr__pfet_01v8__a0_diff_33=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_33=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_33=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_33=-20000.0
+  sky130_fd_pr__pfet_01v8__u0_diff_33=0.0010394
+  sky130_fd_pr__pfet_01v8__vth0_diff_33=-0.016275
+  sky130_fd_pr__pfet_01v8__cgidl_diff_33=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_33=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_33=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_33=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_33=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_33=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_33=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_33=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_33=6.6406e-11
+  sky130_fd_pr__pfet_01v8__bgidl_diff_33=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_33=0.39833
+  sky130_fd_pr__pfet_01v8__ub_diff_33=2.8779e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_33=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_33=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_33=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_33=-0.01555
*
* sky130_fd_pr__pfet_01v8, Bin 034, W = 7.0, L = 0.5
* ---------------------------------
+  sky130_fd_pr__pfet_01v8__pdits_diff_34=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_34=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_34=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_34=-0.020112
+  sky130_fd_pr__pfet_01v8__voff_diff_34=-0.02788
+  sky130_fd_pr__pfet_01v8__a0_diff_34=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_34=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_34=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_34=613.16
+  sky130_fd_pr__pfet_01v8__u0_diff_34=0.0011498
+  sky130_fd_pr__pfet_01v8__vth0_diff_34=-0.0068808
+  sky130_fd_pr__pfet_01v8__cgidl_diff_34=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_34=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_34=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_34=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_34=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_34=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_34=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_34=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_34=1.7924e-11
+  sky130_fd_pr__pfet_01v8__bgidl_diff_34=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_34=0.23722
+  sky130_fd_pr__pfet_01v8__ub_diff_34=1.8181e-19
*
* sky130_fd_pr__pfet_01v8, Bin 035, W = 0.42, L = 1.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__bgidl_diff_35=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_35=-0.090035
+  sky130_fd_pr__pfet_01v8__ub_diff_35=-4.0997e-20
+  sky130_fd_pr__pfet_01v8__pdits_diff_35=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_35=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_35=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_35=0.010808
+  sky130_fd_pr__pfet_01v8__voff_diff_35=0.024377
+  sky130_fd_pr__pfet_01v8__a0_diff_35=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_35=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_35=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_35=-9.3067e-5
+  sky130_fd_pr__pfet_01v8__vsat_diff_35=0.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_35=-0.048783
+  sky130_fd_pr__pfet_01v8__cgidl_diff_35=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_35=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_35=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_35=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_35=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_35=2.2388e-8
+  sky130_fd_pr__pfet_01v8__b1_diff_35=5.046e-8
+  sky130_fd_pr__pfet_01v8__agidl_diff_35=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_35=-8.4106e-12
*
* sky130_fd_pr__pfet_01v8, Bin 036, W = 0.42, L = 20.0
* -----------------------------------
+  sky130_fd_pr__pfet_01v8__agidl_diff_36=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_36=9.6435e-9
+  sky130_fd_pr__pfet_01v8__ua_diff_36=6.4807e-12
+  sky130_fd_pr__pfet_01v8__bgidl_diff_36=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_36=-0.15044
+  sky130_fd_pr__pfet_01v8__ub_diff_36=-5.9248e-21
+  sky130_fd_pr__pfet_01v8__pdits_diff_36=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_36=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_36=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_36=0.020988
+  sky130_fd_pr__pfet_01v8__voff_diff_36=0.048748
+  sky130_fd_pr__pfet_01v8__eta0_diff_36=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_36=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_36=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_36=-3.1063e-5
+  sky130_fd_pr__pfet_01v8__vsat_diff_36=19998.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_36=-0.021127
+  sky130_fd_pr__pfet_01v8__cgidl_diff_36=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_36=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_36=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_36=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_36=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_36=-7.2043e-8
*
* sky130_fd_pr__pfet_01v8, Bin 037, W = 0.42, L = 2.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__b0_diff_37=-4.3049e-8
+  sky130_fd_pr__pfet_01v8__agidl_diff_37=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_37=1.2171e-8
+  sky130_fd_pr__pfet_01v8__ua_diff_37=-5.2171e-12
+  sky130_fd_pr__pfet_01v8__bgidl_diff_37=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_37=-0.038164
+  sky130_fd_pr__pfet_01v8__ub_diff_37=-1.3408e-20
+  sky130_fd_pr__pfet_01v8__tvoff_diff_37=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_37=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_37=0.0092647
+  sky130_fd_pr__pfet_01v8__pdits_diff_37=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_37=0.017086
+  sky130_fd_pr__pfet_01v8__eta0_diff_37=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_37=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_37=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_37=-0.00014879
+  sky130_fd_pr__pfet_01v8__vsat_diff_37=0.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_37=-0.026788
+  sky130_fd_pr__pfet_01v8__cgidl_diff_37=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_37=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_37=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_37=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_37=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 038, W = 0.42, L = 4.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__pclm_diff_38=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_38=-4.5318e-8
+  sky130_fd_pr__pfet_01v8__agidl_diff_38=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_38=4.078e-9
+  sky130_fd_pr__pfet_01v8__ua_diff_38=2.0199e-12
+  sky130_fd_pr__pfet_01v8__bgidl_diff_38=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_38=-0.089367
+  sky130_fd_pr__pfet_01v8__tvoff_diff_38=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_38=0.0
+  sky130_fd_pr__pfet_01v8__ub_diff_38=4.1519e-20
+  sky130_fd_pr__pfet_01v8__k2_diff_38=0.0042115
+  sky130_fd_pr__pfet_01v8__pdits_diff_38=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_38=0.013006
+  sky130_fd_pr__pfet_01v8__eta0_diff_38=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_38=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_38=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_38=0.00083282
+  sky130_fd_pr__pfet_01v8__vsat_diff_38=0.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_38=-0.03433
+  sky130_fd_pr__pfet_01v8__cgidl_diff_38=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_38=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_38=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_38=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 039, W = 0.42, L = 8.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__kt1_diff_39=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_39=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_39=5.0e-10
+  sky130_fd_pr__pfet_01v8__agidl_diff_39=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_39=3.4812e-10
+  sky130_fd_pr__pfet_01v8__bgidl_diff_39=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_39=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_39=1.2806e-11
+  sky130_fd_pr__pfet_01v8__tvoff_diff_39=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_39=0.0
+  sky130_fd_pr__pfet_01v8__ub_diff_39=2.1839e-20
+  sky130_fd_pr__pfet_01v8__k2_diff_39=-0.0011299
+  sky130_fd_pr__pfet_01v8__pdits_diff_39=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_39=0.0063713
+  sky130_fd_pr__pfet_01v8__eta0_diff_39=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_39=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_39=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_39=0.00057373
+  sky130_fd_pr__pfet_01v8__vsat_diff_39=0.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_39=-0.05104
+  sky130_fd_pr__pfet_01v8__cgidl_diff_39=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_39=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_39=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 040, W = 0.42, L = 0.15
* -----------------------------------
+  sky130_fd_pr__pfet_01v8__rdsw_diff_40=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_40=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_40=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_40=-1.2035e-7
+  sky130_fd_pr__pfet_01v8__b1_diff_40=1.1577e-8
+  sky130_fd_pr__pfet_01v8__agidl_diff_40=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_40=2.567e-10
+  sky130_fd_pr__pfet_01v8__bgidl_diff_40=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_40=-1.2
+  sky130_fd_pr__pfet_01v8__ub_diff_40=-4.2123e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_40=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_40=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_40=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_40=-0.029691
+  sky130_fd_pr__pfet_01v8__voff_diff_40=0.1
+  sky130_fd_pr__pfet_01v8__a0_diff_40=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_40=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_40=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_40=18950.0
+  sky130_fd_pr__pfet_01v8__u0_diff_40=6.1346e-5
+  sky130_fd_pr__pfet_01v8__vth0_diff_40=-0.0035207
+  sky130_fd_pr__pfet_01v8__cgidl_diff_40=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_40=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 041, W = 0.42, L = 0.18
* -----------------------------------
+  sky130_fd_pr__pfet_01v8__cgidl_diff_41=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_41=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_41=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_41=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_41=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_41=-4.8814e-8
+  sky130_fd_pr__pfet_01v8__b1_diff_41=-6.4081e-9
+  sky130_fd_pr__pfet_01v8__agidl_diff_41=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_41=5.6529e-11
+  sky130_fd_pr__pfet_01v8__bgidl_diff_41=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_41=-0.14197
+  sky130_fd_pr__pfet_01v8__ub_diff_41=-1.8692e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_41=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_41=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_41=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_41=0.0058397
+  sky130_fd_pr__pfet_01v8__voff_diff_41=0.1
+  sky130_fd_pr__pfet_01v8__a0_diff_41=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_41=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_41=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_41=19265.0
+  sky130_fd_pr__pfet_01v8__u0_diff_41=-0.00038631
+  sky130_fd_pr__pfet_01v8__vth0_diff_41=0.087084
*
* sky130_fd_pr__pfet_01v8, Bin 042, W = 0.42, L = 0.5
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__u0_diff_42=-0.00027392
+  sky130_fd_pr__pfet_01v8__vth0_diff_42=-0.026753
+  sky130_fd_pr__pfet_01v8__cgidl_diff_42=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_42=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_42=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_42=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_42=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_42=2.2186e-8
+  sky130_fd_pr__pfet_01v8__b1_diff_42=7.1375e-10
+  sky130_fd_pr__pfet_01v8__agidl_diff_42=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_42=4.2305e-11
+  sky130_fd_pr__pfet_01v8__bgidl_diff_42=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_42=1.1011
+  sky130_fd_pr__pfet_01v8__ub_diff_42=-1.6872e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_42=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_42=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_42=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_42=0.015644
+  sky130_fd_pr__pfet_01v8__voff_diff_42=0.064149
+  sky130_fd_pr__pfet_01v8__a0_diff_42=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_42=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_42=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_42=19508.0
*
* sky130_fd_pr__pfet_01v8, Bin 043, W = 0.55, L = 1.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__pditsd_diff_43=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_43=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_43=19888.0
+  sky130_fd_pr__pfet_01v8__u0_diff_43=-2.7106e-4
+  sky130_fd_pr__pfet_01v8__vth0_diff_43='-1.7138e-02-0.030'
+  sky130_fd_pr__pfet_01v8__cgidl_diff_43=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_43=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_43=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_43=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_43=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_43=6.2533e-8
+  sky130_fd_pr__pfet_01v8__b1_diff_43=-4.8894e-10
+  sky130_fd_pr__pfet_01v8__agidl_diff_43=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_43=-1.8723e-12
+  sky130_fd_pr__pfet_01v8__bgidl_diff_43=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_43=1.6404
+  sky130_fd_pr__pfet_01v8__ub_diff_43=-6.0808e-20
+  sky130_fd_pr__pfet_01v8__pdits_diff_43=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_43=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_43=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_43=1.3978e-2
+  sky130_fd_pr__pfet_01v8__voff_diff_43=0.059032
+  sky130_fd_pr__pfet_01v8__a0_diff_43=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 044, W = 0.55, L = 2.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__voff_diff_44=-0.0021323
+  sky130_fd_pr__pfet_01v8__a0_diff_44=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_44=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_44=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_44=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_44=1.2479e-4
+  sky130_fd_pr__pfet_01v8__vth0_diff_44=-8.7235e-3
+  sky130_fd_pr__pfet_01v8__cgidl_diff_44=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_44=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_44=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_44=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_44=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_44=-2.0013e-10
+  sky130_fd_pr__pfet_01v8__b1_diff_44=7.8325e-11
+  sky130_fd_pr__pfet_01v8__agidl_diff_44=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_44=9.8128e-11
+  sky130_fd_pr__pfet_01v8__bgidl_diff_44=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_44=4.7747e-1
+  sky130_fd_pr__pfet_01v8__ub_diff_44=-1.5297e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_44=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_44=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_44=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_44=-2.1930e-3
*
* sky130_fd_pr__pfet_01v8, Bin 045, W = 0.55, L = 4.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__pdits_diff_45=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_45=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_45=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_45=0.0079096
+  sky130_fd_pr__pfet_01v8__voff_diff_45=0.012251
+  sky130_fd_pr__pfet_01v8__a0_diff_45=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_45=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_45=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_45=20024.0
+  sky130_fd_pr__pfet_01v8__u0_diff_45=0.00019001
+  sky130_fd_pr__pfet_01v8__vth0_diff_45=-0.0092871
+  sky130_fd_pr__pfet_01v8__cgidl_diff_45=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_45=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_45=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_45=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_45=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_45=-2.9576e-8
+  sky130_fd_pr__pfet_01v8__b1_diff_45=1.6484e-10
+  sky130_fd_pr__pfet_01v8__agidl_diff_45=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_45=-1.0437e-11
+  sky130_fd_pr__pfet_01v8__bgidl_diff_45=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_45=-0.013654
+  sky130_fd_pr__pfet_01v8__ub_diff_45=-1.0391e-21
*
* sky130_fd_pr__pfet_01v8, Bin 046, W = 0.55, L = 8.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__bgidl_diff_46=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_46=-0.082443
+  sky130_fd_pr__pfet_01v8__ub_diff_46=3.384e-22
+  sky130_fd_pr__pfet_01v8__pdits_diff_46=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_46=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_46=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_46=0.0055969
+  sky130_fd_pr__pfet_01v8__voff_diff_46=0.015139
+  sky130_fd_pr__pfet_01v8__a0_diff_46=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_46=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_46=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_46=-0.00011865
+  sky130_fd_pr__pfet_01v8__vsat_diff_46=0.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_46=-0.017083
+  sky130_fd_pr__pfet_01v8__cgidl_diff_46=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_46=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_46=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_46=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_46=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_46=-3.2678e-8
+  sky130_fd_pr__pfet_01v8__b1_diff_46=1.9071e-9
+  sky130_fd_pr__pfet_01v8__agidl_diff_46=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_46=5.1428e-12
*
* sky130_fd_pr__pfet_01v8, Bin 047, W = 0.55, L = 0.15
* -----------------------------------
+  sky130_fd_pr__pfet_01v8__agidl_diff_47=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_47=-1.7747e-9
+  sky130_fd_pr__pfet_01v8__ua_diff_47=4.3611e-11
+  sky130_fd_pr__pfet_01v8__bgidl_diff_47=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_47=-0.19192
+  sky130_fd_pr__pfet_01v8__ub_diff_47=-1.8536e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_47=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_47=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_47=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_47=-0.010015
+  sky130_fd_pr__pfet_01v8__voff_diff_47=0.1
+  sky130_fd_pr__pfet_01v8__eta0_diff_47=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_47=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_47=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_47=-0.00061774
+  sky130_fd_pr__pfet_01v8__vsat_diff_47=19301.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_47=0.078451
+  sky130_fd_pr__pfet_01v8__cgidl_diff_47=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_47=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_47=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_47=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_47=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_47=-1.5389e-7
*
* sky130_fd_pr__pfet_01v8, Bin 048, W = 0.55, L = 0.5
* ----------------------------------
+  sky130_fd_pr__pfet_01v8__b0_diff_48=-5.0000e-11
+  sky130_fd_pr__pfet_01v8__agidl_diff_48=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_48=-8.1786e-9
+  sky130_fd_pr__pfet_01v8__ua_diff_48=-4.5346e-10
+  sky130_fd_pr__pfet_01v8__bgidl_diff_48=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_48=5.7727e-2
+  sky130_fd_pr__pfet_01v8__ub_diff_48=3.2002e-19
+  sky130_fd_pr__pfet_01v8__tvoff_diff_48=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_48=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_48=2.2263e-2
+  sky130_fd_pr__pfet_01v8__pdits_diff_48=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_48=0.07241
+  sky130_fd_pr__pfet_01v8__eta0_diff_48=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_48=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_48=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_48=-1.5000e-3
+  sky130_fd_pr__pfet_01v8__vsat_diff_48=0.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_48='4.9887e-02-0.030'
+  sky130_fd_pr__pfet_01v8__cgidl_diff_48=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_48=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_48=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_48=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_48=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 049, W = 0.64, L = 0.15
* -----------------------------------
+  sky130_fd_pr__pfet_01v8__pclm_diff_49=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_49=-1.0445e-7
+  sky130_fd_pr__pfet_01v8__agidl_diff_49=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_49=2.6323e-8
+  sky130_fd_pr__pfet_01v8__ua_diff_49=7.0e-10
+  sky130_fd_pr__pfet_01v8__bgidl_diff_49=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_49=-1.8
+  sky130_fd_pr__pfet_01v8__tvoff_diff_49=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_49=0.0
+  sky130_fd_pr__pfet_01v8__ub_diff_49=-9.5042e-19
+  sky130_fd_pr__pfet_01v8__k2_diff_49=-0.021554
+  sky130_fd_pr__pfet_01v8__pdits_diff_49=0.0
+  sky130_fd_pr__pfet_01v8__voff_diff_49=0.0045913
+  sky130_fd_pr__pfet_01v8__eta0_diff_49=0.0
+  sky130_fd_pr__pfet_01v8__a0_diff_49=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_49=0.0
+  sky130_fd_pr__pfet_01v8__u0_diff_49=0.00099392
+  sky130_fd_pr__pfet_01v8__vsat_diff_49=19245.0
+  sky130_fd_pr__pfet_01v8__vth0_diff_49=-0.044507
+  sky130_fd_pr__pfet_01v8__cgidl_diff_49=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_49=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_49=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_49=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 050, W = 0.84, L = 0.15
* -----------------------------------
+  sky130_fd_pr__pfet_01v8__kt1_diff_50=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_50=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_50=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_50=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_50=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_50=5.0e-10
+  sky130_fd_pr__pfet_01v8__bgidl_diff_50=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_50=-1.2
+  sky130_fd_pr__pfet_01v8__ub_diff_50=-4.1858e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_50=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_50=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_50=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_50=-0.041886
+  sky130_fd_pr__pfet_01v8__voff_diff_50=0.1
+  sky130_fd_pr__pfet_01v8__a0_diff_50=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_50=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_50=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_50=24936.0
+  sky130_fd_pr__pfet_01v8__u0_diff_50=0.0013713
+  sky130_fd_pr__pfet_01v8__vth0_diff_50=-0.032263
+  sky130_fd_pr__pfet_01v8__cgidl_diff_50=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_50=0.0
+  sky130_fd_pr__pfet_01v8__rdsw_diff_50=0.0
*
* sky130_fd_pr__pfet_01v8, Bin 051, W = 1.65, L = 0.15
* -----------------------------------
+  sky130_fd_pr__pfet_01v8__rdsw_diff_51=0.0
+  sky130_fd_pr__pfet_01v8__kt1_diff_51=0.0
+  sky130_fd_pr__pfet_01v8__pclm_diff_51=0.0
+  sky130_fd_pr__pfet_01v8__b0_diff_51=0.0
+  sky130_fd_pr__pfet_01v8__b1_diff_51=0.0
+  sky130_fd_pr__pfet_01v8__agidl_diff_51=0.0
+  sky130_fd_pr__pfet_01v8__ua_diff_51=1.7718e-11
+  sky130_fd_pr__pfet_01v8__bgidl_diff_51=0.0
+  sky130_fd_pr__pfet_01v8__nfactor_diff_51=-0.37155
+  sky130_fd_pr__pfet_01v8__ub_diff_51=1.9341e-19
+  sky130_fd_pr__pfet_01v8__pdits_diff_51=0.0
+  sky130_fd_pr__pfet_01v8__tvoff_diff_51=0.0
+  sky130_fd_pr__pfet_01v8__ags_diff_51=0.0
+  sky130_fd_pr__pfet_01v8__k2_diff_51=-0.035186
+  sky130_fd_pr__pfet_01v8__voff_diff_51=0.1
+  sky130_fd_pr__pfet_01v8__a0_diff_51=0.0
+  sky130_fd_pr__pfet_01v8__pditsd_diff_51=0.0
+  sky130_fd_pr__pfet_01v8__eta0_diff_51=0.0
+  sky130_fd_pr__pfet_01v8__vsat_diff_51=15169.0
+  sky130_fd_pr__pfet_01v8__u0_diff_51=0.00075953
+  sky130_fd_pr__pfet_01v8__vth0_diff_51=0.041814
+  sky130_fd_pr__pfet_01v8__cgidl_diff_51=0.0
+  sky130_fd_pr__pfet_01v8__keta_diff_51=0.0
.include "sky130_fd_pr__pfet_01v8.pm3.spice"
