* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre=0.0
* statistics {
*   process {
*   }
*   mismatch {
*     vary sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre dist=gauss std = 1.0
*   }
* }
.subckt sky130_fd_pr__pfet_01v8_hvt d g s b
.param l=1 w=1 ad=0 as=0 pd=0 ps=0 nrd=0 nrs=0 sa=0 sb=0 sd=0 mult=1 nf=1.0
msky130_fd_pr__pfet_01v8_hvt d g s b sky130_fd_pr__pfet_01v8_hvt__model l={l} w={w} ad={ad} as={as} pd={pd} ps={ps} nrd={nrd} nrs={nrs} sa={sa} sb={sb} sd={sd} nf={nf}
.model sky130_fd_pr__pfet_01v8_hvt__model.0 pmos
* Model Flag Parameters
+  lmin=2.0e-05 lmax=0.0001 wmin=7.0e-06 wmax=0.0001
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.1148088+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+  k1=0.43657182
+  k2=0.029941288
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-0.19592208+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={2.4926776+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+  eta0=0.08
+  etab=-0.07
+  u0=0.012121798
+  ua=-2.3807897e-10
+  ub=8.2326173e-19
+  uc=-7.7670696e-11
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=200000.0
+  a0=1.4973397
+  ags=0.3863522
+  a1=0.0
+  a2=1.0
+  b0=0.0
+  b1=0.0
+  keta=-0.013169082
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=0.075489662
+  pdiblc1=0.39
+  pdiblc2=0.0036275994
+  pdiblcb=-9.5744039e-5
+  drout=0.56
+  pscbe1=746475130.0
+  pscbe2=9.5049925e-9
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=4.7923891
* Gidl Induced Drain Leakage Model Parameters
+  agidl=9.33252e-11
+  bgidl=1154444600.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-0.44169
+  kt2=-0.037961
+  at=0.0
+  ute=-0.30066
+  ua1=2.2116e-9
+  ub1=-7.9359e-19
+  uc1=1.1985e-10
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.1 pmos
* Model Flag Parameters
+  lmin=8.0e-06 lmax=2.0e-05 wmin=7.0e-06 wmax=0.0001
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.1148088+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+  k1=0.43657182
+  k2=0.029941288
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-0.19592208+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={2.4926776+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+  eta0=0.08
+  etab=-0.07
+  u0=0.012121798
+  ua=-2.3807897e-10
+  ub=8.2326173e-19
+  uc=-7.7670696e-11
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=200000.0
+  a0=1.4973397
+  ags=0.3863522
+  a1=0.0
+  a2=1.0
+  b0=0.0
+  b1=0.0
+  keta=-0.013169082
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=0.075489662
+  pdiblc1=0.39
+  pdiblc2=0.0036275994
+  pdiblcb=-9.5744039e-5
+  drout=0.56
+  pscbe1=746475130.0
+  pscbe2=9.5049925e-9
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=4.7923891
* Gidl Induced Drain Leakage Model Parameters
+  agidl=9.33252e-11
+  bgidl=1154444600.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-0.44169
+  kt2=-0.037961
+  at=0.0
+  ute=-0.30066
+  ua1=2.2116e-9
+  ub1=-7.9359e-19
+  uc1=1.1985e-10
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.2 pmos
* Model Flag Parameters
+  lmin=4.0e-06 lmax=8.0e-06 wmin=7.0e-06 wmax=0.0001
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.114178603e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-5.056396284e-09 wvth0=-6.300787338e-08 pvth0=5.055449322e-13
+  k1=4.360520813e-01 lk1=4.170133487e-09 wk1=5.196413176e-08 pk1=-4.169352504e-13
+  k2=3.027896986e-02 lk2=-2.709397187e-09 wk2=-3.376186226e-08 pk2=2.708889771e-13
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-1.957720726e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-1.203587106e-09 wvoff=-1.499792732e-08 pvoff=1.203361698e-13
+  nfactor={2.490113924e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=2.056970604e-08 wnfactor=2.563195923e-07 pnfactor=-2.056585375e-12
+  eta0=0.08
+  etab=-0.07
+  u0=1.213715227e-02 lu0=-1.231952847e-10 wu0=-1.535139349e-09 pu0=1.231722127e-14
+  ua=-2.364765199e-10 lua=-1.285729009e-17 wua=-1.602149951e-16 pua=1.285488217e-21
+  ub=8.233226294e-19 lub=-4.886274540e-28 wub=-6.088798231e-27 pub=4.885359438e-32
+  uc=-7.712301991e-11 luc=-4.394290090e-18 wuc=-5.475735247e-17 puc=4.393467127e-22
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=1.943910095e+05 lvsat=4.500384746e-02 wvsat=5.607940049e-01 pvsat=-4.499541914e-6
+  a0=1.519489998e+00 la0=-1.777233629e-07 wa0=-2.214615017e-06 pa0=1.776900788e-11
+  ags=4.068572024e-01 lags=-1.645222972e-07 wags=-2.050116227e-06 pags=1.644914855e-11
+  a1=0.0
+  a2=9.848889876e-01 la2=1.211632750e-07 wa2=1.509818428e-06 pa2=-1.211405835e-11
+  b0=0.0
+  b1=0.0
+  keta=-1.635643990e-02 lketa=2.557382988e-08 wketa=3.186760974e-07 pketa=-2.556904041e-12
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=1.175724616e-01 lpclm=-3.376521839e-07 wpclm=-4.207491829e-06 ppclm=3.375889484e-11
+  pdiblc1=0.39
+  pdiblc2=3.389781792e-03 lpdiblc2=1.908134338e-09 wpdiblc2=2.377730700e-08 ppdiblc2=-1.907776982e-13
+  pdiblcb=-1.467376427e-04 lpdiblcb=4.091481994e-10 wpdiblcb=5.098405365e-09 ppdiblcb=-4.090715741e-14
+  drout=0.56
+  pscbe1=7.505167307e+08 lpscbe1=-3.242786410e+01 wpscbe1=-4.040843795e+02 ppscbe1=3.242179101e-3
+  pscbe2=9.463130295e-09 lpscbe2=3.358822405e-16 wpscbe2=4.185436522e-15 ppscbe2=-3.358193364e-20
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=4.831958464e+00 lbeta0=-3.174855852e-07 wbeta0=-3.956195367e-06 pbeta0=3.174261265e-11
* Gidl Induced Drain Leakage Model Parameters
+  agidl=8.808287513e-11 lagidl=4.206189846e-17 wagidl=5.241343089e-16 pagidl=-4.205402110e-21
+  bgidl=1.142782668e+09 lbgidl=9.356974617e+01 wbgidl=1.165974814e+03 pbgidl=-9.355222243e-3
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.425032302e-01 lkt1=6.524968605e-09 wkt1=8.130778772e-08 pkt1=-6.523746609e-13
+  kt2=-3.814108858e-02 lkt2=1.444944301e-09 wkt2=1.800548502e-08 pkt2=-1.444673692e-13
+  at=1.982182491e+04 lat=-1.590408086e-01 wat=-1.981811268e+00 pat=1.590110234e-5
+  ute=-3.004780237e-01 lute=-1.460090468e-09 wute=-1.819422176e-08 pute=1.459817022e-13
+  ua1=2.227215228e-09 lua1=-1.252890908e-16 wua1=-1.561230316e-15 pua1=1.252656266e-20
+  ub1=-8.067459047e-19 lub1=1.055566648e-25 wub1=1.315344090e-24 pub1=-1.055368962e-29
+  uc1=1.211389359e-10 luc1=-1.034180261e-17 wuc1=-1.288694463e-16 puc1=1.033986580e-21
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.3 pmos
* Model Flag Parameters
+  lmin=2.0e-06 lmax=4.0e-06 wmin=7.0e-06 wmax=0.0001
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.123952891e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=3.427064401e-08 wvth0=6.998104626e-08 pvth0=-2.953864571e-14
+  k1=4.495243286e-01 lk1=-5.003572289e-08 wk1=-5.987291272e-07 pk1=2.201142091e-12
+  k2=2.283522063e-02 lk2=2.724067672e-08 wk2=2.580908216e-07 pk2=-9.033861336e-13
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=5.440917032e-01 ldsub=6.400735019e-08 wdsub=1.590531746e-06 pdsub=-6.399536290e-12
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-1.984452484e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=9.551989155e-09 wvoff=5.130896644e-08 pvoff=-1.464509434e-13
+  nfactor={2.496487826e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-5.075814591e-09 wnfactor=3.053533022e-06 pnfactor=-1.331122955e-11
+  eta0=7.396195640e-02 leta0=2.429418919e-08 weta0=6.036912795e-07 peta0=-2.428963937e-12
+  etab=-6.472145874e-02 letab=-2.123831633e-08 wetab=-5.277552695e-07 petab=2.123433882e-12
+  u0=1.171623015e-02 lu0=1.570393268e-09 wu0=1.997950969e-08 pu0=-7.424739945e-14
+  ua=-2.981368707e-10 lua=2.352343645e-16 wua=3.857908333e-15 pua=-1.488151135e-20
+  ub=8.397850866e-19 lub=-6.672565332e-26 wub=-1.733611397e-24 pub=6.999575319e-30
+  uc=-8.628460866e-11 luc=3.246754551e-17 wuc=1.275237878e-16 puc=-2.940651008e-22
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=2.811539150e+05 lvsat=-3.040884381e-01 wvsat=-5.996658712e-01 pvsat=1.695916064e-7
+  a0=1.153198779e+00 la0=1.296056686e-06 wa0=4.733519295e-06 pa0=-1.018694948e-11
+  ags=8.426349409e-02 lags=1.133439940e-06 wags=2.733241817e-06 pags=-2.796788209e-12
+  a1=0.0
+  a2=1.232533907e+00 la2=-8.752410119e-07 wa2=-3.019636855e-06 pa2=6.110295569e-12
+  b0=0.0
+  b1=0.0
+  keta=3.573847254e-02 lketa=-1.840310922e-07 wketa=-6.198263687e-07 pketa=1.219179401e-12
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-5.743551892e-01 lpclm=2.446332558e-06 wpclm=8.595179659e-06 ppclm=-1.775290994e-11
+  pdiblc1=0.39
+  pdiblc2=7.272018917e-03 lpdiblc2=-1.371212438e-08 wpdiblc2=-4.577618178e-08 ppdiblc2=8.907215493e-14
+  pdiblcb=6.311344871e-04 lpdiblcb=-2.720635872e-09 wpdiblcb=-4.359552385e-09 ppdiblcb=-2.852875248e-15
+  drout=0.56
+  pscbe1=6.842376061e+08 lpscbe1=2.342475193e+02 wpscbe1=8.081687591e+02 ppscbe1=-1.635345647e-3
+  pscbe2=1.012851704e-08 lpscbe2=-2.341314636e-15 wpscbe2=-6.259165504e-15 ppscbe2=8.442131502e-21
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=4.333091444e+00 lbeta0=1.689715849e-06 wbeta0=-7.088793101e-06 pbeta0=4.434668229e-11
* Gidl Induced Drain Leakage Model Parameters
+  agidl=1.730263627e-10 lagidl=-2.997099225e-16 wagidl=-9.456294062e-16 pagidl=1.708221593e-21
+  bgidl=1.334029333e+09 lbgidl=-6.759150357e+02 wbgidl=-2.331949629e+03 pbgidl=4.718746713e-3
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.275119288e-01 lkt1=-5.379283214e-08 wkt1=-3.280801412e-07 pkt1=9.948058590e-13
+  kt2=-3.544205663e-02 lkt2=-9.414664724e-09 wkt2=-1.058759390e-08 pkt2=-2.942254429e-14
+  at=-3.182745871e+05 lat=1.201296867e+00 wat=5.266760403e+00 pat=-1.326367075e-5
+  ute=-2.934644332e-01 lute=-2.967941193e-08 wute=-9.632104114e-07 pute=3.948273241e-12
+  ua1=1.926843400e-09 lua1=1.083262963e-15 wua1=7.551048735e-15 pua1=-2.413687434e-20
+  ub1=-5.658354142e-19 lub1=-8.637515121e-25 wub1=-5.146600064e-24 pub1=1.544607193e-29
+  uc1=8.410993789e-11 luc1=1.386451113e-16 wuc1=1.846585998e-15 puc1=-6.914297909e-21
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.4 pmos
* Model Flag Parameters
+  lmin=1.0e-06 lmax=2.0e-06 wmin=7.0e-06 wmax=0.0001
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.105918917e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-2.221462798e-09 wvth0=-5.437815059e-08 pvth0=2.221046763e-13
+  k1=4.209362589e-01 lk1=7.812808045e-09 wk1=8.750771989e-07 pk1=-7.811344862e-13
+  k2=3.762063953e-02 lk2=-2.677914137e-09 wk2=-3.206666877e-07 pk2=2.677412617e-13
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=6.256231254e-01 ldsub=-1.009731133e-07 wdsub=-6.561083554e-06 pdsub=1.009542030e-11
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-1.943410352e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=1.247031615e-09 wvoff=4.054992464e-08 pvoff=-1.246798071e-13
+  nfactor={2.457363595e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=7.409284747e-08 wnfactor=1.361749441e-07 pnfactor=-7.407897137e-12
+  eta0=1.028159145e-01 leta0=-3.409237215e-08 weta0=-2.281164156e-06 peta0=3.408598733e-12
+  etab=-7.525560365e-02 letab=7.773658347e-11 wetab=5.254619384e-07 petab=-7.772202496e-15
+  u0=1.248738789e-02 lu0=9.940161381e-12 wu0=-1.622155057e-08 pu0=-9.938299787e-16
+  ua=-1.795683175e-10 lua=-4.691474330e-18 wua=-3.728164909e-15 pua=4.690595711e-22
+  ub=8.021034188e-19 lub=9.523955049e-27 wub=2.196071759e-24 pub=-9.522171402e-31
+  uc=-6.956153739e-11 luc=-1.371923677e-18 wuc=-8.558592946e-17 puc=1.371666743e-22
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=1.333175302e+05 lvsat=-4.938556796e-03 wvsat=-7.598676897e-01 pvsat=4.937631903e-7
+  a0=1.792548923e+00 la0=2.318882285e-09 wa0=-1.861774140e-07 pa0=-2.318448005e-13
+  ags=6.566084449e-01 lags=-2.471151461e-08 wags=1.301161385e-07 pags=2.470688664e-12
+  a1=0.0
+  a2=0.8
+  b0=0.0
+  b1=0.0
+  keta=-5.399658834e-02 lketa=-2.450401856e-09 wketa=-1.383954429e-07 pketa=2.449942945e-13
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=6.432702753e-01 lpclm=-1.755692243e-08 wpclm=-1.045581678e-06 ppclm=1.755363437e-12
+  pdiblc1=3.865081863e-01 lpdiblc1=7.065754814e-09 wpdiblc1=3.491159731e-07 ppdiblc1=-7.064431539e-13
+  pdiblc2=5.099482136e-04 lpdiblc2=-2.893907100e-11 wpdiblc2=-3.187628269e-09 ppdiblc2=2.893365129e-15
+  pdiblcb=-6.980406594e-04 lpdiblcb=-3.102338003e-11 wpdiblcb=-7.302262240e-09 ppdiblcb=3.101756998e-15
+  drout=5.822361257e-01 ldrout=-4.499524515e-08 wdrout=-2.223196135e-06 pdrout=4.498681844e-12
+  pscbe1=800000000.0
+  pscbe2=9.004637066e-09 lpscbe2=-6.712103110e-17 wpscbe2=-5.403584421e-15 ppscbe2=6.710846068e-21
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=5.284914356e+00 lbeta0=-2.363168505e-07 wbeta0=3.150504249e-06 pbeta0=2.362725931e-11
* Gidl Induced Drain Leakage Model Parameters
+  agidl=2.717963116e-11 lagidl=-4.586144369e-18 wagidl=-3.280456684e-16 pagidl=4.585285476e-22
+  bgidl=1.009722228e+09 lbgidl=-1.967312367e+01 wbgidl=-9.720407651e+02 pbgidl=1.966943929e-3
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.571850165e-01 lkt1=6.251254213e-09 wkt1=4.724131609e-07 pkt1=-6.250083478e-13
+  kt2=-4.036298751e-02 lkt2=5.429373301e-10 wkt2=1.698432722e-09 pkt2=-5.428356488e-14
+  at=2.796575615e+05 lat=-8.630794354e-03 wat=-1.714435011e+00 pat=8.629177979e-7
+  ute=-4.037131370e-01 lute=1.934110450e-07 wute=1.054433858e-05 pute=-1.933748230e-11
+  ua1=2.271623124e-09 lua1=3.855942967e-16 wua1=1.467493875e-14 pua1=-3.855220826e-20
+  ub1=-8.850619598e-19 lub1=-2.177902124e-25 wub1=-8.274254123e-24 pub1=2.177494247e-29
+  uc1=1.581644995e-10 luc1=-1.120577515e-17 wuc1=-2.124052080e-15 puc1=1.120367653e-21
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=2.75e-6
+  sbref=2.74e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.5 pmos
* Model Flag Parameters
+  lmin=5.0e-07 lmax=1.0e-06 wmin=7.0e-06 wmax=0.0001
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.115021394e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=7.095104980e-09 wvth0=8.321207059e-08 pvth0=8.127833310e-14
+  k1=3.579582411e-01 lk1=7.227206883e-08 wk1=3.504394828e-07 pk1=-2.441572911e-13
+  k2=6.235036124e-02 lk2=-2.798927890e-08 wk2=-1.660426236e-07 pk2=1.094804396e-13
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=7.627430442e-01 ldsub=-2.413180925e-07 wdsub=1.656355342e-06 pdsub=1.684707242e-12
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-1.889349318e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-4.286223382e-09 wvoff=-2.061394003e-07 pvoff=1.278116507e-13
+  nfactor={3.159426902e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-6.444829877e-07 wnfactor=-2.089422343e-05 pnfactor=1.411713621e-11
+  eta0=1.428356295e-01 leta0=-7.505335079e-08 weta0=2.040022927e-06 peta0=-1.014222670e-12
+  etab=-1.534115370e-01 letab=8.007189753e-08 wetab=1.064026396e-06 petab=-5.590036962e-13
+  u0=1.482736636e-02 lu0=-2.385074598e-09 wu0=-1.706712528e-08 pu0=-1.283673567e-16
+  ua=2.998072472e-10 lua=-4.953419523e-16 wua=-2.889529493e-15 pua=-3.893005498e-22
+  ub=5.745995099e-19 lub=2.423787559e-25 wub=8.749830476e-25 pub=3.999435780e-31
+  uc=-6.437502238e-11 luc=-6.680425521e-18 wuc=-3.558694348e-16 puc=4.138072477e-22
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=2.073266886e+05 lvsat=-8.068841051e-02 wvsat=-9.642470812e-01 pvsat=7.029495850e-7
+  a0=1.788690308e+00 la0=6.268252188e-09 wa0=4.394503830e-06 pa0=-4.920263667e-12
+  ags=4.249774164e-01 lags=2.123674756e-07 wags=4.443726733e-06 pags=-1.944378052e-12
+  a1=0.0
+  a2=8.157189367e-01 la2=-1.608864606e-08 wa2=-1.571599283e-06 pa2=1.608563298e-12
+  b0=0.0
+  b1=0.0
+  keta=-5.291503915e-02 lketa=-3.557389080e-09 wketa=-4.921358287e-09 pketa=1.083808994e-13
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=6.659649404e-01 lpclm=-4.078536606e-08 wpclm=-8.304646574e-07 ppclm=1.535186864e-12
+  pdiblc1=3.707152219e-01 lpdiblc1=2.323016975e-08 wpdiblc1=1.928116644e-06 ppdiblc1=-2.322581920e-12
+  pdiblc2=7.725462864e-04 lpdiblc2=-2.977134504e-10 wpdiblc2=-4.925283529e-09 ppdiblc2=4.671890040e-15
+  pdiblcb=-1.722688354e-03 lpdiblcb=1.017724028e-09 wpdiblcb=1.756149983e-07 ppdiblcb=-1.841177175e-13
+  drout=5.464353249e-01 ldrout=-8.352409460e-09 wdrout=1.356213473e-06 pdrout=8.350845221e-13
+  pscbe1=7.967747491e+08 lpscbe1=3.301108767e+00 wpscbe1=3.224646842e+02 ppscbe1=-3.300490535e-4
+  pscbe2=9.254539871e-09 lpscbe2=-3.229015507e-16 wpscbe2=-1.277460621e-15 ppscbe2=2.487675836e-21
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=2.850606863e+00 lbeta0=2.255245555e-06 wbeta0=3.973130393e-05 pbeta0=-1.381392078e-11
* Gidl Induced Drain Leakage Model Parameters
+  agidl=3.709516618e-11 lagidl=-1.473489277e-17 wagidl=9.555728686e-17 pagidl=2.496245081e-23
+  bgidl=9.938475275e+08 lbgidl=-3.425049827e+00 wbgidl=6.151320216e+02 pbgidl=3.424408384e-4
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.771376627e-01 lkt1=2.667318659e-08 wkt1=1.862312216e-07 pkt1=-3.320954092e-13
+  kt2=-3.492255148e-02 lkt2=-5.025457758e-09 wkt2=-1.917599409e-07 pkt2=1.437249497e-13
+  at=4.560320206e+05 lat=-1.891535807e-01 wat=-1.383689432e+00 pat=5.243930829e-7
+  ute=-2.606946710e-01 lute=4.702878476e-08 wute=-1.753516874e-05 pute=9.402455039e-12
+  ua1=3.557243351e-09 lua1=-9.302637183e-16 wua1=-5.281107003e-14 pua1=3.052107144e-20
+  ub1=-1.694683912e-18 lub1=6.108740476e-25 wub1=3.798874602e-23 pub1=-2.557616343e-29
+  uc1=3.674054729e-10 luc1=-2.253680963e-16 wuc1=-1.140592200e-15 puc1=1.137767970e-22
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.75e-6
+  sbref=1.74e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.6 pmos
* Model Flag Parameters
+  lmin=2.5e-07 lmax=5.0e-07 wmin=7.0e-06 wmax=0.0001
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.100974240e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-2.588609424e-10 wvth0=1.890286331e-07 pvth0=2.588124630e-14
+  k1=5.180017697e-01 lk1=-1.151391931e-08 wk1=-2.314852367e-06 pk1=1.151176298e-12
+  k2=1.279318065e-03 lk2=3.982633623e-09 wk2=8.036800521e-07 pk2=-3.981887756e-13
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=2.757975244e-01 ldsub=1.360762599e-08 wdsub=7.473162720e-06 pdsub=-1.360507756e-12
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-1.999377088e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=1.473950466e-09 wvoff=3.194930362e-07 pvoff=-1.473674424e-13
+  nfactor={1.856238692e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=3.776210371e-08 wnfactor=1.328334260e-05 pnfactor=-3.775503162e-12
+  eta0=3.855132189e-02 leta0=-2.045843009e-08 weta0=-3.804419564e-06 peta0=2.045459863e-12
+  etab=-4.316676099e-04 letab=-1.612371953e-11 wetab=-6.831959278e-09 petab=1.612069988e-15
+  u0=1.002610540e-02 lu0=1.284815366e-10 wu0=7.224936343e-09 pu0=-1.284574746e-14
+  ua=-7.047379978e-10 lua=3.055757436e-17 wua=2.202701183e-15 pua=-3.055185153e-21
+  ub=1.072875408e-18 lub=-1.847864251e-26 wub=-1.890096806e-24 pub=1.847518183e-30
+  uc=-7.591114001e-11 luc=-6.410372175e-19 wuc=3.121385329e-16 puc=6.409171641e-23
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=5.135536077e+04 lvsat=9.656990086e-04 wvsat=5.629178796e-01 pvsat=-9.655181525e-8
+  a0=1.775864500e+00 la0=1.298281896e-08 wa0=-2.524477132e-06 pa0=-1.298038754e-12
+  ags=9.432344917e-01 lags=-5.895046842e-08 wags=-1.052861600e-05 pags=5.893942818e-12
+  a1=0.0
+  a2=7.685621267e-01 la2=8.598887116e-09 wa2=3.143198565e-06 pa2=-8.597276716e-13
+  b0=0.0
+  b1=0.0
+  keta=-6.437005394e-02 lketa=2.439540263e-09 wketa=6.680027668e-07 pketa=-2.439083386e-13
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=5.743452625e-01 lpclm=7.179367747e-09 wpclm=3.473075195e-06 ppclm=-7.178023195e-13
+  pdiblc1=4.412894919e-01 lpdiblc1=-1.371687206e-08 wpdiblc1=-5.127988638e-06 ppdiblc1=1.371430317e-12
+  pdiblc2=8.357800335e-04 lpdiblc2=-3.308175817e-10 wpdiblc2=-5.918046495e-08 ppdiblc2=3.307556262e-14
+  pdiblcb=2.213138396e-04 wpdiblcb=-1.760768521e-7
+  drout=4.983615438e-01 ldrout=1.681517643e-08 wdrout=6.162691258e-06 pdrout=-1.681202728e-12
+  pscbe1=8.064505017e+08 lpscbe1=-1.764341234e+00 wpscbe1=-6.449293683e+02 ppscbe1=1.764010808e-4
+  pscbe2=7.969590247e-09 lpscbe2=3.497952766e-16 wpscbe2=7.027788115e-14 ppscbe2=-3.497297669e-20
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.387867150e-09 lalpha0=-6.742242102e-16 walpha0=-1.287625958e-13 palpha0=6.740979415e-20
+  alpha1=9.178702143e-11 lalpha1=4.299658541e-18 walpha1=8.211440443e-16 palpha1=-4.298853301e-22
+  beta0=7.780920834e+00 lbeta0=-3.258724150e-07 wbeta0=-4.889006553e-05 pbeta0=3.258113856e-11
* Gidl Induced Drain Leakage Model Parameters
+  agidl=1.099332337e-11 lagidl=-1.070056021e-18 wagidl=-6.111888843e-17 pagidl=1.069855621e-22
+  bgidl=9.933155116e+08 lbgidl=-3.146528817e+00 wbgidl=6.683236567e+02 pbgidl=3.145939535e-4
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.144031702e-01 lkt1=-6.169574881e-09 wkt1=-1.626378332e-06 pkt1=6.168419443e-13
+  kt2=-4.499059075e-02 lkt2=2.453621645e-10 wkt2=1.296347928e-07 pkt2=-2.453162130e-14
+  at=9.515514865e+04 lat=-2.273207112e-04 wat=-4.254351742e-01 pat=2.272781386e-8
+  ute=-1.659350059e-01 lute=-2.579795124e-09 wute=-6.778671376e-08 pute=2.579311980e-13
+  ua1=1.668322807e-09 lua1=5.862396525e-17 wua1=1.668459405e-14 pua1=-5.861298616e-21
+  ub1=-4.176651222e-19 lub1=-5.767082899e-26 wub1=-2.187938944e-23 pub1=5.766002839e-30
+  uc1=-5.312740676e-11 luc1=-5.210723121e-18 wuc1=-1.918399979e-15 puc1=5.209747257e-22
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.25e-6
+  sbref=1.24e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.7 pmos
* Model Flag Parameters
+  lmin=1.8e-07 lmax=2.5e-07 wmin=7.0e-06 wmax=0.0001
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.107392844e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=1.496755479e-09 wvth0=8.307687725e-07 pvth0=-1.496475166e-13
+  k1=5.276136579e-01 lk1=-1.414296297e-08 wk1=-3.275861176e-06 pk1=1.414031427e-12
+  k2=-4.440728611e-03 lk2=5.547180790e-09 wk2=1.375577595e-06 pk2=-5.546141914e-13
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=2.996793189e-01 ldsub=7.075477576e-09 wdsub=5.085430533e-06 pdsub=-7.074152481e-13
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.249216801e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=8.307566293e-09 wvoff=2.817422265e-06 pvoff=-8.306010452e-13
+  nfactor={2.149668309e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-4.249676516e-08 wnfactor=-1.605412375e-05 pnfactor=4.248880636e-12
+  eta0=-3.624551230e-02 weta0=3.673863060e-6
+  etab=-4.906165764e-04 letab=1.790898647e-18 wetab=-9.381666232e-10 petab=-1.790563240e-22
+  u0=1.018777241e-02 lu0=8.426237804e-11 wu0=-8.938736216e-09 pu0=-8.424659738e-15
+  ua=-6.818848042e-10 lua=2.430676884e-17 wua=-8.219018347e-17 pua=-2.430221667e-21
+  ub=1.066803054e-18 lub=-1.681773217e-26 wub=-1.282975103e-24 pub=1.681458255e-30
+  uc=-8.064688196e-11 luc=6.542829207e-19 wuc=7.856240370e-16 puc=-6.541603866e-23
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=5.845092107e+04 lvsat=-9.750786439e-04 wvsat=-1.465052644e-01 pvsat=9.748960311e-8
+  a0=1.784699382e+00 la0=1.056630198e-08 wa0=-3.407799892e-06 pa0=-1.056432313e-12
+  ags=4.971901808e-01 lags=6.305157150e-08 wags=3.406746157e-05 pags=-6.303976320e-12
+  a1=0.0
+  a2=7.835411316e-01 la2=4.501829672e-09 wa2=1.645578594e-06 pa2=-4.500986569e-13
+  b0=0.0
+  b1=0.0
+  keta=-5.560748526e-02 lketa=4.280247753e-11 wketa=-2.080899958e-07 pketa=-4.279446148e-15
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=5.964541114e-01 lpclm=1.132155379e-09 wpclm=1.262604353e-06 ppclm=-1.131943349e-13
+  pdiblc1=3.982918272e-01 lpdiblc1=-1.956150829e-09 wpdiblc1=-8.290274333e-07 ppdiblc1=1.955784481e-13
+  pdiblc2=-2.283667944e-04 lpdiblc2=-3.975214135e-11 wpdiblc2=4.721428849e-08 ppdiblc2=3.974469657e-15
+  pdiblcb=-3.260184720e-02 lpdiblcb=8.977791007e-09 wpdiblcb=3.105624539e-06 ppdiblcb=-8.976109646e-13
+  drout=5.648438079e-01 ldrout=-1.369052466e-09 wdrout=-4.842900782e-07 pdrout=1.368796070e-13
+  pscbe1=7.999776814e+08 lpscbe1=6.104576502e-03 wpscbe1=2.231439469e+00 ppscbe1=-6.103433237e-7
+  pscbe2=1.105607251e-08 lpscbe2=-4.944193516e-16 wpscbe2=-2.383125413e-13 ppscbe2=4.943267567e-20
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=-1.354089340e-09 lalpha0=7.575572888e-17 walpha0=1.453817018e-13 palpha0=-7.574154135e-21
+  alpha1=1.075067441e-10 walpha1=-7.505338223e-16
+  beta0=6.488209541e+00 lbeta0=2.770997771e-08 wbeta0=8.035685382e-05 pbeta0=-2.770478819e-12
* Gidl Induced Drain Leakage Model Parameters
+  agidl=-4.781779655e-12 lagidl=3.244750158e-18 wagidl=1.516095978e-15 pagidl=-3.244142481e-22
+  bgidl=1.015633048e+09 lbgidl=-9.250821265e+00 wbgidl=-1.563011981e+03 pbgidl=9.249088771e-4
+  cgidl=2.452271691e+02 lcgidl=1.498146470e-05 wcgidl=5.476257301e-03 pcgidl=-1.497865897e-9
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.376999320e-01 lkt1=2.025554121e-10 wkt1=7.028615481e-07 pkt1=-2.025174775e-14
+  kt2=-4.730499624e-02 lkt2=8.783983537e-10 wkt2=3.610319975e-07 pkt2=-8.782338473e-14
+  at=9.164850018e+04 lat=7.318177772e-04 wat=-7.483600008e-02 pat=-7.316807224e-8
+  ute=-2.008893713e-01 lute=6.980922904e-09 wute=3.426995202e-06 pute=-6.979615516e-13
+  ua1=1.702500791e-09 lua1=4.927560306e-17 wua1=1.326743573e-14 pua1=-4.926637472e-21
+  ub1=-4.509980178e-19 lub1=-4.855361540e-26 wub1=-1.854672414e-23 pub1=4.854452228e-30
+  uc1=-5.803889983e-11 luc1=-3.867331536e-18 wuc1=-1.427342654e-15 puc1=3.866607262e-22
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.1e-6
+  sbref=1.1e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.8 pmos
* Model Flag Parameters
+  lmin=1.5e-07 lmax=1.8e-07 wmin=7.0e-06 wmax=0.0001
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-2.026e-8
+  vth0={-1.105259107e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=1.151247567e-09 wvth0=6.174350219e-07 pvth0=-1.151031962e-13
+  k1=5.049174235e-01 lk1=-1.031934927e-08 wk1=-1.006662787e-06 pk1=1.031741666e-12
+  k2=-7.961902617e-03 lk2=6.787025396e-09 wk2=1.727629051e-06 pk2=-6.785754322e-13
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=2.125223829e-01 ldsub=2.688633886e-08 wdsub=1.379949186e-05 pdsub=-2.688130359e-12
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-1.681342370e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-3.521270701e-09 wvoff=-2.860258534e-06 pvoff=3.520611238e-13
+  nfactor={1.841029944e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=2.201441778e-08 wnfactor=1.480393263e-05 pnfactor=-2.201029492e-12
+  eta0=-1.649621518e-01 leta0=2.838459334e-08 weta0=1.654311640e-05 peta0=-2.837927747e-12
+  etab=-1.728534057e-02 letab=3.703572536e-09 wetab=1.678219701e-06 petab=-3.702878931e-13
+  u0=1.116013687e-02 lu0=-1.231250069e-10 wu0=-1.061569718e-07 pu0=1.231019481e-14
+  ua=-3.785349030e-10 lua=-4.055761004e-17 wua=-3.041149917e-14 pua=4.055001441e-21
+  ub=8.138861775e-19 lub=3.755071443e-26 wub=2.400397594e-23 pub=-3.754368193e-30
+  uc=-7.937193976e-11 luc=4.277848370e-19 wuc=6.581536942e-16 puc=-4.277047215e-23
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=3.829933133e+04 lvsat=3.387301728e-03 wvsat=1.868276310e+00 pvsat=-3.386667355e-7
+  a0=1.830925004e+00 la0=1.255229794e-09 wa0=-8.029496334e-06 pa0=-1.254994715e-13
+  ags=8.069954653e-01 wags=3.092735154e-6
+  a1=0.0
+  a2=8.339065931e-01 la2=-6.228724624e-09 wa2=-3.390024309e-06 pa2=6.227558109e-13
+  b0=1.004609535e-24 lb0=-2.215364946e-31 wb0=-1.004421392e-28 pb0=2.214950053e-35
+  b1=0.0
+  keta=-2.368520820e-02 lketa=-6.993122774e-09 wketa=-3.399719861e-06 pketa=6.991813102e-13
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=5.660977454e-01 lpclm=7.920910003e-09 wpclm=4.297672438e-06 ppclm=-7.919426574e-13
+  pdiblc1=2.795161891e-01 lpdiblc1=2.407285587e-08 wpdiblc1=1.104631195e-05 ppdiblc1=-2.406834750e-12
+  pdiblc2=-2.940901594e-03 lpdiblc2=5.550955412e-10 wpdiblc2=3.184169681e-07 ppdiblc2=-5.549915829e-14
+  pdiblcb=1.467633113e-02 lpdiblcb=-6.980791245e-10 wpdiblcb=-1.621307868e-06 ppdiblcb=6.979483883e-14
+  drout=7.559186922e-01 ldrout=-4.361924272e-08 wdrout=-1.958820005e-05 pdrout=4.361107370e-12
+  pscbe1=8.000564266e+08 lpscbe1=-1.075040191e-02 wpscbe1=-5.641606431e+00 ppscbe1=1.074838857e-6
+  pscbe2=8.737652132e-09 lpscbe2=-2.446007639e-17 wpscbe2=-6.513923068e-15 ppscbe2=2.445549551e-21
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=-5.214169504e-09 lalpha0=9.333084731e-16 walpha0=5.313174266e-13 palpha0=-9.331336831e-20
+  alpha1=1.075067441e-10 walpha1=-7.505338223e-16
+  beta0=5.510089875e+00 lbeta0=2.457195374e-07 wbeta0=1.781505022e-04 pbeta0=-2.456735190e-11
* Gidl Induced Drain Leakage Model Parameters
+  agidl=5.883420111e-11 lagidl=-1.051281235e-17 wagidl=-4.844310699e-15 pagidl=1.051084351e-21
+  bgidl=9.162852767e+08 lbgidl=1.188462923e+01 wbgidl=8.369904522e+03 pbgidl=-1.188240348e-3
+  cgidl=4.384786632e+02 lcgidl=-2.638295492e-05 wcgidl=-1.384527290e-02 pcgidl=2.637801392e-9
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-1.106e-8
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-6.225285935e-01 lkt1=4.097789125e-08 wkt1=1.918226622e-05 pkt1=-4.097021691e-12
+  kt2=-3.702604909e-02 lkt2=-1.314942569e-09 wkt2=-6.666702137e-07 pkt2=1.314696306e-13
+  at=9.131749198e+04 lat=8.659403532e-04 wat=-4.174137884e-02 pat=-8.657781798e-8
+  ute=-2.204873539e-01 lute=1.188578564e-08 wute=5.386426433e-06 pute=-1.188355967e-12
+  ua1=1.961436525e-09 lua1=-3.708920197e-18 wua1=-1.262128838e-14 pua1=3.708225590e-22
+  ub1=-7.429927856e-19 lub1=1.178139341e-26 wub1=1.064728416e-23 pub1=-1.177918700e-30
+  uc1=-9.002829368e-11 luc1=2.863931878e-18 wuc1=1.770997633e-15 puc1=-2.863395521e-22
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.04e-6
+  sbref=1.04e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.9 pmos
* Model Flag Parameters
+  lmin=2.0e-05 lmax=0.0001 wmin=5.0e-06 wmax=7.0e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.108040143e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-6.770249470e-07 wvth0=-4.725383895e-08 pvth0=4.726495306e-12
+  k1=4.350800323e-01 lk1=1.492138590e-07 wk1=1.041457585e-08 pk1=-1.041702536e-12
+  k2=3.245888784e-02 lk2=-2.518191977e-07 wk2=-1.757604925e-08 pk2=1.758018314e-12
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.203899246e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=2.447359946e-06 wvoff=1.708166785e-07 pvoff=-1.708568546e-11
+  nfactor={1.471364250e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.021553563e-04 wnfactor=7.130066296e-06 pnfactor=-7.131743287e-10
+  eta0=0.08
+  etab=-0.07
+  u0=1.025053831e-02 lu0=1.871699809e-07 wu0=1.306377287e-08 pu0=-1.306684547e-12
+  ua=-6.044964943e-10 lua=3.665037057e-14 wua=2.558060403e-15 pua=-2.558662059e-19
+  ub=9.838180906e-19 lub=-1.605941235e-23 wub=-1.120887625e-24 pub=1.121151258e-28
+  uc=-7.884651350e-11 luc=1.176094057e-16 wuc=8.208701822e-18 puc=-8.210632509e-22
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=1.752591599e+05 lvsat=2.474665916e+00 wvsat=1.727225343e-01 pvsat=-1.727631587e-5
+  a0=1.600990900e+00 la0=-1.036755791e-05 wa0=-7.236172224e-07 pa0=7.237874172e-11
+  ags=4.711848020e-01 lags=-8.485255459e-06 wags=-5.922394688e-07 pags=5.923787635e-11
+  a1=0.0
+  a2=8.753179845e-01 la2=1.247013383e-05 wa2=8.703692509e-07 pa2=-8.705739617e-11
+  b0=0.0
+  b1=0.0
+  keta=-3.618630516e-02 lketa=2.302263681e-06 wketa=1.606894956e-07 pketa=-1.607272898e-11
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=1.378101959e-01 lpclm=-6.233519171e-06 wpclm=-4.350765985e-07 ppclm=4.351789285e-11
+  pdiblc1=0.39
+  pdiblc2=1.469910110e-03 lpdiblc2=2.158196778e-07 wpdiblc2=1.506341582e-08 ppdiblc2=-1.506695874e-12
+  pdiblcb=-1.946926328e-03 lpdiblcb=1.851617687e-07 wpdiblcb=1.292360708e-08 ppdiblcb=-1.292664672e-12
+  drout=0.56
+  pscbe1=7.291872065e+08 lpscbe1=1.729198958e+03 wpscbe1=1.206916960e+02 ppscbe1=-1.207200827e-2
+  pscbe2=9.567285369e-09 lpscbe2=-6.230752035e-15 wpscbe2=-4.348834626e-16 ppscbe2=4.349857472e-20
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=3.334896019e-10 lalpha0=-2.335445187e-14 walpha0=-1.630054420e-15 palpha0=1.630437809e-19
+  alpha1=3.783247579e-11 lalpha1=6.218214601e-15 walpha1=4.340083961e-16 palpha1=-4.341104748e-20
+  beta0=3.808922830e+00 lbeta0=9.836975816e-05 wbeta0=6.865845536e-06 pbeta0=-6.867460383e-10
* Gidl Induced Drain Leakage Model Parameters
+  agidl=3.522350450e-10 lagidl=-2.589707406e-14 wagidl=-1.807520051e-15 pagidl=1.807945180e-19
+  bgidl=1.338946403e+09 lbgidl=-1.845451982e+04 wbgidl=-1.288057274e+03 pbgidl=1.288360225e-1
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-3.731169628e-01 lkt1=-6.858916555e-06 wkt1=-4.787270243e-07 pkt1=4.788396209e-11
+  kt2=-0.037961
+  at=0.0
+  ute=-3.318731997e-01 lute=3.122054108e-06 wute=2.179078374e-07 pute=-2.179590893e-11
+  ua1=2.2116e-9
+  ub1=-8.727419866e-19 lub1=7.917060318e-24 wub1=5.525815480e-25 pub1=-5.527115152e-29
+  uc1=1.1985e-10
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.10 pmos
* Model Flag Parameters
+  lmin=8.0e-06 lmax=2.0e-05 wmin=5.0e-06 wmax=7.0e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.141851628e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} wvth0=1.887933349e-7
+  k1=4.425319618e-01 wk1=-4.160937079e-8
+  k2=1.988271753e-02 wk2=7.022161639e-8
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-9.816566307e-02+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} wvoff=-6.824641364e-7
+  nfactor={6.573132387e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} wnfactor=-2.848676475e-5
+  eta0=0.08
+  etab=-0.07
+  u0=1.959804469e-02 wu0=-5.219371167e-8
+  ua=1.225869524e-09 wua=-1.022022263e-14
+  ub=1.817906574e-19 wub=4.478284038e-24
+  uc=-7.297295053e-11 wuc=-3.279623891e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=2.988471162e+05 wvsat=-6.900786050e-1
+  a0=1.083221901e+00 wa0=2.891068992e-6
+  ags=4.742037597e-02 wags=2.366175253e-6
+  a1=0.0
+  a2=1.498092294e+00 wa2=-3.477387596e-6
+  b0=0.0
+  b1=0.0
+  keta=7.879166481e-02 wketa=-6.420029868e-7
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-1.734996623e-01 wpclm=1.738262198e-6
+  pdiblc1=0.39
+  pdiblc2=1.224821871e-02 wpdiblc2=-6.018288821e-8
+  pdiblcb=7.300287385e-03 wpdiblcb=-5.163370709e-8
+  drout=0.56
+  pscbe1=8.155455970e+08 wpscbe1=-4.821997172e+2
+  pscbe2=9.256113705e-09 wpscbe2=1.737490562e-15
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=-8.328613627e-10 walpha0=6.512558911e-15
+  alpha1=3.483780043e-10 walpha1=-1.733994407e-15
+  beta0=8.721633390e+00 wbeta0=-2.743112314e-5
* Gidl Induced Drain Leakage Model Parameters
+  agidl=-9.410976986e-10 wagidl=7.221587618e-15
+  bgidl=4.173042635e+08 wbgidl=5.146177192e+3
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-7.156599600e-01 wkt1=1.912658811e-6
+  kt2=-0.037961
+  at=0.0
+  ute=-1.759538555e-01 wute=-8.706075150e-7
+  ua1=2.2116e-9
+  ub1=-4.773539471e-19 wub1=-2.207729902e-24
+  uc1=1.1985e-10
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.11 pmos
* Model Flag Parameters
+  lmin=4.0e-06 lmax=8.0e-06 wmin=5.0e-06 wmax=7.0e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.160019051e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=1.457666885e-07 wvth0=2.570167638e-07 pvth0=-5.473920468e-13
+  k1=6.144773880e-01 lk1=-1.379607566e-06 wk1=-1.193671465e-06 pk1=9.243593257e-12
+  k2=-5.621731060e-02 lk2=6.105900977e-07 wk2=5.700921986e-07 pk2=-4.010721614e-12
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-5.937388203e-02+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-3.112466310e-07 wvoff=-9.672307962e-07 pvoff=2.284830991e-12
+  nfactor={7.767593117e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-9.583779558e-06 wnfactor=-3.658719813e-05 pnfactor=6.499398922e-11
+  eta0=0.08
+  etab=-0.07
+  u0=2.238056326e-02 lu0=-2.232559345e-08 wu0=-7.304717772e-08 pu0=1.673182019e-13
+  ua=1.894261785e-09 lua=-5.362858678e-15 wua=-1.503547866e-14 pua=3.863530310e-20
+  ub=-1.720579305e-19 lub=2.839111222e-24 wub=6.942933634e-24 pub=-1.977516533e-29
+  uc=-1.288959178e-10 luc=4.486990467e-16 wuc=3.066833303e-16 puc=-2.723821113e-21
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=3.971096976e+05 lvsat=-7.884117866e-01 wvsat=-8.544402961e-01 pvsat=1.318759316e-6
+  a0=3.067434025e-01 la0=6.230090765e-06 wa0=6.251898837e-06 pa0=-2.696568547e-11
+  ags=-5.501474967e-01 lags=4.794597777e-06 wags=4.630993883e-06 pags=-1.817181758e-11
+  a1=0.0
+  a2=2.200289370e+00 la2=-5.634092286e-06 wa2=-6.975222231e-06 pa2=2.806494615e-11
+  b0=0.0
+  b1=0.0
+  keta=2.232542109e-01 lketa=-1.159098128e-06 wketa=-1.354111030e-06 pketa=5.713613127e-12
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-9.845529400e-01 lpclm=6.507502195e-06 wpclm=3.486745377e-06 ppclm=-1.402898976e-11
+  pdiblc1=0.39
+  pdiblc2=2.342852582e-02 lpdiblc2=-8.970541773e-08 wpdiblc2=-1.161186156e-07 ppdiblc2=4.488014276e-13
+  pdiblcb=9.707473309e-03 lpdiblcb=-1.931410440e-08 wpdiblcb=-6.369652163e-08 ppdiblcb=9.678623372e-14
+  drout=0.56
+  pscbe1=6.407730835e+08 lpscbe1=1.402290758e+03 wpscbe1=3.620658722e+02 ppscbe1=-6.773981842e-3
+  pscbe2=9.820213557e-09 lpscbe2=-4.526066447e-15 wpscbe2=1.692541139e-15 ppscbe2=3.606525906e-22
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=-1.771207950e-09 lalpha0=7.528842612e-15 walpha0=1.306341167e-14 palpha0=-5.256089812e-20
+  alpha1=5.982164713e-10 lalpha1=-2.004583936e-15 walpha1=-3.478184701e-15 palpha1=1.399454571e-20
+  beta0=1.378049567e+01 lbeta0=-4.058988271e-05 wbeta0=-6.642836763e-05 pbeta0=3.128951711e-10
* Gidl Induced Drain Leakage Model Parameters
+  agidl=2.298854359e-07 lagidl=-1.852041309e-12 wagidl=-1.603753692e-12 pagidl=1.292569238e-17
+  bgidl=2.404173694e+09 lbgidl=-1.594168661e+04 wbgidl=-7.640139039e+03 pbgidl=1.025912640e-1
+  cgidl=300.0
+  egidl=6.255642992e-01 legidl=-4.216875666e-06 wegidl=-3.669107326e-06 pegidl=2.943915601e-11
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-9.382687104e-01 lkt1=1.786105761e-06 wkt1=3.542381453e-06 pkt1=-1.307611222e-11
+  kt2=-4.609668255e-02 lkt2=6.527681166e-08 wkt2=7.354565048e-08 pkt2=-5.900949975e-13
+  at=-4.630730766e+05 lat=3.715476092e+00 wat=1.389409387e+00 pat=-1.114795401e-5
+  ute=-2.292033449e+00 lute=1.697840694e-05 wute=1.388539591e-05 pute=-1.183950886e-10
+  ua1=-4.901446257e-09 lua1=5.707166891e-14 wua1=4.820589451e-14 pua1=-3.867809587e-19
+  ub1=4.303583952e-18 lub1=-3.835995085e-23 wub1=-3.436125865e-23 pub1=2.579844810e-28
+  uc1=-8.842320168e-11 luc1=1.671084199e-15 wuc1=1.334140837e-15 puc1=-1.070450569e-20
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.12 pmos
* Model Flag Parameters
+  lmin=2.0e-06 lmax=4.0e-06 wmin=5.0e-06 wmax=7.0e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.134456185e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=4.291398427e-08 wvth0=1.433074019e-07 pvth0=-8.988015505e-14
+  k1=1.429845038e-01 lk1=5.174534834e-07 wk1=1.541308769e-06 pk1=-1.760654415e-12
+  k2=1.466794375e-01 lk2=-2.057690260e-07 wk2=-6.064993416e-07 pk2=7.233179800e-13
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=1.299735799e+00 ldsub=-2.976341784e-06 wdsub=-3.684825225e-06 pdsub=1.482596799e-11
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-1.098479640e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-1.081631528e-07 wvoff=-5.672127749e-07 pvoff=6.753504815e-13
+  nfactor={7.137640313e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-7.049151852e-06 wnfactor=-2.934761488e-05 pnfactor=3.586538125e-11
+  eta0=3.607690274e-01 leta0=-1.129679797e-06 weta0=-1.398586895e-06 peta0=5.627242343e-12
+  etab=-3.154521686e-01 letab=9.875817095e-07 wetab=1.222664015e-06 petab=-4.919413117e-12
+  u0=1.941129734e-02 lu0=-1.037869260e-08 wu0=-3.374184738e-08 pu0=9.172419175e-15
+  ua=9.921942718e-10 lua=-1.733371996e-15 wua=-5.150244343e-15 pua=-1.138134892e-21
+  ub=3.725872679e-19 lub=6.477203732e-25 wub=1.528023653e-24 pub=2.011833279e-30
+  uc=7.102714358e-11 luc=-3.556953894e-16 wuc=-9.707123435e-16 puc=2.415805928e-21
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=2.932006537e+05 lvsat=-3.703316704e-01 wvsat=-6.837674309e-01 pvsat=6.320536295e-7
+  a0=1.768526805e+00 la0=3.485760090e-07 wa0=4.377469720e-07 pa0=-3.572329161e-12
+  ags=5.602000646e-01 lags=3.270921579e-07 wags=-5.894008362e-07 pags=2.832544986e-12
+  a1=0.0
+  a2=0.8
+  b0=0.0
+  b1=0.0
+  keta=-8.725057452e-02 lketa=9.022408639e-08 wketa=2.387936218e-07 pketa=-6.954705980e-13
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=2.722919430e-01 lpclm=1.450561671e-06 wpclm=2.684505740e-06 ppclm=-1.080116254e-11
+  pdiblc1=0.39
+  pdiblc2=1.960393394e-03 lpdiblc2=-3.327957534e-09 wpdiblc2=-8.694279241e-09 ppdiblc2=1.657746168e-14
+  pdiblcb=1.142406264e-02 lpdiblcb=-2.622083591e-08 wpdiblcb=-7.970791951e-08 ppdiblcb=1.612084133e-13
+  drout=0.56
+  pscbe1=1.179482796e+09 lpscbe1=-7.652185455e+02 wpscbe1=-2.649272619e+03 ppscbe1=5.342198806e-3
+  pscbe2=9.703400594e-09 lpscbe2=-4.056067152e-15 wpscbe2=-3.291311963e-15 ppscbe2=2.041328523e-20
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=2.793180190e-03 lalpha0=-1.123841596e-08 walpha0=-1.949994995e-08 palpha0=7.845843863e-14
+  alpha1=-1.519925879e-10 lalpha1=1.013897217e-15 walpha1=1.759228798e-15 palpha1=-7.078292255e-21
+  beta0=6.804964503e+01 lbeta0=-2.589428905e-04 wbeta0=-4.519113846e-04 pbeta0=1.863893800e-9
* Gidl Induced Drain Leakage Model Parameters
+  agidl=-4.633915017e-07 lagidl=9.373723153e-13 wagidl=3.235324431e-12 pagidl=-6.544435233e-18
+  bgidl=-3.303865438e+09 lbgidl=7.024722995e+03 wbgidl=3.004645528e+04 pbgidl=-4.904150195e-2
+  cgidl=300.0
+  egidl=-9.511285983e-01 legidl=2.126979741e-06 wegidl=7.338214652e-06 pegidl=-1.484902411e-11
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-5.884023036e-01 lkt1=3.784112758e-07 wkt1=7.951393273e-07 pkt1=-2.022528578e-12
+  kt2=-2.952864375e-02 lkt2=-1.385023815e-09 wkt2=-5.187073766e-08 pkt2=-8.547965154e-14
+  at=7.388026946e+05 lat=-1.120295111e+00 wat=-2.112983625e+00 pat=2.943994325e-6
+  ute=4.296448953e+00 lute=-9.530483774e-06 wute=-3.300664422e-05 pute=7.027597271e-11
+  ua1=1.782893089e-08 lua1=-3.438445814e-14 wua1=-1.034657494e-13 pua1=2.234729339e-19
+  ub1=-1.144795964e-17 lub1=2.501669983e-23 wub1=7.082446911e-23 pub1=-1.652323984e-28
+  uc1=1.050703613e-09 luc1=-2.912215323e-15 wuc1=-4.901467363e-15 puc1=1.438458862e-20
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.13 pmos
* Model Flag Parameters
+  lmin=1.0e-06 lmax=2.0e-06 wmin=5.0e-06 wmax=7.0e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.147383735e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=6.907314031e-08 wvth0=2.350990250e-07 pvth0=-2.756223402e-13
+  k1=3.433298593e-01 lk1=1.120506495e-07 wk1=1.416868583e-06 pk1=-1.508847210e-12
+  k2=6.036842326e-02 lk2=-3.111696260e-08 wk2=-4.794751533e-07 pk2=4.662819945e-13
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=-1.743627175e+00 ldsub=3.181964063e-06 wdsub=9.979297233e-06 pdsub=-1.282365709e-11
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-1.224464768e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-8.266981023e-08 wvoff=-4.613655432e-07 pvoff=4.611664912e-13
+  nfactor={6.174456768e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-5.100130685e-06 wnfactor=-2.581386354e-05 pnfactor=2.871476473e-11
+  eta0=-6.240498191e-01 leta0=8.631208350e-07 weta0=2.793283238e-06 peta0=-2.855090708e-12
+  etab=-4.212735909e-01 letab=1.201713474e-06 wetab=2.941107624e-06 petab=-8.396718130e-12
+  u0=1.839616428e-02 lu0=-8.324550562e-09 wu0=-5.747232573e-08 pu0=5.719151674e-14
+  ua=1.002142239e-09 lua=-1.753501906e-15 wua=-1.197800773e-14 pua=1.267798087e-20
+  ub=2.892245920e-19 lub=8.164064151e-25 wub=5.776618352e-24 pub=-6.585283066e-30
+  uc=-1.279682227e-10 luc=4.697571425e-17 wuc=3.221670276e-16 puc=-2.003613367e-22
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=9.123788455e+04 lvsat=3.834403225e-02 wvsat=-4.660982375e-01 pvsat=1.915956632e-7
+  a0=6.167977963e-01 la0=2.679122693e-06 wa0=8.022061005e-06 pa0=-1.891934029e-11
+  ags=-5.841844931e-01 lags=2.642777198e-06 wags=8.792429134e-06 pags=-1.615177560e-11
+  a1=0.0
+  a2=0.8
+  b0=0.0
+  b1=0.0
+  keta=2.879347863e-02 lketa=-1.445933760e-07 wketa=-7.163754193e-07 pketa=1.237333060e-12
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=9.620445228e-01 lpclm=5.483353120e-08 wpclm=-3.271031406e-06 ppclm=1.249985990e-12
+  pdiblc1=5.363964344e-01 lpdiblc1=-2.962361130e-07 wpdiblc1=-6.972946565e-07 ppdiblc1=1.410989683e-12
+  pdiblc2=1.988241060e-04 lpdiblc2=2.366131510e-10 wpdiblc2=-1.015586249e-09 ppdiblc2=1.039472837e-15
+  pdiblcb=-6.204607727e-02 lpdiblcb=1.224474616e-07 wpdiblcb=4.209850680e-07 ppdiblcb=-8.519538608e-13
+  drout=-1.104146720e-01 ldrout=1.356597497e-06 wdrout=2.612387485e-06 pdrout=-5.286218323e-12
+  pscbe1=8.026724822e+08 lpscbe1=-2.735338973e+00 wpscbe1=-1.865732510e+01 ppscbe1=1.909614538e-5
+  pscbe2=6.529375979e-09 lpscbe2=2.366635137e-15 wpscbe2=1.187688650e-14 ppscbe2=-1.027986772e-20
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=-5.550299118e-03 lalpha0=5.644781295e-09 walpha0=3.874814853e-08 palpha0=-3.940775360e-14
+  alpha1=3.490636000e-10 walpha1=-1.738780737e-15
+  beta0=-8.113928659e+01 lbeta0=4.294389638e-05 wbeta0=6.065013585e-04 pbeta0=-2.778255543e-10
* Gidl Induced Drain Leakage Model Parameters
+  agidl=-2.009077583e-10 lagidl=9.688451904e-17 wagidl=1.264294437e-15 pagidl=-2.498657537e-22
+  bgidl=-1.176512912e+08 lbgidl=5.773549445e+02 wbgidl=6.898460421e+03 pbgidl=-2.201071407e-3
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-3.539925581e-01 lkt1=-9.592153241e-08 wkt1=-2.480014596e-07 pkt1=8.828766663e-14
+  kt2=-1.126756896e-02 lkt2=-3.833667387e-08 wkt2=-2.014245981e-07 pkt2=2.171455762e-13
+  at=1.295071730e+05 lat=1.126265628e-01 wat=-6.661943077e-01 pat=1.638720589e-8
+  ute=5.476944561e-01 lute=-1.944804073e-06 wute=3.902303394e-06 pute=-4.410020968e-12
+  ua1=3.005299628e-09 lua1=-4.388543816e-15 wua1=9.552943513e-15 pua1=-5.222651534e-21
+  ub1=-5.867946440e-20 lub1=1.970263605e-24 wub1=-1.404345510e-23 pub1=6.499543617e-30
+  uc1=-6.996263011e-10 luc1=6.296122650e-16 wuc1=3.864418818e-15 puc1=-3.353357387e-21
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=2.75e-6
+  sbref=2.74e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.14 pmos
* Model Flag Parameters
+  lmin=5.0e-07 lmax=1.0e-06 wmin=5.0e-06 wmax=7.0e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.068182483e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-1.199092545e-08 wvth0=-2.437831103e-07 pvth0=2.145231029e-13
+  k1=4.353011249e-01 lk1=1.791621972e-08 wk1=-1.895122268e-07 pk1=1.353156763e-13
+  k2=4.430925493e-02 lk2=-1.468008263e-08 wk2=-4.009275317e-08 pk2=1.656532028e-14
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=1.747613553e+00 ldsub=-3.913906473e-07 wdsub=-5.219293564e-06 pdsub=2.732404567e-12
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.920389307e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=9.091145818e-08 wvoff=5.136576603e-07 pvoff=-5.367892580e-13
+  nfactor={-4.807464680e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=6.140085555e-06 wnfactor=3.472481369e-05 pnfactor=-3.324778219e-11
+  eta0=5.400164911e-01 leta0=-3.283243147e-07 weta0=-7.328047011e-07 peta0=7.539308192e-13
+  etab=1.544391921e+00 letab=-8.101844905e-07 wetab=-1.078880134e-05 petab=5.656118298e-12
+  u0=1.010599306e-02 lu0=1.606054853e-10 wu0=1.589406592e-08 pu0=-1.790045244e-14
+  ua=-6.837859573e-10 lua=-2.792067872e-17 wua=3.977202205e-15 pua=-3.652495599e-21
+  ub=1.060784935e-18 lub=2.669897289e-26 wub=-2.519209648e-24 pub=1.905662808e-30
+  uc=-1.416036312e-10 luc=6.093182749e-17 wuc=1.832844893e-16 puc=-5.821228112e-23
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=1.800908601e+05 lvsat=-5.259876526e-02 wvsat=-7.741063545e-01 pvsat=5.068481311e-7
+  a0=5.968410662e+00 la0=-2.798360107e-06 wa0=-2.478526085e-05 pa0=1.465960977e-11
+  ags=3.542808022e+00 lags=-1.581282181e-06 wags=-1.732269678e-05 pags=1.057757808e-11
+  a1=0.0
+  a2=1.506618902e-01 la2=6.646105421e-07 wa2=3.071344854e-06 pa2=-3.143582885e-12
+  b0=0.0
+  b1=0.0
+  keta=-2.019073207e-01 lketa=9.153350609e-08 wketa=1.035234285e-06 pketa=-5.554745045e-13
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=4.746650055e-01 lpclm=5.536762148e-07 wpclm=5.050522222e-07 ppclm=-2.614911125e-12
+  pdiblc1=1.335071147e+00 lpdiblc1=-1.113695655e-06 wpdiblc1=-4.804314372e-06 ppdiblc1=5.614606503e-12
+  pdiblc2=2.229783483e-03 lpdiblc2=-1.842114391e-09 wpdiblc2=-1.509865277e-08 ppdiblc2=1.545377308e-14
+  pdiblcb=1.440601212e-01 lpdiblcb=-8.850635464e-08 wpdiblcb=-8.421344480e-07 ppdiblcb=4.408742262e-13
+  drout=8.452348106e-01 ldrout=3.784711386e-07 wdrout=-7.297870108e-07 pdrout=-1.865435883e-12
+  pscbe1=9.499741653e+08 lpscbe1=-1.535015577e+02 wpscbe1=-7.470621103e+02 ppscbe1=7.646330112e-4
+  pscbe2=8.944163672e-09 lpscbe2=-1.049483623e-16 wpscbe2=8.893600510e-16 ppscbe2=9.660853449e-22
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=-7.212182280e-05 lalpha0=3.775726902e-11 walpha0=5.035027602e-10 palpha0=-2.635937650e-16
+  alpha1=6.098431517e-10 lalpha1=-2.669130868e-16 walpha1=-3.559353720e-15 palpha1=1.863392859e-21
+  beta0=-8.949517053e+01 lbeta0=5.149631071e-05 wbeta0=6.844222940e-04 pbeta0=-3.575791902e-10
* Gidl Induced Drain Leakage Model Parameters
+  agidl=-2.813310970e-10 lagidl=1.791994147e-16 wagidl=2.318577642e-15 pagidl=-1.328945700e-21
+  bgidl=-3.220042723e+08 lbgidl=7.865143077e+02 wbgidl=9.801451348e+03 pbgidl=-5.172340680e-3
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.055005721e-01 lkt1=-4.320204996e-08 wkt1=-3.138867931e-07 pkt1=1.557226232e-13
+  kt2=-6.961287253e-02 lkt2=2.138091124e-08 wkt2=5.042262617e-08 pkt2=-4.062509483e-14
+  at=4.762483034e+05 lat=-2.422699190e-01 wat=-1.524824801e+00 pat=8.952126882e-7
+  ute=-2.653281287e+00 lute=1.331458619e-06 wute=-8.318707952e-07 pute=4.355009987e-13
+  ua1=-5.460209246e-09 lua1=4.276073828e-15 wua1=1.014221930e-14 pua1=-5.825787089e-21
+  ub1=6.418331373e-18 lub1=-4.659086527e-24 wub1=-1.865042043e-23 pub1=1.121486477e-29
+  uc1=6.646302350e-11 luc1=-1.544954805e-16 wuc1=9.603688960e-16 puc1=-3.810042108e-22
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.75e-6
+  sbref=1.74e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.15 pmos
* Model Flag Parameters
+  lmin=2.5e-07 lmax=5.0e-07 wmin=5.0e-06 wmax=7.0e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.117628391e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=1.389499659e-08 wvth0=3.052957900e-07 pvth0=-7.293068296e-14
+  k1=2.016500546e-01 lk1=1.402372280e-07 wk1=-1.063149961e-07 pk1=9.176026209e-14
+  k2=1.041084279e-01 lk2=-4.598614566e-08 wk2=8.580206686e-08 pk2=-4.934313591e-14
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=1.450662923e+00 ldsub=-2.359310533e-07 wdsub=-7.288921885e-07 pdsub=3.815896385e-13
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.691331461e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=7.891982185e-08 wvoff=8.025652050e-07 pvoff=-6.880381358e-13
+  nfactor={1.373776762e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-3.568714456e-06 wnfactor=-6.966484259e-05 pnfactor=2.140229067e-11
+  eta0=-7.185587252e-01 leta0=3.305649825e-07 weta0=1.481171609e-06 peta0=-4.051300584e-13
+  etab=-5.973928727e-03 letab=1.463038985e-09 wetab=3.186007308e-08 petab=-8.714367188e-15
+  u0=1.668495700e-02 lu0=-3.283613714e-09 wu0=-3.926231784e-08 pu0=1.097501758e-14
+  ua=6.662618483e-10 lua=-7.346977059e-16 wua=-7.368621654e-15 pua=2.287270107e-21
+  ub=3.314638057e-19 lub=4.085131705e-25 wub=3.285899257e-24 pub=-1.133427806e-30
+  uc=-8.980501514e-11 luc=3.381421602e-17 wuc=4.091354543e-16 puc=-1.764497783e-22
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=8.302198147e+04 lvsat=-1.781265927e-03 wvsat=3.418445872e-01 pvsat=-7.737450586e-8
+  a0=3.465333115e-01 la0=1.448051234e-07 wa0=7.454072674e-06 pa0=-2.218326117e-12
+  ags=-2.364577166e+00 lags=1.511352112e-06 wags=1.256411690e-05 pags=-5.068766621e-12
+  a1=0.0
+  a2=2.098676220e+00 la2=-3.552139196e-07 wa2=-6.142689708e-06 pa2=1.680148489e-12
+  b0=0.0
+  b1=0.0
+  keta=3.954702331e-03 lketa=-1.623938021e-08 wketa=1.910090590e-07 pketa=-1.135057141e-13
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=2.188538802e+00 lpclm=-3.435709955e-07 wpclm=-7.796048969e-06 ppclm=1.730881370e-12
+  pdiblc1=-2.214995844e+00 lpdiblc1=7.448354167e-07 wpdiblc1=1.341626181e-05 ppdiblc1=-3.924229537e-12
+  pdiblc2=-1.180361173e-02 lpdiblc2=5.504648669e-09 wpdiblc2=2.905856684e-08 ppdiblc2=-7.663414525e-15
+  pdiblcb=-0.025
+  drout=2.347480820e+00 ldrout=-4.079846921e-07 wdrout=-6.746513369e-06 pdrout=1.284440700e-12
+  pscbe1=5.000516694e+08 lpscbe1=8.204186738e+01 wpscbe1=1.494124221e+03 ppscbe1=-4.086728568e-4
+  pscbe2=1.721592081e-08 lpscbe2=-4.435378661e-15 wpscbe2=5.726732475e-15 ppscbe2=-1.566375867e-21
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=-5.978582246e-08 lalpha0=3.135142577e-14 walpha0=2.983075706e-13 palpha0=-1.561699794e-19
+  alpha1=4.819035035e-10 lalpha1=-1.999341221e-16 walpha1=-1.902365229e-15 palpha1=9.959262445e-22
+  beta0=-2.097858390e+01 lbeta0=1.562650728e-05 wbeta0=1.518878596e-04 pbeta0=-7.878676314e-11
* Gidl Induced Drain Leakage Model Parameters
+  agidl=1.785666659e-11 lagidl=2.256863670e-17 wagidl=-1.090337543e-16 pagidl=-5.804258153e-23
+  bgidl=9.928906596e+08 lbgidl=9.814051296e+01 wbgidl=6.712896636e+02 pbgidl=-3.925184352e-4
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-9.981063204e-01 lkt1=2.670389114e-07 wkt1=2.448612126e-06 pkt1=-1.290500811e-12
+  kt2=-2.320283450e-02 lkt2=-2.915671869e-09 wkt2=-2.247145986e-08 pkt2=-2.463582914e-15
+  at=-4.305382275e+04 lat=2.959513005e-02 wat=5.394392480e-01 pat=-1.854708266e-7
+  ute=-1.129708342e-01 lute=1.555291119e-09 wute=-4.375440026e-07 pute=2.290630362e-13
+  ua1=4.427681481e-09 lua1=-9.004347262e-16 wua1=-2.579239406e-15 pua1=8.341509731e-22
+  ub1=-4.781699273e-18 lub1=1.204353517e-24 wub1=8.587119985e-24 pub1=-3.044532387e-30
+  uc1=-3.387452462e-10 luc1=5.763915280e-17 wuc1=7.557584605e-17 puc1=8.220264674e-23
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.25e-6
+  sbref=1.24e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.16 pmos
* Model Flag Parameters
+  lmin=1.8e-07 lmax=2.5e-07 wmin=5.0e-06 wmax=7.0e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.033836982e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-9.023629721e-09 wvth0=3.172552923e-07 pvth0=-7.620184602e-14
+  k1=-7.179019438e-01 lk1=3.917530906e-07 wk1=5.419422020e-06 pk1=-1.419639327e-12
+  k2=4.547178430e-01 lk2=-1.418848329e-07 wk2=-1.829933285e-06 pk2=4.746487974e-13
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=3.805262131e+00 ldsub=-8.799610287e-07 wdsub=-1.938799660e-05 pdsub=5.485227876e-12
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={1.043886688e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-2.802173631e-07 wvoff=-6.040474065e-06 pvoff=1.183669965e-12
+  nfactor={-5.454426575e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.680734499e-06 wnfactor=3.703213095e-05 pnfactor=-7.781465534e-12
+  eta0=0.49
+  etab=-6.249996955e-04 letab=-8.327678673e-17 wetab=-1.516614237e-15 petab=4.148243259e-22
+  u0=2.502012850e-02 lu0=-5.563449825e-09 wu0=-1.124874485e-07 pu0=3.100355533e-14
+  ua=3.876963028e-09 lua=-1.612888693e-15 wua=-3.190874691e-14 pua=8.999485166e-21
+  ub=-2.324599821e-18 lub=1.134999694e-24 wub=2.239333083e-23 pub=-6.359692490e-30
+  uc=6.986948201e-11 luc=-9.859952434e-18 wuc=-2.651716403e-16 puc=7.986698224e-24
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=1.603207695e+05 lvsat=-2.292403043e-02 wvsat=-8.576863849e-01 pvsat=2.507212056e-7
+  a0=3.791647055e+00 la0=-7.975023878e-07 wa0=-1.741884749e-05 pa0=4.584915005e-12
+  ags=8.717042371e+00 lags=-1.519692463e-06 wags=-2.331756237e-05 pags=4.745590294e-12
+  a1=0.0
+  a2=-1.020052651e-01 la2=2.467164801e-07 wa2=7.827818858e-06 pa2=-2.141065014e-12
+  b0=0.0
+  b1=0.0
+  keta=3.845372347e-01 lketa=-1.203363145e-07 wketa=-3.280860005e-06 pketa=8.361199123e-13
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=1.233741352e+00 lpclm=-8.241479669e-08 wpclm=-3.186471212e-06 ppclm=4.700696623e-13
+  pdiblc1=9.266435940e-01 lpdiblc1=-1.144658025e-07 wpdiblc1=-4.517594829e-06 ppdiblc1=9.810389291e-13
+  pdiblc2=5.066555978e-03 lpdiblc2=8.903203988e-10 wpdiblc2=1.024899240e-08 ppdiblc2=-2.518619725e-15
+  pdiblcb=9.241277873e-01 lpdiblcb=-2.596054324e-07 wpdiblcb=-3.573565269e-06 ppdiblcb=9.774415725e-13
+  drout=4.483823127e-01 ldrout=1.114567316e-07 wdrout=3.287592976e-07 pdrout=-6.507878801e-13
+  pscbe1=7.984893667e+08 lpscbe1=4.131884139e-01 wpscbe1=1.262176923e+01 ppscbe1=-3.452306319e-6
+  pscbe2=-6.562293270e-08 lpscbe2=1.822270455e-14 wpscbe2=2.970044507e-13 ppscbe2=-8.123665736e-20
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=6.771515431e-08 lalpha0=-3.522641393e-15 walpha0=-3.368094750e-13 palpha0=1.754723494e-20
+  alpha1=-2.490636000e-10 walpha1=1.738780737e-15
+  beta0=4.308361785e+01 lbeta0=-1.895786144e-06 wbeta0=-1.751256456e-04 pbeta0=1.065797080e-11
* Gidl Induced Drain Leakage Model Parameters
+  agidl=3.921827450e-10 lagidl=-7.981703225e-17 wagidl=-1.255221343e-15 pagidl=2.554626477e-22
+  bgidl=-1.259459367e+09 lbgidl=7.142032922e+02 wbgidl=1.432002699e+04 pbgidl=-4.125721069e-3
+  cgidl=2.846936635e+03 lcgidl=-6.966381084e-04 wcgidl=-1.268698415e-02 pcgidl=3.470143904e-9
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=1.097822318e+00 lkt1=-3.062394899e-07 wkt1=-1.001703694e-05 pkt1=2.119103523e-12
+  kt2=2.202787940e-02 lkt2=-1.528717674e-08 wkt2=-1.229996659e-07 pkt2=2.503289201e-14
+  at=1.223245529e+05 lat=-1.563916325e-02 wat=-2.889938678e-01 pat=4.112219920e-8
+  ute=-1.648664105e+00 lute=4.215981144e-07 wute=1.353430441e-05 pute=-3.592516942e-12
+  ua1=3.339621791e-09 lua1=-6.028286398e-16 wua1=1.838248726e-15 pua1=-3.741203808e-22
+  ub1=-1.683862502e-18 lub1=3.570332029e-25 wub1=-9.939761842e-24 pub1=2.022940330e-30
+  uc1=-4.730024479e-10 luc1=9.436118261e-17 wuc1=1.469630745e-15 puc1=-2.990992492e-22
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.1e-6
+  sbref=1.1e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.17 pmos
* Model Flag Parameters
+  lmin=1.5e-07 lmax=1.8e-07 wmin=5.0e-06 wmax=7.0e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-2.026e-8
+  vth0={-7.864545651e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-6.433014291e-08 wvth0=-1.608226198e-06 pvth0=3.420402017e-13
+  k1=2.231797383e+00 lk1=-2.259915185e-07 wk1=-1.306248150e-05 pk1=2.537407742e-12
+  k2=-9.539460961e-02 lk2=-3.242565707e-08 wk2=2.338020560e-06 pk2=-4.048210300e-13
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=-5.967321931e+00 ldsub=1.201586175e-06 wdsub=5.694266594e-05 pdsub=-1.088902943e-11
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-5.979759371e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=5.843966186e-08 wvoff=1.405832923e-07 pvoff=-8.050499979e-14
+  nfactor={4.225575476e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-3.135080126e-07 wnfactor=-1.843228334e-06 pnfactor=1.413438568e-13
+  eta0=2.203525186e+00 leta0=-3.778665741e-07 weta0=8.062068554e-09 peta0=-1.777847358e-15
+  etab=3.717098228e-01 letab=-8.210727516e-08 wetab=-1.037461342e-06 petab=2.287809752e-13
+  u0=-6.278305794e-02 lu0=1.333419458e-08 wu0=4.100605836e-07 pu0=-8.163901365e-14
+  ua=-2.252968576e-08 lua=4.075581108e-15 wua=1.242317101e-13 pua=-2.468088254e-20
+  ub=1.746716558e-17 lub=-3.134674032e-24 wub=-9.225709729e-23 pub=1.839179561e-29
+  uc=3.276711830e-10 luc=-6.753398413e-17 wuc=-2.183525062e-15 puc=4.316891226e-22
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=-8.000231262e+04 lvsat=2.815717426e-02 wvsat=2.694172265e+00 pvsat=-5.115919530e-7
+  a0=-8.390843776e-01 la0=1.570512336e-07 wa0=1.061056540e-05 pa0=-1.213153751e-12
+  ags=1.25
+  a1=0.0
+  a2=3.288562375e+00 la2=-4.803632994e-07 wa2=-2.052664399e-05 pa2=3.932818242e-12
+  b0=-4.671434337e-23 lb0=1.030144700e-29 wb0=2.326968506e-28 pb0=-5.131430950e-35
+  b1=0.0
+  keta=-1.167657057e+00 lketa=2.119018935e-07 wketa=4.586658775e-06 pketa=-8.289843380e-13
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=2.086595653e+00 lpclm=-2.773703249e-07 wpclm=-6.317337034e-06 ppclm=1.199753053e-12
+  pdiblc1=1.111623739e+00 lpdiblc1=-1.648189381e-07 wpdiblc1=5.237142818e-06 ppdiblc1=-1.088129758e-12
+  pdiblc2=3.731465057e-02 lpdiblc2=-6.146661070e-09 wpdiblc2=3.738200889e-08 ppdiblc2=-8.712372510e-15
+  pdiblcb=-2.846287229e+00 lpdiblcb=5.501616779e-07 wpdiblcb=1.835185693e-05 ppdiblcb=-3.775906959e-12
+  drout=9.707988652e-01 ldrout=5.563400195e-09 wdrout=-2.108833699e-05 pdrout=4.017749963e-12
+  pscbe1=8.038192380e+08 lpscbe1=-7.276412232e-01 wpscbe1=-3.191081606e+01 ppscbe1=6.079648675e-6
+  pscbe2=1.134615031e-07 lpscbe2=-1.974685501e-14 wpscbe2=-7.376196116e-13 ppscbe2=1.401329531e-19
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=2.472088819e-07 lalpha0=-4.339884400e-14 walpha0=-1.230916555e-12 palpha0=2.161814465e-19
+  alpha1=-2.490636000e-10 walpha1=1.738780737e-15
+  beta0=6.936154958e+01 lbeta0=-7.848950426e-06 wbeta0=-2.676139056e-04 pbeta0=3.194374086e-11
* Gidl Induced Drain Leakage Model Parameters
+  agidl=-2.216786569e-09 lagidl=4.888457742e-16 wagidl=1.104241687e-14 pagidl=-2.435073767e-21
+  bgidl=5.108109374e+09 lbgidl=-6.303156553e+02 wbgidl=-2.089435968e+04 pbgidl=3.295134517e-3
+  cgidl=-6.139257841e+03 lcgidl=1.226807404e-03 wcgidl=3.207569478e-02 pcgidl=-6.111061370e-9
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-1.106e-8
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=2.991625939e+00 lkt1=-7.494412103e-07 wkt1=-6.049129622e-06 pkt1=1.421109051e-12
+  kt2=-9.113273842e-01 lkt2=1.892593900e-07 wkt2=5.437065217e-06 pkt2=-1.198981622e-12
+  at=4.886346092e+05 lat=-9.772419421e-02 wat=-2.815520245e+00 pat=6.017067279e-7
+  ute=5.965435931e+00 lute=-1.222247188e-06 wute=-3.779918659e-05 pute=7.427462005e-12
+  ua1=-3.402938721e-09 lua1=8.336866039e-16 wua1=2.482887432e-14 pua1=-5.475263366e-21
+  ub1=5.647008248e-18 lub1=-1.229747476e-24 wub1=-3.396305113e-23 pub1=7.489532036e-30
+  uc1=5.840870338e-10 luc1=-1.308662122e-16 wuc1=-2.935184827e-15 puc1=6.472669581e-22
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.04e-6
+  sbref=1.04e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.18 pmos
* Model Flag Parameters
+  lmin=2.0e-05 lmax=0.0001 wmin=3.0e-06 wmax=5.0e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.105023953e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-9.787147949e-07 wvth0=-6.227829712e-08 pvth0=6.229294498e-12
+  k1=4.564604659e-01 lk1=-1.989332367e-06 wk1=-9.608717931e-08 pk1=9.610977902e-12
+  k2=2.113654736e-02 lk2=8.806811518e-07 wk2=3.882360836e-08 pk2=-3.883273967e-12
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-1.671824734e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-2.874636618e-06 wvoff=-9.422410853e-08 pvoff=9.424627004e-12
+  nfactor={3.519822945e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.027386930e-04 wnfactor=-3.073863648e-06 pnfactor=3.074586621e-10
+  eta0=0.08
+  etab=-0.07
+  u0=1.252691333e-02 lu0=-4.052106141e-08 wu0=1.724529722e-09 pu0=-1.724935331e-13
+  ua=1.115990911e-10 lua=-3.497603054e-14 wua=-1.009006486e-15 pua=1.009243805e-19
+  ub=4.293807568e-19 lub=3.939736140e-23 wub=1.640915542e-24 pub=-1.641301485e-28
+  uc=-8.825926672e-11 luc=1.059106115e-15 wuc=5.509618585e-17 puc=-5.510914448e-21
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=2.099335431e+05 lvsat=-9.935879494e-1
+  a0=1.456412825e+00 la0=4.093650064e-06 wa0=-3.434505911e-09 pa0=3.435313707e-13
+  ags=3.081280271e-01 lags=7.824257127e-06 wags=2.199906785e-07 pags=-2.200424203e-11
+  a1=0.0
+  a2=1.050046297e+00 la2=-5.006807030e-6
+  b0=0.0
+  b1=0.0
+  keta=3.107433122e-03 lketa=-1.628034336e-06 wketa=-3.504330271e-08 pketa=3.505154490e-12
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=7.444511586e-03 lpclm=6.806115463e-06 wpclm=2.143103346e-07 ppclm=-2.143607404e-11
+  pdiblc1=0.39
+  pdiblc2=4.538916351e-03 lpdiblc2=-9.115312932e-08 wpdiblc2=-2.241390338e-10 ppdiblc2=2.241917513e-14
+  pdiblcb=1.220200939e-03 lpdiblcb=-1.316254488e-07 wpdiblcb=-2.852715292e-09 ppdiblcb=2.853386251e-13
+  drout=0.56
+  pscbe1=7.800989187e+08 lpscbe1=-3.363169700e+03 wpscbe1=-1.329133902e+02 ppscbe1=1.329446514e-2
+  pscbe2=9.388803122e-09 lpscbe2=1.162167058e-14 wpscbe2=4.541851576e-16 ppscbe2=-4.542919819e-20
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=-1.334896019e-10 lalpha0=2.335445187e-14 walpha0=6.960960125e-16 palpha0=-6.962597342e-20
+  alpha1=1.621675242e-10 lalpha1=-6.218214601e-15 walpha1=-1.853382992e-16 palpha1=1.853818908e-20
+  beta0=5.107119932e+00 lbeta0=-3.148048563e-05 wbeta0=3.991726618e-07 pbeta0=-3.992665472e-11
* Gidl Induced Drain Leakage Model Parameters
+  agidl=-1.840057134e-10 lagidl=2.773961416e-14 wagidl=8.636410237e-16 pagidl=-8.638441521e-20
+  bgidl=9.123199415e+08 lbgidl=2.421816062e+04 wbgidl=8.370851749e+02 pbgidl=-8.372820574e-2
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-5.154304340e-01 lkt1=7.375777779e-06 wkt1=2.301750850e-07 pkt1=-2.302292222e-11
+  kt2=-0.037961
+  at=0.0
+  ute=-2.802778133e-01 lute=-2.038698055e-06 wute=-3.910281622e-08 pute=3.911201320e-12
+  ua1=2.318865459e-09 lua1=-1.072906873e-14 wua1=-5.343184250e-16 pua1=5.344440967e-20
+  ub1=-1.045453622e-18 lub1=2.519228602e-23 wub1=1.412905181e-24 pub1=-1.413237496e-28
+  uc1=2.340289505e-10 luc1=-1.142058054e-14 wuc1=-5.687564091e-16 puc1=5.688901806e-20
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.19 pmos
* Model Flag Parameters
+  lmin=8.0e-06 lmax=2.0e-05 wmin=3.0e-06 wmax=5.0e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.153902212e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} wvth0=2.488205755e-7
+  k1=3.571106828e-01 wk1=3.838972541e-7
+  k2=6.511888172e-02 wk2=-1.551120217e-7
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-3.107454742e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} wvoff=3.764537246e-7
+  nfactor={-1.611077765e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} wnfactor=1.228101212e-5
+  eta0=0.08
+  etab=-0.07
+  u0=1.050324010e-02 wu0=-6.890016229e-9
+  ua=-1.635148261e-09 wua=4.031285154e-15
+  ub=2.396934983e-18 wub=-6.555952368e-24
+  uc=-3.536616325e-11 wuc=-2.201258754e-16
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=160312.5
+  a0=1.660854905e+00 wa0=1.372188671e-8
+  ags=6.988813575e-01 wags=-8.789290933e-7
+  a1=0.0
+  a2=0.8
+  b0=0.0
+  b1=0.0
+  keta=-7.819866770e-02 wketa=1.400085608e-7
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=3.473505552e-01 wpclm=-8.562344069e-7
+  pdiblc1=0.39
+  pdiblc2=-1.338660609e-05 wpdiblc2=8.955030236e-10
+  pdiblcb=-5.353341015e-03 wpdiblcb=1.139745776e-8
+  drout=0.56
+  pscbe1=6.121379558e+08 wpscbe1=5.310290705e+2
+  pscbe2=9.969204099e-09 wpscbe2=-1.814606653e-15
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.032861363e-09 walpha0=-2.781113460e-15
+  alpha1=-1.483780043e-10 walpha1=7.404823896e-16
+  beta0=3.534944529e+00 wbeta0=-1.594815144e-6
* Gidl Induced Drain Leakage Model Parameters
+  agidl=1.201345821e-09 wagidl=-3.450506299e-15
+  bgidl=2.121805617e+09 wbgidl=-3.344407676e+3
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-1.470747314e-01 wkt1=-9.196188682e-7
+  kt2=-0.037961
+  at=0.0
+  ute=-3.820929814e-01 wute=1.562275413e-7
+  ua1=1.783042150e-09 wua1=2.134763219e-15
+  ub1=2.126811126e-19 wub1=-5.644982224e-24
+  uc1=-3.363293351e-10 wuc1=2.272353349e-15
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.20 pmos
* Model Flag Parameters
+  lmin=4.0e-06 lmax=8.0e-06 wmin=3.0e-06 wmax=5.0e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.143929921e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-8.001287539e-08 wvth0=1.768724314e-07 pvth0=5.772773731e-13
+  k1=2.598280247e-01 lk1=7.805493535e-07 wk1=5.729334777e-07 pk1=-1.516735921e-12
+  k2=1.131204395e-01 lk2=-3.851414589e-07 wk2=-2.734251945e-07 pk2=9.492881083e-13
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-3.466078850e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=2.877427706e-07 wvoff=4.635599004e-07 pvoff=-6.988981437e-13
+  nfactor={-2.982470790e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.100339936e-05 wnfactor=1.696179421e-05 pnfactor=-3.755634870e-11
+  eta0=0.08
+  etab=-0.07
+  u0=3.622134379e-03 lu0=5.521068938e-08 wu0=2.039365886e-08 pu0=-2.189111127e-13
+  ua=-3.362611847e-09 lua=1.386033863e-14 wua=1.115043877e-14 pua=-5.712067140e-20
+  ub=3.394594119e-18 lub=-8.004738034e-24 wub=-1.082353036e-23 pub=3.424099734e-29
+  uc=4.490116745e-11 luc=-6.440265333e-16 wuc=-5.590472244e-16 puc=2.719342222e-21
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=2.312313388e+05 lvsat=-5.690187217e-01 wvsat=-2.815507220e-02 pvsat=2.259027849e-7
+  a0=1.352419069e+00 la0=2.474741098e-06 wa0=1.043103919e-06 pa0=-8.259267323e-12
+  ags=3.434426014e-01 lags=2.851869968e-06 wags=1.797785483e-07 pags=-8.494561936e-12
+  a1=0.0
+  a2=0.8
+  b0=0.0
+  b1=0.0
+  keta=-6.512733318e-02 lketa=-1.048781139e-07 wketa=8.239588087e-08 pketa=4.622564896e-13
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=6.021009426e-02 lpclm=2.303877232e-06 wpclm=-1.717503472e-06 ppclm=6.910409570e-12
+  pdiblc1=0.39
+  pdiblc2=-2.431161254e-04 lpdiblc2=1.843239393e-09 wpdiblc2=1.796271605e-09 ppdiblc2=-7.227334728e-15
+  pdiblcb=-7.019781344e-03 lpdiblcb=1.337071731e-08 wpdiblcb=1.962648361e-08 ppdiblcb=-6.602575347e-14
+  drout=0.56
+  pscbe1=6.135808014e+08 lpscbe1=-1.157670052e+01 wpscbe1=4.975180255e+02 ppscbe1=2.688765398e-4
+  pscbe2=1.166373232e-08 lpscbe2=-1.359608106e-14 wpscbe2=-7.490527251e-15 ppscbe2=4.554086244e-20
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.971207950e-09 lalpha0=-7.528842612e-15 walpha0=-5.578579868e-15 palpha0=2.244552767e-20
+  alpha1=-3.982164713e-10 lalpha1=2.004583936e-15 walpha1=1.485318816e-15 palpha1=-5.976209961e-21
+  beta0=2.172240540e+00 lbeta0=1.093368271e-05 wbeta0=-8.604491362e-06 pbeta0=5.624227732e-11
* Gidl Induced Drain Leakage Model Parameters
+  agidl=-2.293026917e-07 lagidl=1.849453755e-12 wagidl=6.835872708e-13 pagidl=-5.512461346e-18
+  bgidl=9.745385433e+08 lbgidl=9.205120314e+03 wbgidl=-5.187374917e+02 pbgidl=-2.267182124e-2
+  cgidl=300.0
+  egidl=-4.255642992e-01 legidl=4.216875666e-06 wegidl=1.566850129e-06 pegidl=-1.257165335e-11
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=1.954414237e-01 lkt1=-2.748185221e-06 wkt1=-2.104937094e-06 pkt1=9.510424490e-12
+  kt2=-3.133225080e-02 lkt2=-5.318590178e-8
+  at=-1.896342590e+05 lat=1.521534270e+00 wat=2.733626154e-02 pat=-2.193330412e-7
+  ute=9.866349256e-01 lute=-1.098201574e-05 wute=-2.446543066e-06 pute=2.088338202e-11
+  ua1=3.916344793e-09 lua1=-1.711659642e-14 wua1=4.282078845e-15 pua1=-1.722902987e-20
+  ub1=-1.318203050e-19 lub1=2.764114014e-24 wub1=-1.226730362e-23 pub1=5.313432813e-29
+  uc1=-7.356328499e-10 luc1=3.203819737e-15 wuc1=4.558068135e-15 puc1=-1.833947830e-20
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.21 pmos
* Model Flag Parameters
+  lmin=2.0e-06 lmax=4.0e-06 wmin=3.0e-06 wmax=5.0e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.218135999e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=2.185567614e-07 wvth0=5.601393161e-07 pvth0=-9.648046027e-13
+  k1=2.337095284e-01 lk1=8.856376457e-07 wk1=1.089382744e-06 pk1=-3.594679874e-12
+  k2=8.144511033e-02 lk2=-2.576951385e-07 wk2=-2.815494145e-07 pk2=9.819760698e-13
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-3.453449132e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=2.826611782e-07 wvoff=6.058615845e-07 pvoff=-1.271451816e-12
+  nfactor={-1.651034109e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=5.646337247e-06 wnfactor=1.443116293e-05 pnfactor=-2.737430312e-11
+  eta0=0.08
+  etab=-0.07
+  u0=2.637391328e-02 lu0=-3.633154807e-08 wu0=-6.842453122e-08 pu0=1.384506514e-13
+  ua=2.071881725e-09 lua=-8.005454944e-15 wua=-1.052846122e-14 pua=3.010481628e-20
+  ub=4.022273774e-19 lub=4.035109401e-24 wub=1.380378206e-24 pub=-1.486167284e-29
+  uc=-2.088903783e-10 luc=3.771088269e-16 wuc=4.236329707e-16 puc=-1.234491196e-21
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=1.714936062e+05 lvsat=-3.286627596e-01 wvsat=-7.751152270e-02 pvsat=4.244894506e-7
+  a0=1.504063772e+00 la0=1.864595602e-06 wa0=1.755109275e-06 pa0=-1.112403511e-11
+  ags=3.994891645e-01 lags=2.626365500e-06 wags=2.111438702e-07 pags=-8.620760936e-12
+  a1=0.0
+  a2=0.8
+  b0=0.0
+  b1=0.0
+  keta=-3.610420826e-02 lketa=-2.216532375e-07 wketa=-1.598034031e-08 pketa=8.580751830e-13
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=6.209306932e-01 lpclm=4.780668739e-08 wpclm=9.478412961e-07 ppclm=-3.813658412e-12
+  pdiblc1=0.39
+  pdiblc2=0.000215
+  pdiblcb=-4.125487681e-02 lpdiblcb=1.511163086e-07 wpdiblcb=1.827002066e-07 ppdiblcb=-7.221561393e-13
+  drout=0.56
+  pscbe1=4.205172038e+08 lpscbe1=7.652185455e+02 wpscbe1=1.131341435e+03 ppscbe1=-2.281324624e-3
+  pscbe2=-2.585559726e-09 lpscbe2=4.373623047e-14 wpscbe2=5.792334199e-14 ppscbe2=-2.176531487e-19
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=-2.793179990e-03 lalpha0=1.123841596e-08 walpha0=8.327229593e-09 palpha0=-3.350477481e-14
+  alpha1=3.519925879e-10 lalpha1=-1.013897217e-15 walpha1=-7.512584466e-16 palpha1=3.022703385e-21
+  beta0=-6.473634889e+01 lbeta0=2.801417305e-04 wbeta0=2.095317689e-04 pbeta0=-8.214333287e-10
* Gidl Induced Drain Leakage Model Parameters
+  agidl=4.633682952e-07 lagidl=-9.375218141e-13 wagidl=-1.381118197e-12 pagidl=2.794922397e-18
+  bgidl=5.092119605e+09 lbgidl=-7.362049439e+03 wbgidl=-1.177622993e+04 pbgidl=2.262292474e-2
+  cgidl=300.0
+  egidl=1.151128598e+00 legidl=-2.126979741e-06 wegidl=-3.133700259e-06 pegidl=6.341105147e-12
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-5.574049919e-01 lkt1=2.809073892e-07 wkt1=6.407332863e-07 pkt1=-1.536835198e-12
+  kt2=-3.970993539e-02 lkt2=-1.947812028e-08 wkt2=-1.154954685e-09 pkt2=4.646983276e-15
+  at=3.718000333e+05 lat=-7.374078337e-01 wat=-2.848435442e-01 pat=1.036728651e-6
+  ute=-3.335977105e+00 lute=6.410100220e-06 wute=5.012545996e-06 pute=-9.128412000e-12
+  ua1=-2.370081736e-09 lua1=8.176966447e-15 wua1=-2.848973367e-15 pua1=1.146290132e-20
+  ub1=2.114256973e-18 lub1=-6.273022835e-24 wub1=3.267379227e-24 pub1=-9.369778976e-30
+  uc1=2.798421021e-11 luc1=1.313912233e-16 wuc1=1.929761629e-16 puc1=-7.764434508e-22
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.22 pmos
* Model Flag Parameters
+  lmin=1.0e-06 lmax=2.0e-06 wmin=3.0e-06 wmax=5.0e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.119575034e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=1.911667783e-08 wvth0=9.657632174e-08 pvth0=-2.677561239e-14
+  k1=9.195973498e-01 lk1=-5.022700787e-07 wk1=-1.453676532e-06 pk1=1.551251432e-12
+  k2=-1.285370450e-01 lk2=1.672079526e-07 wk2=4.615143665e-07 pk2=-5.216283524e-13
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=7.186915507e-02 ldsub=9.877425273e-07 wdsub=9.358161955e-07 pdsub=-1.893642788e-12
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.049227550e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-1.485867303e-09 wvoff=-5.052876758e-08 pvoff=5.676718944e-14
+  nfactor={8.443078793e-01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=5.969628277e-07 wnfactor=7.370578731e-07 pnfactor=3.359923365e-13
+  eta0=-6.482533088e-02 leta0=2.930569535e-07 weta0=7.633953140e-09 peta0=-1.544745686e-14
+  etab=-6.381137200e-01 letab=1.149589475e-06 wetab=4.021247288e-06 petab=-8.137074312e-12
+  u0=4.604665615e-03 lu0=7.718959966e-09 wu0=1.122688041e-08 pu0=-2.272557303e-14
+  ua=-3.413120761e-09 lua=3.093557285e-15 wua=1.001561823e-14 pua=-1.146653936e-20
+  ub=3.828436208e-18 lub=-2.897892692e-24 wub=-1.185315737e-23 pub=1.191665108e-29
+  uc=2.528989018e-11 luc=-9.675962994e-17 wuc=-4.412533190e-16 puc=5.156235087e-22
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=-6.532160438e+04 lvsat=1.505375553e-01 wvsat=3.137671611e-01 pvsat=-3.672707916e-7
+  a0=3.787851474e+00 la0=-2.756694489e-06 wa0=-7.773819892e-06 pa0=8.157943634e-12
+  ags=2.843619634e+00 lags=-2.319381388e-06 wags=-8.282395587e-06 pags=8.566086027e-12
+  a1=0.0
+  a2=0.8
+  b0=0.0
+  b1=0.0
+  keta=-2.828745321e-01 lketa=2.776914481e-07 wketa=8.361277157e-07 pketa=-8.661825104e-13
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=7.144552896e-01 lpclm=-1.414422040e-07 wpclm=-2.037722091e-06 ppclm=2.227688814e-12
+  pdiblc1=3.769599201e-01 lpdiblc1=2.638686241e-08 wpdiblc1=9.690198789e-08 ppdiblc1=-1.960831105e-13
+  pdiblc2=-5.056800000e-06 lpdiblc2=4.452893359e-10
+  pdiblcb=9.322424029e-02 lpdiblcb=-1.210048744e-07 wpdiblcb=-3.524586173e-07 ppdiblcb=3.607484440e-13
+  drout=8.530688465e-01 ldrout=-5.930306722e-07 wdrout=-2.186985988e-06 pdrout=4.425409887e-12
+  pscbe1=7.973275178e+08 lpscbe1=2.735338973e+00 wpscbe1=7.967396330e+00 ppscbe1=-8.154789491e-6
+  pscbe2=2.919713530e-08 lpscbe2=-2.057668856e-14 wpscbe2=-1.010373883e-13 ppscbe2=1.040070682e-19
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=5.550299318e-03 lalpha0=-5.644781295e-09 walpha0=-1.654695165e-08 palpha0=1.682862842e-14
+  alpha1=-1.490636000e-10 walpha1=7.425263369e-16
+  beta0=9.108816238e+01 lbeta0=-3.517228460e-05 wbeta0=-2.514104108e-04 pbeta0=1.112923908e-10
* Gidl Induced Drain Leakage Model Parameters
+  agidl=-1.440503678e-11 lagidl=1.423475334e-16 wagidl=3.352736525e-16 pagidl=-4.763293941e-22
+  bgidl=1.263660399e+09 lbgidl=3.849143340e+02 wbgidl=1.777117686e+01 pbgidl=-1.242472382e-3
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-3.438673538e-01 lkt1=-1.511902922e-07 wkt1=-2.984378561e-07 pkt1=3.635963920e-13
+  kt2=-3.813431627e-02 lkt2=-2.266641708e-08 wkt2=-6.759402200e-08 pkt2=1.390877648e-13
+  at=-1.063506058e+05 lat=2.301395475e-01 wat=5.086774417e-01 pat=-5.689769345e-7
+  ute=3.315259227e+00 lute=-7.048809522e-06 wute=-9.883689505e-06 pute=2.101441846e-11
+  ua1=8.040603263e-09 lua1=-1.288926286e-14 wua1=-1.552927350e-14 pua1=3.712174224e-20
+  ub1=-4.887192482e-18 lub1=7.894550165e-24 wub1=1.000868160e-23 pub1=-2.301093915e-29
+  uc1=-4.461870145e-11 luc1=2.783046671e-16 wuc1=6.016478023e-16 puc1=-1.603398687e-21
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=2.75e-6
+  sbref=2.74e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.23 pmos
* Model Flag Parameters
+  lmin=5.0e-07 lmax=1.0e-06 wmin=3.0e-06 wmax=5.0e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.125210011e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=2.488418900e-08 wvth0=4.028651773e-08 pvth0=3.083812781e-14
+  k1=5.055959375e-01 lk1=-7.853135321e-08 wk1=-5.396698085e-07 pk1=6.157472708e-13
+  k2=1.039530254e-02 lk2=2.500791618e-08 wk2=1.288418683e-07 pk2=-1.811313969e-13
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=1.075564090e+00 ldsub=-3.955931233e-08 wdsub=-1.871632391e-06 pdsub=9.798369894e-13
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-1.416533944e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-6.624332326e-08 wvoff=-2.354536005e-07 pvoff=2.460414544e-13
+  nfactor={4.585070823e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-3.231782860e-06 wnfactor=-1.206196041e-05 pnfactor=1.343604353e-11
+  eta0=4.298444042e-01 leta0=-2.132474137e-07 weta0=-1.840075693e-07 peta0=1.807014742e-13
+  etab=9.924805620e-01 letab=-5.193563848e-07 wetab=-8.039580747e-06 petab=4.207424399e-12
+  u0=1.607401453e-02 lu0=-4.020148031e-09 wu0=-1.383427230e-08 pu0=2.925017987e-15
+  ua=6.848944077e-10 lua=-1.100843200e-15 wua=-2.840566974e-15 pua=1.692023315e-21
+  ub=2.107514272e-19 lub=8.048800346e-25 wub=1.715038464e-24 pub=-1.970668725e-30
+  uc=-1.636235744e-10 luc=9.659707935e-17 wuc=2.929718161e-16 puc=-2.358706016e-22
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=-1.304478408e+04 lvsat=9.703118417e-02 wvsat=1.879548220e-01 pvsat=-2.384993463e-7
+  a0=7.739346593e-01 la0=3.281096490e-07 wa0=1.089837019e-06 pa0=-9.141864873e-13
+  ags=2.667888633e-01 lags=3.180564430e-07 wags=-1.003954268e-06 pags=1.116455768e-12
+  a1=0.0
+  a2=1.030543051e+00 la2=-2.359654231e-07 wa2=-1.311582533e-06 pa2=1.342430954e-12
+  b0=0.0
+  b1=0.0
+  keta=-1.288042003e-02 lketa=1.347074567e-09 wketa=9.363987754e-08 pketa=-1.062313584e-13
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=6.419291245e-01 lpclm=-6.721022351e-08 wpclm=-3.281358507e-07 ppclm=4.778931049e-13
+  pdiblc1=1.351757863e+00 lpdiblc1=-9.713383280e-07 wpdiblc1=-4.887435445e-06 ppdiblc1=4.905485939e-12
+  pdiblc2=-1.719686927e-03 lpdiblc2=2.200247563e-09 wpdiblc2=4.574733600e-09 ppdiblc2=-4.682331334e-15
+  pdiblcb=1.349796040e-02 lpdiblcb=-3.940343243e-08 wpdiblcb=-1.917688122e-07 ppdiblcb=1.962792147e-13
+  drout=2.340769612e-01 ldrout=4.051990225e-08 wdrout=2.314556472e-06 pdrout=-1.820088520e-13
+  pscbe1=7.863501317e+08 lpscbe1=1.397091322e+01 wpscbe1=6.799370684e+01 ppscbe1=-6.959291882e-5
+  pscbe2=8.798412926e-09 lpscbe2=3.018117566e-16 wpscbe2=1.615384159e-15 ppscbe2=-1.060097446e-21
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=7.212202280e-05 lalpha0=-3.775726902e-11 walpha0=-2.150150690e-10 palpha0=1.125646889e-16
+  alpha1=-4.098431517e-10 lalpha1=2.669130868e-16 walpha1=1.519981113e-15 palpha1=-7.957405121e-22
+  beta0=1.067416489e+02 lbeta0=-5.119394112e-05 wbeta0=-2.930866800e-04 pbeta0=1.539488859e-10
* Gidl Induced Drain Leakage Model Parameters
+  agidl=2.748904206e-10 lagidl=-1.537521531e-16 wagidl=-4.521130291e-16 pagidl=3.295766223e-22
+  bgidl=2.185674947e+09 lbgidl=-5.587859968e+02 wbgidl=-2.689980934e+03 pbgidl=1.528966058e-3
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.920101620e-01 lkt1=4.368348712e-10 wkt1=1.170410050e-07 pkt1=-6.165453190e-14
+  kt2=-1.084289843e-01 lkt2=4.928158154e-08 wkt2=2.437762368e-07 pkt2=-1.796059226e-13
+  at=1.651193588e+05 lat=-4.771539069e-02 wat=2.499309910e-02 pat=-7.391633617e-8
+  ute=-7.055508399e+00 lute=3.565878559e-06 wute=2.109681986e-05 pute=-1.069475248e-11
+  ua1=-1.250648107e-08 lua1=8.141088891e-15 wua1=4.524161583e-14 pua1=-2.507847841e-20
+  ub1=8.192226211e-18 lub1=-5.492496455e-24 wub1=-2.748667311e-23 pub1=1.536630631e-29
+  uc1=8.301520091e-10 luc1=-6.170406505e-16 wuc1=-2.843773665e-15 puc1=1.923059093e-21
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.75e-6
+  sbref=1.74e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.24 pmos
* Model Flag Parameters
+  lmin=2.5e-07 lmax=5.0e-07 wmin=3.0e-06 wmax=5.0e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.090977311e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=6.962685976e-09 wvth0=1.725395091e-07 pvth0=-3.839895822e-14
+  k1=-2.259010367e-01 lk1=3.044219427e-07 wk1=2.023433284e-06 pk1=-7.260884600e-13
+  k2=2.714927548e-01 lk2=-1.116818220e-07 wk2=-7.479847939e-07 pk2=2.779048973e-13
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=1.082878138e+00 ldsub=-4.338836296e-08 wdsub=1.103143860e-06 pdsub=-5.775178734e-13
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-1.835178484e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-4.432644431e-08 wvoff=3.760921199e-07 pvoff=-7.411496111e-14
+  nfactor={-5.941624088e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=2.279152460e-06 wnfactor=2.836356028e-05 pnfactor=-7.727525062e-12
+  eta0=-4.889602848e-01 leta0=2.677652171e-07 weta0=3.374793261e-07 peta0=-9.230734528e-14
+  etab=1.591956038e-03 letab=-6.063818155e-10 wetab=-5.827656859e-09 petab=1.593980704e-15
+  u0=1.339511380e-02 lu0=-2.617689922e-09 wu0=-2.287471403e-08 pu0=7.657870040e-15
+  ua=-4.734947761e-10 lua=-4.944032948e-16 wua=-1.691183894e-15 pua=1.090298285e-21
+  ub=1.453488264e-18 lub=1.542824458e-25 wub=-2.303209761e-24 pub=1.329645852e-31
+  uc=4.882544602e-11 luc=-1.462423183e-17 wuc=-2.814205802e-16 puc=6.483530573e-23
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=2.456116777e+05 lvsat=-3.838064673e-02 wvsat=-4.680589143e-01 pvsat=1.049369650e-7
+  a0=2.170576841e+00 la0=-4.030604657e-07 wa0=-1.631984284e-06 pa0=5.107414016e-13
+  ags=1.713448526e-01 lags=3.680232914e-07 wags=-6.800044313e-08 pags=6.264652216e-13
+  a1=0.0
+  a2=3.389138989e-01 la2=1.261162704e-07 wa2=2.623165067e-06 pa2=-7.174881090e-13
+  b0=0.0
+  b1=0.0
+  keta=1.422262750e-01 lketa=-7.985438240e-08 wketa=-4.977592543e-07 pketa=2.033779151e-13
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=3.790229365e-01 lpclm=7.042642404e-08 wpclm=1.217641748e-06 ppclm=-3.313523837e-13
+  pdiblc1=-1.314805471e+00 lpdiblc1=4.246609087e-07 wpdiblc1=8.932168704e-06 ppdiblc1=-2.329353226e-12
+  pdiblc2=-4.971783760e-03 lpdiblc2=3.902785297e-09 wpdiblc2=-4.972626522e-09 ppdiblc2=3.159026370e-16
+  pdiblcb=-1.019959208e-01 lpdiblcb=2.105992426e-08 wpdiblcb=3.835376244e-07 ppdiblcb=-1.049052110e-13
+  drout=1.567527797e-01 ldrout=8.100065770e-08 wdrout=4.166098877e-06 pdrout=-1.151328332e-12
+  pscbe1=8.270594435e+08 lpscbe1=-7.341225704e+00 wpscbe1=-1.347904482e+02 ppscbe1=3.656864205e-5
+  pscbe2=3.181440245e-08 lpscbe2=-1.174751908e-14 wpscbe2=-6.699227535e-14 ppscbe2=3.485738446e-20
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=8.936650713e+00 lbeta0=8.931534583e-09 wbeta0=2.871939058e-06 pbeta0=-9.913703680e-13
* Gidl Induced Drain Leakage Model Parameters
+  agidl=-1.096577597e-10 lagidl=4.756651021e-17 wagidl=5.261502869e-16 pagidl=-1.825637889e-22
+  bgidl=7.722061918e+08 lbgidl=1.811931661e+02 wbgidl=1.770579024e+03 pbgidl=-8.062262910e-4
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-5.250421389e-01 lkt1=1.772973540e-08 wkt1=9.215076497e-08 pkt1=-4.862399343e-14
+  kt2=-1.826391978e-03 lkt2=-6.527007592e-09 wkt2=-1.289533345e-07 pkt2=1.552546260e-14
+  at=1.247866472e+05 lat=-2.660040950e-02 wat=-2.966197853e-01 pat=9.445444106e-8
+  ute=-4.377110072e-01 lute=1.013292682e-07 wute=1.180075128e-06 pute=-2.679382821e-13
+  ua1=5.926249790e-09 lua1=-1.508814368e-15 wua1=-1.004401576e-14 pua1=3.864655446e-21
+  ub1=-4.746666054e-18 lub1=1.281272423e-24 wub1=8.412609992e-24 pub1=-3.427686385e-30
+  uc1=-7.780917943e-10 luc1=2.249071454e-16 wuc1=2.264080504e-15 puc1=-7.510047214e-22
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.25e-6
+  sbref=1.24e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.25 pmos
* Model Flag Parameters
+  lmin=1.8e-07 lmax=2.5e-07 wmin=3.0e-06 wmax=5.0e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-9.469552240e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-3.243023519e-08 wvth0=-1.155263751e-07 pvth0=4.039282241e-14
+  k1=1.154733366e+00 lk1=-7.320917920e-08 wk1=-3.908683817e-06 pk1=8.964642093e-13
+  k2=-2.113185875e-01 lk2=2.037673632e-08 wk2=1.487775337e-06 pk2=-3.336202139e-13
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=-1.192934348e+00 ldsub=5.790918683e-07 wdsub=5.509379574e-06 pdsub=-1.782711466e-12
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-1.932227810e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-4.167195115e-08 wvoff=1.219046915e-07 pvoff=-4.589615699e-15
+  nfactor={2.775418974e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.051331588e-07 wnfactor=-3.962968250e-06 pnfactor=1.114427023e-12
+  eta0=0.49
+  etab=-0.000625
+  u0=-9.946903891e-03 lu0=3.766818756e-09 wu0=6.169285085e-08 pu0=-1.547305031e-14
+  ua=-6.595232335e-09 lua=1.180014362e-15 wua=2.025610664e-14 pua=-4.912724620e-21
+  ub=5.273967078e-18 lub=-8.906949194e-25 wub=-1.545719770e-23 pub=3.730843367e-30
+  uc=1.190954363e-10 luc=-3.384447956e-17 wuc=-5.103795080e-16 puc=1.274601517e-22
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=4.966738497e+04 lvsat=1.521403623e-02 wvsat=-3.064917789e-01 pvsat=6.074512207e-8
+  a0=-4.995392958e-01 la0=3.272696999e-07 wa0=3.956718930e-06 pa0=-1.017880702e-12
+  ags=2.292707650e+00 lags=-2.122118610e-07 wags=8.683796291e-06 pags=-1.767326221e-12
+  a1=0.0
+  a2=1.873052142e+00 la2=-2.935012220e-07 wa2=-2.010479305e-06 pa2=5.499062995e-13
+  b0=0.0
+  b1=0.0
+  keta=-6.074305790e-01 lketa=1.251917603e-07 wketa=1.660401490e-06 pketa=-3.869222117e-13
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=9.441754329e-01 lpclm=-8.415408679e-08 wpclm=-1.744064610e-06 ppclm=4.787335394e-13
+  pdiblc1=-1.481867710e-01 lpdiblc1=1.055673618e-07 wpdiblc1=8.364275731e-07 ppdiblc1=-1.150061114e-13
+  pdiblc2=1.386804803e-02 lpdiblc2=-1.250285494e-09 wpdiblc2=-3.359363353e-08 ppdiblc2=8.144320474e-15
+  pdiblcb=-3.129714574e-01 lpdiblcb=7.876595303e-08 wpdiblcb=2.588762559e-06 ppdiblcb=-7.080783353e-13
+  drout=1.693827719e+00 ldrout=-3.394200796e-07 wdrout=-5.875143032e-06 pdrout=1.595152155e-12
+  pscbe1=8.034066367e+08 lpscbe1=-8.717099974e-01 wpscbe1=-1.187249019e+01 ppscbe1=2.948122160e-6
+  pscbe2=-2.778975791e-08 lpscbe2=4.555410864e-15 wpscbe2=1.085471165e-13 ppscbe2=-1.315614999e-20
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=7.743796531e+00 lbeta0=3.352010105e-07 wbeta0=9.116168817e-07 pbeta0=-4.551830465e-13
* Gidl Induced Drain Leakage Model Parameters
+  agidl=2.510417111e-10 lagidl=-5.109200904e-17 wagidl=-5.521594628e-16 pagidl=1.123754939e-22
+  bgidl=2.300401376e+09 lbgidl=-2.367987808e+02 wbgidl=-3.412607655e+03 pbgidl=6.114789294e-4
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-1.005052610e+00 lkt1=1.490221996e-07 wkt1=4.579550579e-07 pkt1=-1.486787836e-13
+  kt2=7.257413394e-02 lkt2=-2.687703944e-08 wkt2=-3.747843083e-07 pkt2=8.276515058e-14
+  at=-5.259389146e+04 lat=2.191671543e-02 wat=5.823224812e-01 pat=-1.459538477e-7
+  ute=2.574251680e+00 lute=-7.225027661e-07 wute=-7.501187748e-06 pute=2.106560740e-12
+  ua1=2.565980705e-09 lua1=-5.897135675e-16 wua1=5.691965406e-15 pua1=-4.394501231e-22
+  ub1=-2.786617816e-18 lub1=7.451600294e-25 wub1=-4.446637674e-24 pub1=8.957503701e-32
+  uc1=1.265632042e-10 luc1=-2.253408975e-17 wuc1=-1.516968850e-15 puc1=2.831878979e-22
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.1e-6
+  sbref=1.1e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.26 pmos
* Model Flag Parameters
+  lmin=1.5e-07 lmax=1.8e-07 wmin=3.0e-06 wmax=5.0e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-2.026e-8
+  vth0={-1.162477536e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=1.238785152e-08 wvth0=2.648464967e-07 pvth0=-4.011299589e-14
+  k1=-1.230503357e+00 lk1=4.466680696e-07 wk1=4.184180238e-06 pk1=-8.132926295e-13
+  k2=6.565337073e-01 lk2=-1.692999855e-07 wk2=-1.407538911e-06 pk2=2.769872298e-13
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=1.021009696e+01 ldsub=-1.887133126e-06 wdsub=-2.364145784e-05 pdsub=4.496721537e-12
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-5.365070073e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=3.054823359e-08 wvoff=-1.656101669e-07 pvoff=5.842979087e-14
+  nfactor={2.447141143e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-4.152309106e-08 wnfactor=7.015636815e-06 pnfactor=-1.213487017e-12
+  eta0=2.205658168e+00 leta0=-3.783369393e-07 weta0=-2.562894499e-09 peta0=5.651694949e-16
+  etab=4.097131148e-01 letab=-9.048776107e-08 wetab=-1.226766076e-06 petab=2.705264550e-13
+  u0=3.906903833e-02 lu0=-6.727534925e-09 wu0=-9.729241162e-08 pu0=1.829391783e-14
+  ua=7.986081489e-09 lua=-1.936890511e-15 wua=-2.777562689e-14 pua=5.268873986e-21
+  ub=-4.994636342e-18 lub=1.299337872e-24 wub=1.963124772e-23 pub=-3.695223740e-30
+  uc=-2.772734064e-10 luc=5.073575250e-17 wuc=8.298684831e-16 puc=-1.574446049e-22
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=4.568163537e+05 lvsat=-7.329962783e-02 wvsat=2.013247298e-02 pvsat=-6.208025547e-9
+  a0=3.432086684e+00 la0=-5.123956642e-07 wa0=-1.066529941e-05 pa0=2.121543337e-12
+  ags=1.25
+  a1=0.0
+  a2=-2.131395663e+00 la2=5.650434880e-07 wa2=6.471641229e-06 pa2=-1.274637317e-12
+  b0=0.0
+  b1=0.0
+  keta=8.486824401e-02 lketa=-1.701672416e-08 wketa=-1.652510436e-06 pketa=3.113215625e-13
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-6.081563001e-02 lpclm=1.304371621e-07 wpclm=4.379502665e-06 ppclm=-8.316469638e-13
+  pdiblc1=1.847189028e+00 lpdiblc1=-3.256348810e-07 wpdiblc1=1.573092037e-06 ppdiblc1=-2.870618050e-13
+  pdiblc2=3.653656943e-02 lpdiblc2=-6.353584024e-09 wpdiblc2=4.125784267e-08 ppdiblc2=-7.681632994e-15
+  pdiblcb=-6.234950264e+00 lpdiblcb=1.391260030e-06 wpdiblcb=3.523170922e-05 ppdiblcb=-7.965646627e-12
+  drout=-6.158963588e+00 ldrout=1.363925743e-06 wdrout=1.442694909e-05 pdrout=-2.748622341e-12
+  pscbe1=7.935569236e+08 lpscbe1=1.227534912e+00 wpscbe1=1.920856321e+01 ppscbe1=-3.659615462e-6
+  pscbe2=-1.002993965e-07 lpscbe2=2.092574925e-14 wpscbe2=3.271815721e-13 ppscbe2=-6.246835170e-20
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=1.702609762e+01 lbeta0=-1.683732728e-06 wbeta0=-6.916784160e-06 pbeta0=1.233114569e-12
* Gidl Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=7.846252603e+08 lbgidl=7.768039600e+01 wbgidl=6.420906811e+02 pbgidl=-2.315863895e-4
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-1.106e-8
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=1.425385136e+00 lkt1=-3.744901267e-07 wkt1=1.752741834e-06 pkt1=-4.466242835e-13
+  kt2=4.803089799e-01 lkt2=-1.190357634e-07 wkt2=-1.495054038e-06 pkt2=3.367203940e-13
+  at=-9.938417231e+04 lat=3.406560864e-02 wat=1.135612473e-01 pat=-5.477412691e-8
+  ute=-6.463882970e+00 lute=1.210236122e-06 wute=2.411463163e-05 pute=-4.689398996e-12
+  ua1=-1.454946324e-09 lua1=2.477225610e-16 wua1=1.512539435e-14 pua1=-2.556417086e-21
+  ub1=8.817910418e-19 lub1=-1.554368342e-27 wub1=-1.022620809e-23 pub1=1.371568096e-30
+  uc1=2.696402911e-11 luc1=-2.452749352e-18 wuc1=-1.600036035e-16 puc1=7.604571328e-24
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.04e-6
+  sbref=1.04e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.27 pmos
* Model Flag Parameters
+  lmin=2.0e-05 lmax=0.0001 wmin=2.0e-06 wmax=3.0e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.152810438e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=1.649326082e-06 wvth0=8.018621018e-08 pvth0=-1.605610183e-12
+  k1=4.301581266e-01 lk1=1.115754053e-06 wk1=-1.767275182e-08 pk1=3.538706995e-13
+  k2=2.415484789e-02 lk2=-2.215556813e-07 wk2=2.982523348e-08 pk2=-5.972061590e-13
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-1.015598312e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-1.660205885e-06 wvoff=-2.898630543e-07 pvoff=5.804078665e-12
+  nfactor={6.547162456e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-8.087206496e-05 wnfactor=-1.209918617e-05 pnfactor=2.422682962e-10
+  eta0=0.08
+  etab=-0.07
+  u0=2.054120039e-02 lu0=-2.472716456e-07 wu0=-2.216823987e-08 pu0=4.438861945e-13
+  ua=1.229185677e-09 lua=-3.027818265e-14 wua=-4.340836081e-15 pua=8.691881809e-20
+  ub=3.417851123e-19 lub=-2.881294268e-24 wub=1.902061984e-24 pub=-3.808597618e-29
+  uc=-6.510615108e-11 luc=-8.829619220e-16 wuc=-1.392954952e-17 puc=2.789186133e-22
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=3.082463265e+05 lvsat=-2.962155933e+00 wvsat=-2.930971483e-01 pvsat=5.868836610e-6
+  a0=1.043381575e+00 la0=1.245615172e-05 wa0=1.227923994e-06 pa0=-2.458736066e-11
+  ags=4.481922779e-02 lags=7.193355894e-06 wags=1.004985829e-06 pags=-2.012335385e-11
+  a1=0.0
+  a2=1.545456024e+00 la2=-1.492665361e-05 wa2=-1.476951148e-06 pa2=2.957376085e-11
+  b0=0.0
+  b1=0.0
+  keta=8.281659213e-02 lketa=-2.283733859e-06 wketa=-2.726779866e-07 pketa=5.459973119e-12
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-1.683133279e-01 lpclm=4.574563226e-06 wpclm=7.382922603e-07 ppclm=-1.478320984e-11
+  pdiblc1=0.39
+  pdiblc2=1.303775326e-02 lpdiblc2=-2.553151722e-07 wpdiblc2=-2.556148355e-08 ppdiblc2=5.118308771e-13
+  pdiblcb=7.619373436e-03 lpdiblcb=-1.832091216e-07 wpdiblcb=-2.193038908e-08 ppdiblcb=4.391235844e-13
+  drout=0.56
+  pscbe1=8.042132361e+08 lpscbe1=-2.794009115e+02 wpscbe1=-2.048047295e+02 ppscbe1=4.100911597e-3
+  pscbe2=9.293615777e-09 lpscbe2=1.339968409e-15 wpscbe2=7.379645233e-16 ppscbe2=-1.477664739e-20
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=-8.278186408e-10 lalpha0=1.857819511e-14 walpha0=2.766079735e-15 palpha0=-5.538665289e-20
+  alpha1=3.470353598e-10 lalpha1=-4.946517467e-15 walpha1=-7.364796011e-16 palpha1=1.474691402e-20
+  beta0=9.149017509e+00 lbeta0=-1.231249751e-04 wbeta0=-1.165082341e-05 pbeta0=2.332904956e-10
* Gidl Induced Drain Leakage Model Parameters
+  agidl=-9.231481124e-10 lagidl=1.936474504e-14 wagidl=3.067225562e-15 pagidl=-6.141665238e-20
+  bgidl=4.599455427e+08 lbgidl=1.081379123e+04 wbgidl=2.185736304e+03 pbgidl=-4.376613459e-2
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-7.107124024e-01 lkt1=5.109449704e-06 wkt1=8.123637495e-07 pkt1=-1.626638179e-11
+  kt2=-0.037961
+  at=0.0
+  ute=-1.693619384e-01 lute=-3.210332148e-06 wute=-3.697732085e-07 pute=7.404161236e-12
+  ua1=2.139640475e-09 lua1=7.197644988e-15
+  ub1=-2.570000687e-19 lub1=-2.850948640e-23 wub1=-9.376893207e-25 pub1=1.877584087e-29
+  uc1=4.325252718e-11 luc1=7.661548855e-15 puc1=-3.308722450e-36
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.28 pmos
* Model Flag Parameters
+  lmin=8.0e-06 lmax=2.0e-05 wmin=2.0e-06 wmax=3.0e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.070441+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+  k1=0.4858803
+  k2=0.013090076
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-0.18447262+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={2.5083089+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+  eta0=0.08
+  etab=-0.07
+  u0=0.0081921406
+  ua=-2.8294519e-10
+  ub=1.9788962e-19
+  uc=-1.0920239e-10
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=160312.5
+  a0=1.6654576
+  ags=0.40406455
+  a1=0.0
+  a2=0.8
+  b0=0.0
+  b1=0.0
+  keta=-0.031235975
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=0.060146165
+  pdiblc1=0.39
+  pdiblc2=0.00028698955
+  pdiblcb=-0.0015303226
+  drout=0.56
+  pscbe1=790259600.0
+  pscbe2=9.3605355e-9
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=3.0
* Gidl Induced Drain Leakage Model Parameters
+  agidl=4.395183e-11
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-0.45554
+  kt2=-0.037961
+  at=0.0
+  ute=-0.32969
+  ua1=2.4991e-9
+  ub1=-1.6808e-18
+  uc1=4.2588e-10
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.29 pmos
* Model Flag Parameters
+  lmin=4.0e-06 lmax=8.0e-06 wmin=2.0e-06 wmax=3.0e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.084602080e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=1.136217118e-7
+  k1=4.520055508e-01 lk1=2.717947275e-7
+  k2=2.140616637e-02 lk2=-6.672431739e-8
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-1.911172420e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=5.331325740e-8
+  nfactor={2.706977945e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.594025058e-6
+  eta0=0.08
+  etab=-0.07
+  u0=1.046272419e-02 lu0=-1.821807282e-8
+  ua=3.775496570e-10 lua=-5.299493615e-15 pua=-3.308722450e-36
+  ub=-2.359133808e-19 lub=3.480627053e-24 pub=1.540743956e-45
+  uc=-1.426185303e-10 luc=2.681150701e-16
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=2.217873591e+05 lvsat=-4.932447618e-1
+  a0=1.702304594e+00 la0=-2.956425918e-7
+  ags=4.037452334e-01 lags=2.562043175e-9
+  a1=0.0
+  a2=0.8
+  b0=0.0
+  b1=0.0
+  keta=-3.748950581e-02 lketa=5.017532955e-8
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-5.158874480e-01 lpclm=4.621817215e-06 wpclm=1.110223025e-22 ppclm=1.332267630e-27
+  pdiblc1=0.39
+  pdiblc2=3.594023986e-04 lpdiblc2=-5.810059386e-10
+  pdiblcb=-4.365230551e-04 lpdiblcb=-8.776122525e-9
+  drout=0.56
+  pscbe1=7.804619264e+08 lpscbe1=7.861182970e+1
+  pscbe2=9.151205032e-09 lpscbe2=1.679567196e-15
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=-7.139407148e-01 lbeta0=2.979887760e-5
* Gidl Induced Drain Leakage Model Parameters
+  agidl=-8.863176868e-12 lagidl=4.237622639e-16
+  bgidl=8.005398301e+08 lbgidl=1.600372662e+3
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-5.106119300e-01 lkt1=4.418707318e-7
+  kt2=-3.133225080e-02 lkt2=-5.318590178e-8
+  at=-1.804649308e+05 lat=1.447963982e+0
+  ute=1.659976052e-01 lute=-3.977159414e-6
+  ua1=5.352670913e-09 lua1=-2.289568329e-14
+  ub1=-4.246608763e-18 lub1=2.058681792e-23 pub1=-1.232595164e-44
+  uc1=7.932676112e-10 luc1=-2.947741846e-15
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.30 pmos
* Model Flag Parameters
+  lmin=2.0e-06 lmax=4.0e-06 wmin=2.0e-06 wmax=3.0e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.030249984e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-1.050650359e-7
+  k1=5.991182345e-01 lk1=-3.201160977e-7
+  k2=-1.299424793e-02 lk2=7.168643753e-08 wk2=-6.938893904e-24 pk2=1.387778781e-29
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-1.421224013e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-1.438184639e-7
+  nfactor={3.189571823e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-3.535751178e-6
+  eta0=0.08
+  etab=-0.07
+  u0=3.422457921e-03 lu0=1.010857931e-8
+  ua=-1.459651534e-09 lua=2.092522121e-15
+  ub=8.652439039e-19 lub=-9.499013051e-25
+  uc=-6.679231726e-11 luc=-3.697321461e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=1.454941258e+05 lvsat=-1.862774118e-1
+  a0=2.092775327e+00 la0=-1.866709395e-6
+  ags=4.703125816e-01 lags=-2.652730136e-7
+  a1=0.0
+  a2=0.8
+  b0=0.0
+  b1=0.0
+  keta=-4.146445057e-02 lketa=6.616859927e-8
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=9.388625344e-01 lpclm=-1.231398434e-6
+  pdiblc1=0.39
+  pdiblc2=0.000215
+  pdiblcb=2.002775912e-02 lpdiblcb=-9.111457113e-08 ppdiblcb=2.775557562e-29
+  drout=0.56
+  pscbe1=800000000.0
+  pscbe2=1.684351014e-08 lpscbe2=-2.927057626e-14 wpscbe2=1.323488980e-29
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=5.546325391e+00 lbeta0=4.610571722e-6
* Gidl Induced Drain Leakage Model Parameters
+  agidl=1.035556976e-10 lagidl=-2.855732580e-17
+  bgidl=1.142050664e+09 lbgidl=2.262969922e+2
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-3.424855594e-01 lkt1=-2.345890828e-7
+  kt2=-4.009733871e-02 lkt2=-1.791939525e-8
+  at=2.762557340e+05 lat=-3.896607476e-1
+  ute=-1.654632365e+00 lute=3.348181683e-6
+  ua1=-3.325705164e-09 lua1=1.202193642e-14 wua1=-1.654361225e-30 pua1=1.654361225e-36
+  ub1=3.210225146e-18 lub1=-9.415902443e-24 wub1=1.540743956e-39 pub1=-6.162975822e-45
+  uc1=9.271368235e-11 luc1=-1.290491024e-16
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.31 pmos
* Model Flag Parameters
+  lmin=1.0e-06 lmax=2.0e-06 wmin=2.0e-06 wmax=3.0e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.087180700e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=1.013540662e-8
+  k1=4.319945642e-01 lk1=1.806199173e-8
+  k2=2.626747013e-02 lk2=-7.760434200e-9
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=3.857674493e-01 ldsub=3.525630509e-7
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.218714828e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=1.755539745e-8
+  nfactor={1.091537207e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=7.096638280e-7
+  eta0=-6.226469463e-02 leta0=2.878754549e-07 peta0=1.110223025e-28
+  etab=7.107223768e-01 letab=-1.579807344e-06 wetab=3.330669074e-22 petab=1.110223025e-28
+  u0=8.370467731e-03 lu0=9.618249656e-11
+  ua=-5.360904043e-11 lua=-7.526329856e-16
+  ub=-1.474362962e-19 lub=1.099277333e-24
+  uc=-1.227185167e-10 luc=7.619456839e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=3.992446544e+04 lvsat=2.734490745e-2
+  a0=1.180300103e+00 la0=-2.029753060e-8
+  ags=6.547809364e-02 lags=5.539176694e-7
+  a1=0.0
+  a2=0.8
+  b0=0.0
+  b1=0.0
+  keta=-2.414474864e-03 lketa=-1.284980757e-8
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=3.094768240e-02 lpclm=6.057854269e-7
+  pdiblc1=4.094634917e-01 lpdiblc1=-3.938476478e-8
+  pdiblc2=-5.056800000e-06 lpdiblc2=4.452893359e-10
+  pdiblcb=-0.025
+  drout=1.194940541e-01 ldrout=8.913725917e-7
+  pscbe1=800000000.0
+  pscbe2=-4.693562463e-09 lpscbe2=1.431012090e-14 ppscbe2=3.308722450e-36
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=6.758248586e+00 lbeta0=2.158220897e-6
* Gidl Induced Drain Leakage Model Parameters
+  agidl=9.805489728e-11 lagidl=-1.742634638e-17
+  bgidl=1.269621336e+09 lbgidl=-3.184481508e+1
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.439715564e-01 lkt1=-2.923013823e-8
+  kt2=-6.080719617e-02 lkt2=2.398741550e-8
+  at=6.427369205e+04 lat=3.928915392e-2
+  ute=0.0
+  ua1=2.831661075e-09 lua1=-4.376173113e-16
+  ub1=-1.530007496e-18 lub1=1.760531127e-25
+  uc1=1.571903929e-10 luc1=-2.595190157e-16 puc1=1.033975766e-37
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=2.75e-6
+  sbref=2.74e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.32 pmos
* Model Flag Parameters
+  lmin=5.0e-07 lmax=1.0e-06 wmin=2.0e-06 wmax=3.0e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.111696813e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=3.522813877e-8
+  k1=3.245759539e-01 lk1=1.280070877e-7
+  k2=5.361238178e-02 lk2=-3.574849817e-8
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=4.477675013e-01 ldsub=2.891047577e-7
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.206309585e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=1.628569604e-8
+  nfactor={5.391600791e-01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.275032866e-6
+  eta0=3.681232431e-01 leta0=-1.526352071e-7
+  etab=-1.704214254e+00 letab=8.919285964e-7
+  u0=1.143362200e-02 lu0=-3.039017162e-09 wu0=-1.387778781e-23
+  ua=-2.679092862e-10 lua=-5.332923980e-16
+  ub=7.860221385e-19 lub=1.438639564e-25
+  uc=-6.535283089e-11 luc=1.747964170e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=5.000039328e+04 lvsat=1.703199379e-2
+  a0=1.139495742e+00 la0=2.146654927e-8
+  ags=-6.996480032e-02 lags=6.925461803e-07 pags=-4.440892099e-28
+  a1=0.0
+  a2=5.906024704e-01 la2=2.143225595e-7
+  b0=0.0
+  b1=0.0
+  keta=1.852895072e-02 lketa=-3.428582252e-8
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=5.318634040e-01 lpclm=9.308816755e-8
+  pdiblc1=-2.876213835e-01 lpdiblc1=6.740955467e-7
+  pdiblc2=-1.851964142e-04 lpdiblc2=6.296658339e-10
+  pdiblcb=-5.082653338e-02 lpdiblcb=2.643397344e-8
+  drout=1.010442376e+00 ldrout=-2.053083449e-8
+  pscbe1=8.091570768e+08 lpscbe1=-9.372451233e+0
+  pscbe2=9.340256864e-09 lpscbe2=-5.377386132e-17
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=8.432376873e+00 lbeta0=4.447171140e-7
* Gidl Induced Drain Leakage Model Parameters
+  agidl=1.232393706e-10 lagidl=-4.320315848e-17
+  bgidl=1.283381922e+09 lbgidl=-4.592904908e+1
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.527514144e-01 lkt1=-2.024377793e-8
+  kt2=-2.665978080e-02 lkt2=-1.096314708e-8
+  at=1.735027264e+05 lat=-7.250894732e-2
+  ute=2.094080000e-02 lute=-2.143332762e-8
+  ua1=2.668791712e-09 lua1=-2.709172611e-16
+  ub1=-1.027554176e-18 lub1=-3.382179098e-25
+  uc1=-1.237272963e-10 luc1=2.800585753e-17
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.75e-6
+  sbref=1.74e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.33 pmos
* Model Flag Parameters
+  lmin=2.5e-07 lmax=5.0e-07 wmin=2.0e-06 wmax=3.0e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.033102850e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-5.917372677e-9
+  k1=4.528137145e-01 lk1=6.087205529e-8
+  k2=2.059823932e-02 lk2=-1.846493431e-8
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=1.452902698e+00 ldsub=-2.371036206e-07 wdsub=-1.776356839e-21
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-5.736628630e-02+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-6.918662517e-8
+  nfactor={3.572288190e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-3.128703623e-7
+  eta0=-3.757605076e-01 leta0=2.368028140e-07 weta0=1.110223025e-22 peta0=-5.551115123e-29
+  etab=-3.627991333e-04 letab=-7.171718105e-11
+  u0=5.722310368e-03 lu0=-4.903129582e-11
+  ua=-1.040764014e-09 lua=-1.286874911e-16
+  ub=6.809288462e-19 lub=1.988823968e-25
+  uc=-4.557069771e-11 luc=7.123299332e-18
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=8.861194262e+04 lvsat=-3.181924523e-3
+  a0=1.623164768e+00 la0=-2.317438593e-7
+  ags=1.485356480e-01 lags=5.781568256e-7
+  a1=0.0
+  a2=1.218795059e+00 la2=-1.145488246e-7
+  b0=0.0
+  b1=0.0
+  keta=-2.473576480e-02 lketa=-1.163587865e-8
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=7.874532133e-01 lpclm=-4.071820942e-8
+  pdiblc1=1.681287708e+00 lpdiblc1=-3.566677408e-7
+  pdiblc2=-6.639738419e-03 lpdiblc2=4.008747664e-09 wpdiblc2=1.734723476e-24 ppdiblc2=1.734723476e-30
+  pdiblcb=2.665306675e-02 lpdiblcb=-1.412814682e-08 wpdiblcb=5.204170428e-24 ppdiblcb=-8.673617380e-31
+  drout=1.554176053e+00 ldrout=-3.051862892e-7
+  pscbe1=7.818470482e+08 lpscbe1=4.924894947e+0
+  pscbe2=9.343364803e-09 lpscbe2=-5.540092987e-17
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=9.899977460e+00 lbeta0=-3.236011454e-7
* Gidl Induced Drain Leakage Model Parameters
+  agidl=6.682740736e-11 lagidl=-1.367036750e-17
+  bgidl=1.366106723e+09 lbgidl=-8.923713710e+1
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.941322571e-01 lkt1=1.419920859e-9
+  kt2=-4.508086002e-02 lkt2=-1.319343681e-9
+  at=2.529227521e+04 lat=5.082188084e-3
+  ute=-4.188160000e-02 lute=1.145545523e-8
+  ua1=2.557212761e-09 lua1=-2.125034486e-16
+  ub1=-1.924847048e-18 lub1=1.315328544e-25
+  uc1=-1.865739702e-11 luc1=-2.700033615e-17
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.25e-6
+  sbref=1.24e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.34 pmos
* Model Flag Parameters
+  lmin=1.8e-07 lmax=2.5e-07 wmin=2.0e-06 wmax=3.0e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-9.857058982e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-1.888138695e-08 wvth0=-7.506586996e-14 pvth0=2.053201698e-20
+  k1=-1.563457235e-01 lk1=2.274893448e-07 wk1=-4.360840187e-13 pk1=1.192777006e-19
+  k2=2.877218865e-01 lk2=-9.152859427e-08 wk2=-5.440924422e-14 pk2=1.488201651e-20
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=6.550619064e-01 ldsub=-1.887820719e-08 wdsub=8.519164929e-14 pdsub=-2.330161930e-20
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-1.523326051e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-4.321143764e-08 wvoff=-4.482349780e-14 pvoff=1.226012336e-20
+  nfactor={1.446131443e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=2.686760312e-07 wnfactor=-5.535431029e-13 pnfactor=1.514051107e-19
+  eta0=0.49
+  etab=-0.000625
+  u0=1.074656242e-02 lu0=-1.423264717e-09 wu0=-8.424656528e-16 pu0=2.304312054e-22
+  ua=1.992187916e-10 lua=-4.678475880e-16 wua=-2.646207226e-22 pua=7.237906130e-29
+  ub=8.920119077e-20 lub=3.607317451e-25 wub=-3.377424088e-31 pub=9.237930208e-38
+  uc=-5.209978104e-11 luc=8.909134205e-18 wuc=-8.100667627e-26 puc=2.215693744e-32
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=-5.313832696e+04 lvsat=3.558960921e-02 wvsat=1.155693620e-08 pvsat=-3.161053290e-15
+  a0=8.276522243e-01 la0=-1.415526839e-08 wa0=1.269099315e-14 pa0=-3.471240628e-21
+  ags=5.205489786e+00 lags=-8.050212702e-07 wags=4.684864692e-13 pags=-1.281404192e-19
+  a1=0.0
+  a2=1.198682166e+00 la2=-1.090475461e-07 wa2=1.022839776e-12 pa2=-2.797671352e-19
+  b0=0.0
+  b1=0.0
+  keta=-5.048659977e-02 lketa=-4.592510270e-09 wketa=-6.750531245e-16 pketa=1.846405806e-22
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=3.591685616e-01 lpclm=7.642620852e-08 wpclm=-4.455349867e-15 ppclm=1.218626977e-21
+  pdiblc1=1.323738849e-01 lpdiblc1=6.699116803e-08 wpdiblc1=-5.467926023e-14 ppdiblc1=1.495587121e-20
+  pdiblc2=2.599826658e-03 lpdiblc2=1.481541824e-09 wpdiblc2=-6.561512167e-16 ppdiblc2=1.794704871e-22
+  pdiblcb=5.553700604e-01 lpdiblcb=-1.587428189e-07 wpdiblcb=3.059338559e-13 ppdiblcb=-8.367902840e-20
+  drout=-2.768556477e-01 ldrout=1.956375016e-07 wdrout=1.098985702e-13 pdrout=-3.005945715e-20
+  pscbe1=7.994242825e+08 lpscbe1=1.171698239e-01 wpscbe1=-8.910694122e-06 ppscbe1=2.437253475e-12
+  pscbe2=8.619907344e-09 lpscbe2=1.424791544e-16 wpscbe2=9.140212890e-22 ppscbe2=-2.500030979e-28
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=8.049577549e+00 lbeta0=1.825202381e-07 wbeta0=4.927884731e-13 pbeta0=-1.347874985e-19
* Gidl Induced Drain Leakage Model Parameters
+  agidl=6.583253563e-11 lagidl=-1.339825019e-17 wagidl=-5.338316465e-22 pagidl=1.460136320e-28
+  bgidl=1.155719483e+09 lbgidl=-3.169201929e+01 wbgidl=4.225829544e-04 pbgidl=-1.155848913e-10
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.00074326333
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.5407449e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-8.514419438e-01 lkt1=9.915126636e-08 wkt1=-1.212394487e-13 pkt1=3.316141406e-20
+  kt2=-5.313874957e-02 lkt2=8.846502693e-10 wkt2=-8.687927044e-15 pkt2=2.376321862e-21
+  at=1.427329404e+05 lat=-2.704018266e-02 wat=6.656019215e-08 pat=-1.820554378e-14
+  ute=5.814857624e-02 lute=-1.590479857e-08 wute=-1.433811908e-14 pute=3.921762332e-21
+  ua1=4.475221582e-09 lua1=-7.371172213e-16 wua1=-9.599248698e-22 pua1=2.625586491e-28
+  ub1=-4.278141744e-18 lub1=7.752060197e-25 wub1=8.505663633e-31 pub1=-2.326469116e-37
+  uc1=-3.822695268e-10 luc1=7.245485357e-17 wuc1=-7.628095000e-23 puc1=2.086436547e-29
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.1e-6
+  sbref=1.1e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.35 pmos
* Model Flag Parameters
+  lmin=1.5e-07 lmax=1.8e-07 wmin=2.0e-06 wmax=3.0e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-2.026e-8
+  vth0={-1.073640688e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-1.067167064e-09 wvth0=-3.110260636e-13 pvth0=7.428099735e-20
+  k1=1.729847659e-01 lk1=1.738675416e-07 wk1=3.937183379e-13 pk1=-5.374706369e-20
+  k2=1.844069818e-01 lk2=-7.639096347e-08 wk2=-7.240327706e-13 pk2=1.637904892e-19
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=2.280106903e+00 ldsub=-3.788100242e-07 wdsub=-5.130828171e-13 pdsub=1.066834843e-19
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-5.920571879e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=5.014718140e-08 wvoff=3.118175407e-14 pvoff=-3.476468446e-21
+  nfactor={4.800376943e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-4.485597115e-07 wnfactor=8.148020072e-13 pnfactor=-1.376955083e-19
+  eta0=2.204798408e+00 leta0=-3.781473450e-07 weta0=2.836796433e-13 peta0=-6.255703422e-20
+  etab=-1.777710849e-03 letab=2.541957964e-10 wetab=9.724808840e-16 petab=-2.144514843e-22
+  u0=6.434507574e-03 lu0=-5.912555053e-10 wu0=1.150462309e-15 pu0=-1.898013795e-22
+  ua=-1.330622280e-09 lua=-1.695662852e-16 wua=1.191177007e-21 pua=-2.426076433e-28
+  ub=1.590219695e-18 lub=5.985902195e-26 wub=7.908878833e-31 pub=-1.487898163e-37
+  uc=1.087131029e-12 luc=-2.075464785e-18 wuc=6.964443600e-24 puc=-1.529654985e-30
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=4.635692546e+05 lvsat=-7.538195110e-02 wvsat=2.385521978e-07 pvsat=-5.348209082e-14
+  a0=-1.453461285e-01 la0=1.992279406e-07 wa0=8.602212773e-13 pa0=-1.906585707e-19
+  ags=1.250000397e+00 lags=-7.569264771e-14 wags=-1.184444535e-12 pags=2.256603722e-19
+  a1=0.0
+  a2=3.937021919e-02 la2=1.374951966e-07 wa2=-2.315453383e-12 pa2=4.330243577e-19
+  b0=0.0
+  b1=0.0
+  keta=-4.694290232e-01 lketa=8.740906114e-08 wketa=4.866082697e-13 pketa=-1.072556547e-19
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=1.408188788e+00 lpclm=-1.485198601e-07 wpclm=9.272768580e-13 ppclm=-2.041451674e-19
+  pdiblc1=2.374847504e+00 lpdiblc1=-4.219233505e-07 wpdiblc1=-1.401834279e-12 ppdiblc1=3.132797581e-19
+  pdiblc2=5.037555360e-02 lpdiblc2=-8.930208479e-09 wpdiblc2=6.666580060e-14 ppdiblc2=-1.465137520e-20
+  pdiblcb=5.582731366e+00 lpdiblcb=-1.280636302e-06 wpdiblcb=-1.412657732e-11 ppdiblcb=3.091988638e-18
+  drout=-1.319771726e+00 ldrout=4.419629311e-07 wdrout=1.889519506e-12 pdrout=-4.250123284e-19
+  pscbe1=7.999999924e+08 lpscbe1=1.439687252e-06 wpscbe1=2.252834320e-05 ppscbe1=-4.292099953e-12
+  pscbe2=9.446233704e-09 lpscbe2=-2.784106864e-17 wpscbe2=-2.237618583e-21 ppscbe2=4.241138171e-28
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=1.470601929e+01 lbeta0=-1.270112403e-06 wbeta0=3.946046263e-13 pbeta0=-1.243947878e-19
* Gidl Induced Drain Leakage Model Parameters
+  agidl=-4.632401722e-15 lagidl=1.007955918e-21 wagidl=1.381044955e-20 pagidl=-3.004990757e-27
+  bgidl=1.000000358e+09 lbgidl=-6.827608728e-05 wbgidl=-1.068389603e-03 pbgidl=2.035495872e-10
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-1.106e-8
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.00074326333
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.5407449e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=2.013303222e+00 lkt1=-5.243002449e-07 wkt1=-1.894948491e-12 pkt1=4.270697014e-19
+  kt2=-2.117299069e-02 lkt2=-6.090544155e-09 wkt2=1.193077246e-13 pkt2=-2.565078544e-20
+  at=-6.129262404e+04 lat=1.569287175e-02 wat=-1.895824913e-08 pat=-8.677238802e-16
+  ute=1.624822846e+00 lute=-3.627163344e-07 wute=-5.347319205e-13 pute=1.190065875e-19
+  ua1=3.618522564e-09 lua1=-6.097692625e-16 wua1=3.606683984e-21 pua1=-7.225384435e-28
+  ub1=-2.548357211e-18 lub1=4.585067958e-25 wub1=-3.146698016e-30 pub1=6.293968617e-37
+  uc1=-2.670561116e-11 luc1=9.804371184e-20 wuc1=1.922656008e-22 puc1=-3.661272209e-29
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.04e-6
+  sbref=1.04e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.36 pmos
* Model Flag Parameters
+  lmin=2.0e-05 lmax=0.0001 wmin=1.68e-06 wmax=2.0e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.112338352e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=8.389324645e-7
+  k1=4.212382248e-01 lk1=1.294361886e-6
+  k2=3.920842634e-02 lk2=-5.229813104e-7
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.478613255e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=1.269265013e-6
+  nfactor={4.403855138e-01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=4.140710528e-05 pnfactor=2.842170943e-26
+  eta0=0.08
+  etab=-0.07
+  u0=9.352307657e-03 lu0=-2.323062827e-8
+  ua=-9.617482694e-10 lua=1.359202704e-14
+  ub=1.301805738e-18 lub=-2.210428646e-23
+  uc=-7.213676046e-11 luc=-7.421843743e-16
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=160312.5
+  a0=1.663147057e+00 la0=4.626521022e-8
+  ags=5.520619633e-01 lags=-2.963429165e-6
+  a1=0.0
+  a2=0.8
+  b0=0.0
+  b1=0.0
+  keta=-5.481114733e-02 lketa=4.720579346e-7
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=2.043221610e-01 lpclm=-2.886910939e-6
+  pdiblc1=0.39
+  pdiblc2=1.362013555e-04 lpdiblc2=3.019310429e-9
+  pdiblcb=-3.449469752e-03 lpdiblcb=3.842808139e-8
+  drout=0.56
+  pscbe1=7.008429116e+08 lpscbe1=1.790436848e+3
+  pscbe2=9.666085849e-09 lpscbe2=-6.118193515e-15
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=5.682944295e-10 lalpha0=-9.376902874e-15
+  alpha1=-2.468523241e-11 lalpha1=2.496637245e-15 walpha1=-1.252080029e-32 palpha1=4.523643975e-37
+  beta0=3.268541021e+00 lbeta0=-5.377136505e-6
* Gidl Induced Drain Leakage Model Parameters
+  agidl=6.249611638e-10 lagidl=-1.163385201e-14
+  bgidl=1.563144045e+09 lbgidl=-1.127612605e+4
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-3.006910881e-01 lkt1=-3.100620284e-6
+  kt2=-0.037961
+  at=0.0
+  ute=-3.559961858e-01 lute=5.267424367e-7
+  ua1=2.139640475e-09 lua1=7.197644988e-15
+  ub1=-7.302764894e-19 lub1=-1.903282652e-23 wub1=1.540743956e-39
+  uc1=4.325252718e-11 luc1=7.661548855e-15
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.37 pmos
* Model Flag Parameters
+  lmin=8.0e-06 lmax=2.0e-05 wmin=1.68e-06 wmax=2.0e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.070441+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+  k1=0.4858803
+  k2=0.013090076
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-0.18447262+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={2.5083089+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+  eta0=0.08
+  etab=-0.07
+  u0=0.0081921406
+  ua=-2.8294519e-10
+  ub=1.9788962e-19
+  uc=-1.0920239e-10
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=160312.5
+  a0=1.6654576
+  ags=0.40406455
+  a1=0.0
+  a2=0.8
+  b0=0.0
+  b1=0.0
+  keta=-0.031235975
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=0.060146165
+  pdiblc1=0.39
+  pdiblc2=0.00028698955
+  pdiblcb=-0.0015303226
+  drout=0.56
+  pscbe1=790259600.0
+  pscbe2=9.3605355e-9
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=3.0
* Gidl Induced Drain Leakage Model Parameters
+  agidl=4.395183e-11
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-0.45554
+  kt2=-0.037961
+  at=0.0
+  ute=-0.32969
+  ua1=2.4991e-9
+  ub1=-1.6808e-18
+  uc1=4.2588e-10
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.38 pmos
* Model Flag Parameters
+  lmin=4.0e-06 lmax=8.0e-06 wmin=1.68e-06 wmax=2.0e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.084602080e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=1.136217118e-7
+  k1=4.520055508e-01 lk1=2.717947275e-7
+  k2=2.140616637e-02 lk2=-6.672431739e-8
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-1.911172420e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=5.331325740e-8
+  nfactor={2.706977945e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.594025058e-6
+  eta0=0.08
+  etab=-0.07
+  u0=1.046272419e-02 lu0=-1.821807282e-8
+  ua=3.775496570e-10 lua=-5.299493615e-15 pua=-3.308722450e-36
+  ub=-2.359133808e-19 lub=3.480627053e-24
+  uc=-1.426185303e-10 luc=2.681150701e-16
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=2.217873591e+05 lvsat=-4.932447618e-1
+  a0=1.702304594e+00 la0=-2.956425918e-7
+  ags=4.037452334e-01 lags=2.562043175e-9
+  a1=0.0
+  a2=0.8
+  b0=0.0
+  b1=0.0
+  keta=-3.748950581e-02 lketa=5.017532955e-8
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-5.158874480e-01 lpclm=4.621817215e-06 ppclm=-1.776356839e-27
+  pdiblc1=0.39
+  pdiblc2=3.594023986e-04 lpdiblc2=-5.810059386e-10
+  pdiblcb=-4.365230551e-04 lpdiblcb=-8.776122525e-9
+  drout=0.56
+  pscbe1=7.804619264e+08 lpscbe1=7.861182970e+1
+  pscbe2=9.151205032e-09 lpscbe2=1.679567196e-15
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=-7.139407148e-01 lbeta0=2.979887760e-5
* Gidl Induced Drain Leakage Model Parameters
+  agidl=-8.863176868e-12 lagidl=4.237622639e-16
+  bgidl=8.005398301e+08 lbgidl=1.600372662e+3
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-5.106119300e-01 lkt1=4.418707318e-7
+  kt2=-3.133225080e-02 lkt2=-5.318590178e-8
+  at=-1.804649308e+05 lat=1.447963982e+0
+  ute=1.659976052e-01 lute=-3.977159414e-06 pute=3.552713679e-27
+  ua1=5.352670913e-09 lua1=-2.289568329e-14
+  ub1=-4.246608763e-18 lub1=2.058681792e-23 wub1=6.162975822e-39 pub1=-2.465190329e-44
+  uc1=7.932676112e-10 luc1=-2.947741846e-15 puc1=-6.617444900e-36
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.39 pmos
* Model Flag Parameters
+  lmin=2.0e-06 lmax=4.0e-06 wmin=1.68e-06 wmax=2.0e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.030249984e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-1.050650359e-7
+  k1=5.991182345e-01 lk1=-3.201160977e-7
+  k2=-1.299424793e-02 lk2=7.168643753e-8
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-1.421224013e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-1.438184639e-7
+  nfactor={3.189571823e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-3.535751178e-6
+  eta0=0.08
+  etab=-0.07
+  u0=3.422457921e-03 lu0=1.010857931e-8
+  ua=-1.459651534e-09 lua=2.092522121e-15 wua=-3.308722450e-30
+  ub=8.652439039e-19 lub=-9.499013051e-25 wub=1.540743956e-39
+  uc=-6.679231726e-11 luc=-3.697321461e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=1.454941258e+05 lvsat=-1.862774118e-1
+  a0=2.092775327e+00 la0=-1.866709395e-6
+  ags=4.703125816e-01 lags=-2.652730136e-7
+  a1=0.0
+  a2=0.8
+  b0=0.0
+  b1=0.0
+  keta=-4.146445057e-02 lketa=6.616859927e-8
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=9.388625344e-01 lpclm=-1.231398434e-06 wpclm=1.776356839e-21
+  pdiblc1=0.39
+  pdiblc2=0.000215
+  pdiblcb=2.002775912e-02 lpdiblcb=-9.111457113e-08 wpdiblcb=6.938893904e-24 ppdiblcb=2.775557562e-29
+  drout=0.56
+  pscbe1=800000000.0
+  pscbe2=1.684351014e-08 lpscbe2=-2.927057626e-14 ppscbe2=5.293955920e-35
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=5.546325391e+00 lbeta0=4.610571722e-6
* Gidl Induced Drain Leakage Model Parameters
+  agidl=1.035556976e-10 lagidl=-2.855732580e-17
+  bgidl=1.142050664e+09 lbgidl=2.262969922e+2
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-3.424855594e-01 lkt1=-2.345890828e-7
+  kt2=-4.009733871e-02 lkt2=-1.791939525e-8
+  at=2.762557340e+05 lat=-3.896607476e-1
+  ute=-1.654632365e+00 lute=3.348181683e-6
+  ua1=-3.325705164e-09 lua1=1.202193642e-14 wua1=3.308722450e-30 pua1=-1.158052858e-35
+  ub1=3.210225146e-18 lub1=-9.415902443e-24 wub1=3.081487911e-39
+  uc1=9.271368235e-11 luc1=-1.290491024e-16
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.40 pmos
* Model Flag Parameters
+  lmin=1.0e-06 lmax=2.0e-06 wmin=1.68e-06 wmax=2.0e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.087180700e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=1.013540662e-8
+  k1=4.319945642e-01 lk1=1.806199173e-8
+  k2=2.626747013e-02 lk2=-7.760434200e-09 wk2=-5.551115123e-23
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=3.857674493e-01 ldsub=3.525630509e-7
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.218714828e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=1.755539745e-8
+  nfactor={1.091537207e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=7.096638280e-7
+  eta0=-6.226469463e-02 leta0=2.878754549e-07 peta0=2.220446049e-28
+  etab=7.107223768e-01 letab=-1.579807344e-06 wetab=4.440892099e-22 petab=1.332267630e-27
+  u0=8.370467731e-03 lu0=9.618249656e-11
+  ua=-5.360904043e-11 lua=-7.526329856e-16
+  ub=-1.474362962e-19 lub=1.099277333e-24
+  uc=-1.227185167e-10 luc=7.619456839e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=3.992446544e+04 lvsat=2.734490745e-2
+  a0=1.180300103e+00 la0=-2.029753060e-8
+  ags=6.547809364e-02 lags=5.539176694e-7
+  a1=0.0
+  a2=0.8
+  b0=0.0
+  b1=0.0
+  keta=-2.414474864e-03 lketa=-1.284980757e-8
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=3.094768240e-02 lpclm=6.057854269e-7
+  pdiblc1=4.094634917e-01 lpdiblc1=-3.938476478e-8
+  pdiblc2=-5.056800000e-06 lpdiblc2=4.452893359e-10
+  pdiblcb=-0.025
+  drout=1.194940541e-01 ldrout=8.913725917e-7
+  pscbe1=800000000.0
+  pscbe2=-4.693562463e-09 lpscbe2=1.431012090e-14 ppscbe2=-1.323488980e-35
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=6.758248586e+00 lbeta0=2.158220897e-6
* Gidl Induced Drain Leakage Model Parameters
+  agidl=9.805489728e-11 lagidl=-1.742634638e-17
+  bgidl=1.269621336e+09 lbgidl=-3.184481508e+1
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.439715564e-01 lkt1=-2.923013823e-8
+  kt2=-6.080719617e-02 lkt2=2.398741550e-8
+  at=6.427369205e+04 lat=3.928915392e-2
+  ute=0.0
+  ua1=2.831661075e-09 lua1=-4.376173113e-16
+  ub1=-1.530007496e-18 lub1=1.760531127e-25
+  uc1=1.571903929e-10 luc1=-2.595190157e-16 wuc1=1.033975766e-31 puc1=1.033975766e-37
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=2.75e-6
+  sbref=2.74e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.41 pmos
* Model Flag Parameters
+  lmin=5.0e-07 lmax=1.0e-06 wmin=1.68e-06 wmax=2.0e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.111696813e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=3.522813877e-8
+  k1=3.245759539e-01 lk1=1.280070877e-7
+  k2=5.361238178e-02 lk2=-3.574849817e-08 wk2=5.551115123e-23
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=4.477675013e-01 ldsub=2.891047577e-7
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.206309585e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=1.628569604e-8
+  nfactor={5.391600791e-01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.275032866e-6
+  eta0=3.681232431e-01 leta0=-1.526352071e-7
+  etab=-1.704214254e+00 letab=8.919285964e-7
+  u0=1.143362200e-02 lu0=-3.039017162e-9
+  ua=-2.679092862e-10 lua=-5.332923980e-16
+  ub=7.860221385e-19 lub=1.438639564e-25
+  uc=-6.535283089e-11 luc=1.747964170e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=5.000039328e+04 lvsat=1.703199379e-2
+  a0=1.139495742e+00 la0=2.146654927e-8
+  ags=-6.996480032e-02 lags=6.925461803e-7
+  a1=0.0
+  a2=5.906024704e-01 la2=2.143225595e-7
+  b0=0.0
+  b1=0.0
+  keta=1.852895072e-02 lketa=-3.428582252e-8
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=5.318634040e-01 lpclm=9.308816755e-8
+  pdiblc1=-2.876213835e-01 lpdiblc1=6.740955467e-7
+  pdiblc2=-1.851964142e-04 lpdiblc2=6.296658339e-10
+  pdiblcb=-5.082653338e-02 lpdiblcb=2.643397344e-8
+  drout=1.010442376e+00 ldrout=-2.053083449e-8
+  pscbe1=8.091570768e+08 lpscbe1=-9.372451233e+0
+  pscbe2=9.340256864e-09 lpscbe2=-5.377386132e-17
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=8.432376873e+00 lbeta0=4.447171140e-7
* Gidl Induced Drain Leakage Model Parameters
+  agidl=1.232393706e-10 lagidl=-4.320315848e-17
+  bgidl=1.283381922e+09 lbgidl=-4.592904908e+1
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.527514144e-01 lkt1=-2.024377793e-8
+  kt2=-2.665978080e-02 lkt2=-1.096314708e-8
+  at=1.735027264e+05 lat=-7.250894732e-2
+  ute=2.094080000e-02 lute=-2.143332762e-8
+  ua1=2.668791712e-09 lua1=-2.709172611e-16
+  ub1=-1.027554176e-18 lub1=-3.382179098e-25
+  uc1=-1.237272963e-10 luc1=2.800585753e-17
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.75e-6
+  sbref=1.74e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.42 pmos
* Model Flag Parameters
+  lmin=2.5e-07 lmax=5.0e-07 wmin=1.68e-06 wmax=2.0e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.167960429e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=6.468326705e-08 wvth0=2.671895451e-07 pvth0=-1.398790707e-13
+  k1=2.077624821e+00 lk1=-7.897490553e-07 wk1=-3.219192751e-06 pk1=1.685311789e-12
+  k2=-6.331318294e-01 lk2=3.237758313e-07 wk2=1.295217081e-06 pk2=-6.780720461e-13
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=1.318067672e+00 ldsub=-1.665147878e-07 wdsub=2.671448616e-07 pdsub=-1.398556779e-13
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-3.659978631e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=9.238817790e-08 wvoff=6.114831014e-07 pvoff=-3.201236332e-13
+  nfactor={5.491269532e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.317495475e-06 wnfactor=-3.802024002e-06 pnfactor=1.990435606e-12
+  eta0=-3.757605076e-01 leta0=2.368028140e-7
+  etab=-3.627991333e-04 letab=-7.171718105e-11
+  u0=-4.443157036e-03 lu0=5.272794200e-09 wu0=2.014055593e-08 pu0=-1.054398384e-14
+  ua=-4.382299405e-09 lua=1.620673117e-15 wua=6.620490508e-15 pua=-3.465959191e-21
+  ub=3.257404976e-18 lub=-1.149954387e-24 wub=-5.104700015e-24 pub=2.672412552e-30
+  uc=1.806154146e-11 luc=-2.618945052e-17 wuc=-1.260727738e-16 puc=6.600161852e-23
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=3.428057138e+05 lvsat=-1.362574476e-01 wvsat=-5.036270013e-01 pvsat=2.636588077e-7
+  a0=1.522062740e+00 la0=-1.788149257e-07 wa0=2.003106169e-07 pa0=-1.048666141e-13
+  ags=-5.601216109e+00 lags=3.588266866e-06 wags=1.139182216e-05 pags=-5.963846739e-12
+  a1=0.0
+  a2=4.399372766e-01 la2=2.931988017e-07 wa2=1.543129117e-06 pa2=-8.078589551e-13
+  b0=0.0
+  b1=0.0
+  keta=-5.753712337e-02 lketa=5.536288585e-09 wketa=6.498841329e-08 pketa=-3.402273413e-14
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=1.333316672e+00 lpclm=-3.264886474e-07 wpclm=-1.081503987e-06 ppclm=5.661889671e-13
+  pdiblc1=2.159762765e+00 lpdiblc1=-6.071590029e-07 wpdiblc1=-9.479892342e-07 ppdiblc1=4.962913239e-13
+  pdiblc2=3.941966512e-03 lpdiblc2=-1.530986501e-09 wpdiblc2=-2.096523569e-08 ppdiblc2=1.097572019e-14
+  pdiblcb=-1.107145511e+00 lpdiblcb=5.794380848e-07 wpdiblcb=2.246363377e-06 ppdiblcb=-1.176016155e-12
+  drout=2.951489307e+00 ldrout=-1.036707724e-06 wdrout=-2.768457626e-06 pdrout=1.449342936e-12
+  pscbe1=7.826839260e+08 lpscbe1=4.486772688e+00 wpscbe1=-1.658082528e+00 ppscbe1=8.680393651e-7
+  pscbe2=1.036100124e-08 lpscbe2=-5.881539572e-16 wpscbe2=-2.016214578e-15 ppscbe2=1.055528656e-21
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=1.120360213e+01 lbeta0=-1.006074730e-06 wbeta0=-2.582835048e-06 pbeta0=1.352165804e-12
* Gidl Induced Drain Leakage Model Parameters
+  agidl=-2.886718541e-11 lagidl=3.642766571e-17 wagidl=1.895970172e-16 pagidl=-9.925783045e-23
+  bgidl=1.139750512e+09 lbgidl=2.926486643e+01 wbgidl=4.484732227e+02 pbgidl=-2.347847015e-4
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.00074326333
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.5407449e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=2.140418490e-01 lkt1=-3.693233872e-07 wkt1=-1.403085528e-06 pkt1=7.345433354e-13
+  kt2=-3.876236123e-02 lkt2=-4.627204171e-09 wkt2=-1.251866475e-08 pkt2=6.553771370e-15
+  at=-1.678384952e+05 lat=1.061900090e-01 wat=3.826445877e-01 pat=-2.003220946e-7
+  ute=-1.554793746e-01 lute=7.092616220e-08 wute=2.250680901e-07 pute=-1.178276465e-13
+  ua1=-2.707542461e-09 lua1=2.543701205e-15 wua1=1.043091211e-14 pua1=-5.460791107e-21
+  ub1=3.611952172e-18 lub1=-2.767092273e-24 wub1=-1.096990526e-23 pub1=5.742964804e-30
+  uc1=4.988412880e-10 luc1=-2.979212477e-16 wuc1=-1.025305655e-15 puc1=5.367680163e-22
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.1e-6
+  sbref=1.1e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.43 pmos
* Model Flag Parameters
+  lmin=1.8e-07 lmax=2.5e-07 wmin=1.68e-06 wmax=2.0e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-5.040717256e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-1.169035711e-07 wvth0=-9.542483755e-07 pvth0=1.942086294e-13
+  k1=-5.959242754e+00 lk1=1.408494964e-06 wk1=1.149711697e-05 pk1=-2.339893245e-12
+  k2=2.622472104e+00 lk2=-5.666969567e-07 wk2=-4.625775288e-06 pk2=9.414377867e-13
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=1.136615614e+00 ldsub=-1.168840207e-07 wdsub=-9.540887914e-07 pdsub=1.941761508e-13
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={9.499230035e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-2.675424975e-07 wvoff=-2.183868219e-06 pvoff=4.444608600e-13
+  nfactor={-5.407373631e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.663501403e-06 wnfactor=1.357865715e-05 pnfactor=-2.763528303e-12
+  eta0=0.49
+  etab=-0.000625
+  u0=4.705180272e-02 lu0=-8.812107194e-09 wu0=-7.193055691e-08 pu0=1.463930694e-14
+  ua=1.213327363e-08 lua=-2.896666419e-15 wua=-2.364460896e-14 pua=4.812150815e-21
+  ub=-9.112499444e-18 lub=2.233461870e-24 wub=1.823107148e-23 pub=-3.710387668e-30
+  uc=-2.793577781e-10 luc=5.516068177e-17 wuc=4.502599063e-16 puc=-9.163689613e-23
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=-9.609732180e+05 lvsat=2.203521658e-01 wvsat=1.798667862e+00 pvsat=-3.660648832e-7
+  a0=1.188730902e+00 la0=-8.764200123e-08 wa0=-7.153950603e-07 pa0=1.455972027e-13
+  ags=2.574031773e+01 lags=-4.984269469e-06 wags=-4.068507916e-05 pags=8.280227310e-12
+  a1=0.0
+  a2=3.980317620e+00 la2=-6.751660299e-07 wa2=-5.511175416e-06 pa2=1.121634421e-12
+  b0=0.0
+  b1=0.0
+  keta=6.666110905e-02 lketa=-2.843441195e-08 wketa=-2.321014760e-07 pketa=4.723729240e-14
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-1.590343793e+00 lpclm=4.731909632e-07 wpclm=3.862514238e-06 ppclm=-7.860988978e-13
+  pdiblc1=-1.576465634e+00 lpdiblc1=4.147741888e-07 wpdiblc1=3.385675836e-06 ppdiblc1=-6.890527462e-13
+  pdiblc2=-3.519197700e-02 lpdiblc2=9.172929728e-09 wpdiblc2=7.487584176e-08 ppdiblc2=-1.523873131e-14
+  pdiblcb=4.604650851e+00 lpdiblcb=-9.828524563e-07 wpdiblcb=-8.022726345e-06 ppdiblcb=1.632785266e-12
+  drout=-5.267260071e+00 ldrout=1.211284606e-06 wdrout=9.887348663e-06 pdrout=-2.012273200e-12
+  pscbe1=7.964354287e+08 lpscbe1=7.254616517e-01 wpscbe1=5.921723315e+00 ppscbe1=-1.205189129e-6
+  pscbe2=4.985491960e-09 lpscbe2=8.821553410e-16 wpscbe2=7.200766350e-15 ppscbe2=-1.465499968e-21
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=3.393775422e+00 lbeta0=1.130069070e-06 wbeta0=9.224410886e-06 pbeta0=-1.877352104e-12
* Gidl Induced Drain Leakage Model Parameters
+  agidl=4.075986690e-10 lagidl=-8.295447478e-17 wagidl=-6.771322043e-16 pagidl=1.378099462e-22
+  bgidl=1.964134735e+09 lbgidl=-1.962207064e+02 wbgidl=-1.601690081e+03 pbgidl=3.259759653e-4
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.00074326333
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.5407449e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-3.380635241e+00 lkt1=6.138926905e-07 wkt1=5.011019741e-06 pkt1=-1.019842738e-12
+  kt2=-7.570482109e-02 lkt2=5.477297452e-09 wkt2=4.470951696e-08 pkt2=-9.099280893e-15
+  at=8.324857254e+05 lat=-1.674186718e-01 wat=-1.366587813e+00 pat=2.781279518e-7
+  ute=4.638549069e-01 lute=-9.847415049e-08 wute=-8.038146075e-07 pute=1.635923489e-13
+  ua1=2.327791832e-08 lua1=-4.563842027e-15 wua1=-3.725325753e-14 pua1=7.581782972e-21
+  ub1=-2.405242424e-17 lub1=4.799667964e-24 wub1=3.917823309e-23 pub1=-7.973553998e-30
+  uc1=-2.230479155e-09 luc1=4.486024797e-16 wuc1=3.661805910e-15 puc1=-7.452507387e-22
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.1e-6
+  sbref=1.1e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.44 pmos
* Model Flag Parameters
+  lmin=1.5e-07 lmax=1.8e-07 wmin=1.68e-06 wmax=2.0e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-2.026e-8
+  vth0={-1.224871589e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=3.228227414e-08 wvth0=2.996292390e-07 pvth0=-6.607423978e-14
+  k1=2.797653987e-01 lk1=1.503202932e-07 wk1=-2.115610842e-07 pk1=4.665345028e-14
+  k2=1.283850377e-01 lk2=-6.403700226e-08 wk2=1.109939853e-07 pk2=-2.447639364e-14
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=2.414027790e+00 ldsub=-4.083422614e-07 wdsub=-2.653342159e-07 pdsub=5.851150130e-14
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-1.912617931e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=3.413572381e-07 wvoff=2.616390055e-06 pvoff=-5.769663349e-13
+  nfactor={7.939716180e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.140846779e-06 wnfactor=-6.219884113e-06 pnfactor=1.371608845e-12
+  eta0=-2.894334393e-02 leta0=1.144373862e-07 weta0=4.425650273e-06 peta0=-9.759443981e-13
+  etab=-1.484481651e+00 letab=3.272200687e-07 wetab=2.937639802e-06 petab=-6.478083292e-13
+  u0=3.520255316e-02 lu0=-6.935184885e-09 wu0=-5.699732206e-08 pu0=1.256904946e-14
+  ua=1.128551715e-08 lua=-2.951677342e-15 wua=-2.499600261e-14 pua=5.512118496e-21
+  ub=-9.137699022e-18 lub=2.425579670e-24 wub=2.125492576e-23 pub=-4.687136229e-30
+  uc=-6.568264105e-11 luc=1.264860536e-17 wuc=1.322890868e-16 puc=-2.917238943e-23
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=8.698934900e+05 lvsat=-1.649845719e-01 wvsat=-8.050385919e-01 pvsat=1.775271103e-7
+  a0=-8.285801497e+00 la0=1.994361158e-06 wa0=1.612845715e-05 pa0=-3.556647371e-12
+  ags=1.249999799e+00 lags=3.820406569e-14
+  a1=0.0
+  a2=-2.017380650e+00 la2=5.910498591e-07 wa2=4.074980592e-06 pa2=-8.986147202e-13
+  b0=6.947626328e-23 lb0=-1.532090558e-29 wb0=-1.376513751e-28 pb0=3.035488124e-35
+  b1=0.0
+  keta=-7.038732374e-01 lketa=1.391086993e-07 wketa=4.644982437e-07 pketa=-1.024311527e-13
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=2.659451529e+00 lpclm=-4.244483197e-07 wpclm=-2.479090907e-06 ppclm=5.466891268e-13
+  pdiblc1=2.566595050e+00 lpdiblc1=-4.642075173e-07 wpdiblc1=-3.799054459e-07 ppdiblc1=8.377674893e-14
+  pdiblc2=6.707207329e-02 lpdiblc2=-1.261212498e-08 wpdiblc2=-3.308028028e-08 ppdiblc2=7.294863408e-15
+  pdiblcb=4.066413726e+01 lpdiblcb=-9.016787941e-06 wpdiblcb=-6.950582134e-05 ppdiblcb=1.532742372e-11
+  drout=-1.319768868e+00 ldrout=4.419622965e-07 wdrout=-3.774175028e-12 pdrout=8.322810761e-19
+  pscbe1=7.876846413e+08 lpscbe1=2.715783011e+00 wpscbe1=2.440008288e+01 ppscbe1=-5.380706277e-6
+  pscbe2=-4.116811368e-08 lpscbe2=1.113363478e-14 wpscbe2=1.002807870e-13 ppscbe2=-2.211391916e-20
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=2.181320232e+01 lbeta0=-2.837388423e-06 wbeta0=-1.408126234e-05 pbeta0=3.105199971e-12
* Gidl Induced Drain Leakage Model Parameters
+  agidl=1.329003043e-14 lagidl=-2.923862667e-21 wagidl=-2.169876345e-20 pagidl=4.785011316e-27
+  bgidl=9.999998191e+08 lbgidl=3.446073341e-5
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-1.106e-8
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=2.783463815e+00 lkt1=-6.941360542e-07 wkt1=-1.525899513e-06 pkt1=3.364913606e-13
+  kt2=-2.117284491e-02 lkt2=-6.090575968e-09 wkt2=-1.695087293e-13 pkt2=3.738006504e-20
+  at=2.087262877e+05 lat=-4.385170120e-02 wat=-5.349809282e-01 pat=1.179739943e-7
+  ute=1.624822074e+00 lute=-3.627161636e-07 wute=9.942867174e-13 pute=-2.192601080e-19
+  ua1=5.596685055e-09 lua1=-1.045993618e-15 wua1=-3.919274349e-15 pua1=8.642783794e-22
+  ub1=-2.548359675e-18 lub1=4.585073066e-25 wub1=1.734858761e-30 pub1=-3.825710544e-37
+  uc1=-8.905018881e-10 luc1=1.905824016e-16 wuc1=1.711415570e-15 puc1=-3.774013614e-22
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.04e-6
+  sbref=1.04e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.45 pmos
* Model Flag Parameters
+  lmin=2.0e-05 lmax=0.0001 wmin=1.65e-06 wmax=1.68e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.112338352e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=8.389324645e-7
+  k1=4.212382248e-01 lk1=1.294361886e-6
+  k2=3.920842634e-02 lk2=-5.229813104e-7
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.478613255e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=1.269265013e-06 wvoff=3.552713679e-21
+  nfactor={4.403855138e-01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=4.140710528e-5
+  eta0=0.08
+  etab=-0.07
+  u0=9.352307657e-03 lu0=-2.323062827e-8
+  ua=-9.617482694e-10 lua=1.359202704e-14
+  ub=1.301805738e-18 lub=-2.210428646e-23
+  uc=-7.213676046e-11 luc=-7.421843743e-16
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=160312.5
+  a0=1.663147057e+00 la0=4.626521022e-8
+  ags=5.520619633e-01 lags=-2.963429165e-6
+  a1=0.0
+  a2=0.8
+  b0=0.0
+  b1=0.0
+  keta=-5.481114733e-02 lketa=4.720579346e-7
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=2.043221610e-01 lpclm=-2.886910939e-6
+  pdiblc1=0.39
+  pdiblc2=1.362013555e-04 lpdiblc2=3.019310429e-9
+  pdiblcb=-3.449469752e-03 lpdiblcb=3.842808139e-8
+  drout=0.56
+  pscbe1=7.008429116e+08 lpscbe1=1.790436848e+3
+  pscbe2=9.666085849e-09 lpscbe2=-6.118193515e-15
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=5.682944295e-10 lalpha0=-9.376902874e-15
+  alpha1=-2.468523241e-11 lalpha1=2.496637245e-15 walpha1=-3.231174268e-32 palpha1=1.096014312e-35
+  beta0=3.268541021e+00 lbeta0=-5.377136505e-6
* Gidl Induced Drain Leakage Model Parameters
+  agidl=6.249611638e-10 lagidl=-1.163385201e-14
+  bgidl=1.563144045e+09 lbgidl=-1.127612605e+4
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-3.006910881e-01 lkt1=-3.100620284e-6
+  kt2=-0.037961
+  at=0.0
+  ute=-3.559961858e-01 lute=5.267424367e-7
+  ua1=2.139640475e-09 lua1=7.197644988e-15
+  ub1=-7.302764894e-19 lub1=-1.903282652e-23 wub1=1.232595164e-38
+  uc1=4.325252718e-11 luc1=7.661548855e-15
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.46 pmos
* Model Flag Parameters
+  lmin=8.0e-06 lmax=2.0e-05 wmin=1.65e-06 wmax=1.68e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.070441+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+  k1=0.4858803
+  k2=0.013090076
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-0.18447262+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={2.5083089+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+  eta0=0.08
+  etab=-0.07
+  u0=0.0081921406
+  ua=-2.8294519e-10
+  ub=1.9788962e-19
+  uc=-1.0920239e-10
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=160312.5
+  a0=1.6654576
+  ags=0.40406455
+  a1=0.0
+  a2=0.8
+  b0=0.0
+  b1=0.0
+  keta=-0.031235975
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=0.060146165
+  pdiblc1=0.39
+  pdiblc2=0.00028698955
+  pdiblcb=-0.0015303226
+  drout=0.56
+  pscbe1=790259600.0
+  pscbe2=9.3605355e-9
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=3.0
* Gidl Induced Drain Leakage Model Parameters
+  agidl=4.395183e-11
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-0.45554
+  kt2=-0.037961
+  at=0.0
+  ute=-0.32969
+  ua1=2.4991e-9
+  ub1=-1.6808e-18
+  uc1=4.2588e-10
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.47 pmos
* Model Flag Parameters
+  lmin=4.0e-06 lmax=8.0e-06 wmin=1.65e-06 wmax=1.68e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.084602080e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=1.136217118e-7
+  k1=4.520055508e-01 lk1=2.717947275e-7
+  k2=2.140616637e-02 lk2=-6.672431739e-8
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-1.911172420e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=5.331325740e-8
+  nfactor={2.706977945e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.594025058e-6
+  eta0=0.08
+  etab=-0.07
+  u0=1.046272419e-02 lu0=-1.821807282e-8
+  ua=3.775496570e-10 lua=-5.299493615e-15 pua=2.646977960e-35
+  ub=-2.359133808e-19 lub=3.480627053e-24
+  uc=-1.426185303e-10 luc=2.681150701e-16
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=2.217873591e+05 lvsat=-4.932447618e-01 wvsat=3.725290298e-15
+  a0=1.702304594e+00 la0=-2.956425918e-7
+  ags=4.037452334e-01 lags=2.562043175e-9
+  a1=0.0
+  a2=0.8
+  b0=0.0
+  b1=0.0
+  keta=-3.748950581e-02 lketa=5.017532955e-8
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-5.158874480e-01 lpclm=4.621817215e-06 ppclm=2.842170943e-26
+  pdiblc1=0.39
+  pdiblc2=3.594023986e-04 lpdiblc2=-5.810059386e-10
+  pdiblcb=-4.365230551e-04 lpdiblcb=-8.776122525e-9
+  drout=0.56
+  pscbe1=7.804619264e+08 lpscbe1=7.861182970e+1
+  pscbe2=9.151205032e-09 lpscbe2=1.679567196e-15
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=-7.139407148e-01 lbeta0=2.979887760e-5
* Gidl Induced Drain Leakage Model Parameters
+  agidl=-8.863176868e-12 lagidl=4.237622639e-16
+  bgidl=8.005398301e+08 lbgidl=1.600372662e+3
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-5.106119300e-01 lkt1=4.418707318e-7
+  kt2=-3.133225080e-02 lkt2=-5.318590178e-8
+  at=-1.804649308e+05 lat=1.447963982e+0
+  ute=1.659976052e-01 lute=-3.977159414e-6
+  ua1=5.352670913e-09 lua1=-2.289568329e-14 wua1=5.293955920e-29
+  ub1=-4.246608763e-18 lub1=2.058681792e-23 pub1=-1.972152263e-43
+  uc1=7.932676112e-10 luc1=-2.947741846e-15
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.48 pmos
* Model Flag Parameters
+  lmin=2.0e-06 lmax=4.0e-06 wmin=1.65e-06 wmax=1.68e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.030249984e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-1.050650359e-7
+  k1=5.991182345e-01 lk1=-3.201160977e-7
+  k2=-1.299424793e-02 lk2=7.168643753e-08 pk2=-2.220446049e-28
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-1.421224013e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-1.438184639e-7
+  nfactor={3.189571823e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-3.535751178e-6
+  eta0=0.08
+  etab=-0.07
+  u0=3.422457921e-03 lu0=1.010857931e-8
+  ua=-1.459651534e-09 lua=2.092522121e-15
+  ub=8.652439039e-19 lub=-9.499013051e-25
+  uc=-6.679231726e-11 luc=-3.697321461e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=1.454941258e+05 lvsat=-1.862774118e-1
+  a0=2.092775327e+00 la0=-1.866709395e-6
+  ags=4.703125816e-01 lags=-2.652730136e-7
+  a1=0.0
+  a2=0.8
+  b0=0.0
+  b1=0.0
+  keta=-4.146445057e-02 lketa=6.616859927e-8
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=9.388625344e-01 lpclm=-1.231398434e-6
+  pdiblc1=0.39
+  pdiblc2=0.000215
+  pdiblcb=2.002775912e-02 lpdiblcb=-9.111457113e-08 wpdiblcb=-5.551115123e-23 ppdiblcb=3.330669074e-28
+  drout=0.56
+  pscbe1=800000000.0
+  pscbe2=1.684351014e-08 lpscbe2=-2.927057626e-14
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=5.546325391e+00 lbeta0=4.610571722e-6
* Gidl Induced Drain Leakage Model Parameters
+  agidl=1.035556976e-10 lagidl=-2.855732580e-17
+  bgidl=1.142050664e+09 lbgidl=2.262969922e+2
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-3.424855594e-01 lkt1=-2.345890828e-7
+  kt2=-4.009733871e-02 lkt2=-1.791939525e-8
+  at=2.762557340e+05 lat=-3.896607476e-1
+  ute=-1.654632365e+00 lute=3.348181683e-6
+  ua1=-3.325705164e-09 lua1=1.202193642e-14 wua1=1.323488980e-29
+  ub1=3.210225146e-18 lub1=-9.415902443e-24 wub1=-2.465190329e-38 pub1=-4.930380658e-44
+  uc1=9.271368235e-11 luc1=-1.290491024e-16
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.49 pmos
* Model Flag Parameters
+  lmin=1.0e-06 lmax=2.0e-06 wmin=1.65e-06 wmax=1.68e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.087180700e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=1.013540662e-8
+  k1=4.319945642e-01 lk1=1.806199173e-8
+  k2=2.626747013e-02 lk2=-7.760434200e-9
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=3.857674493e-01 ldsub=3.525630509e-7
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.218714828e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=1.755539745e-8
+  nfactor={1.091537207e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=7.096638280e-7
+  eta0=-6.226469463e-02 leta0=2.878754549e-7
+  etab=7.107223768e-01 letab=-1.579807344e-06 wetab=-1.776356839e-21 petab=-7.105427358e-27
+  u0=8.370467731e-03 lu0=9.618249656e-11
+  ua=-5.360904043e-11 lua=-7.526329856e-16
+  ub=-1.474362962e-19 lub=1.099277333e-24
+  uc=-1.227185167e-10 luc=7.619456839e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=3.992446544e+04 lvsat=2.734490745e-2
+  a0=1.180300103e+00 la0=-2.029753060e-8
+  ags=6.547809364e-02 lags=5.539176694e-7
+  a1=0.0
+  a2=0.8
+  b0=0.0
+  b1=0.0
+  keta=-2.414474864e-03 lketa=-1.284980757e-8
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=3.094768240e-02 lpclm=6.057854269e-7
+  pdiblc1=4.094634917e-01 lpdiblc1=-3.938476478e-8
+  pdiblc2=-5.056800000e-06 lpdiblc2=4.452893359e-10
+  pdiblcb=-0.025
+  drout=1.194940541e-01 ldrout=8.913725917e-7
+  pscbe1=800000000.0
+  pscbe2=-4.693562463e-09 lpscbe2=1.431012090e-14 ppscbe2=5.293955920e-35
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=6.758248586e+00 lbeta0=2.158220897e-6
* Gidl Induced Drain Leakage Model Parameters
+  agidl=9.805489728e-11 lagidl=-1.742634638e-17
+  bgidl=1.269621336e+09 lbgidl=-3.184481508e+1
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.439715564e-01 lkt1=-2.923013823e-8
+  kt2=-6.080719617e-02 lkt2=2.398741550e-8
+  at=6.427369205e+04 lat=3.928915392e-2
+  ute=0.0
+  ua1=2.831661075e-09 lua1=-4.376173113e-16
+  ub1=-1.530007496e-18 lub1=1.760531127e-25
+  uc1=1.571903929e-10 luc1=-2.595190157e-16 wuc1=8.271806126e-31 puc1=8.271806126e-37
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=2.75e-6
+  sbref=2.74e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.50 pmos
* Model Flag Parameters
+  lmin=5.0e-07 lmax=1.0e-06 wmin=1.65e-06 wmax=1.68e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.111696813e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=3.522813877e-8
+  k1=3.245759539e-01 lk1=1.280070877e-7
+  k2=5.361238178e-02 lk2=-3.574849817e-8
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=4.477675013e-01 ldsub=2.891047577e-7
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.206309585e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=1.628569604e-8
+  nfactor={5.391600791e-01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.275032866e-6
+  eta0=3.681232431e-01 leta0=-1.526352071e-7
+  etab=-1.704214254e+00 letab=8.919285964e-7
+  u0=1.143362200e-02 lu0=-3.039017162e-9
+  ua=-2.679092862e-10 lua=-5.332923980e-16
+  ub=7.860221385e-19 lub=1.438639564e-25
+  uc=-6.535283089e-11 luc=1.747964170e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=5.000039328e+04 lvsat=1.703199379e-2
+  a0=1.139495742e+00 la0=2.146654927e-8
+  ags=-6.996480032e-02 lags=6.925461803e-7
+  a1=0.0
+  a2=5.906024704e-01 la2=2.143225595e-7
+  b0=0.0
+  b1=0.0
+  keta=1.852895072e-02 lketa=-3.428582252e-08 pketa=2.220446049e-28
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=5.318634040e-01 lpclm=9.308816755e-8
+  pdiblc1=-2.876213835e-01 lpdiblc1=6.740955467e-7
+  pdiblc2=-1.851964142e-04 lpdiblc2=6.296658339e-10
+  pdiblcb=-5.082653338e-02 lpdiblcb=2.643397344e-8
+  drout=1.010442376e+00 ldrout=-2.053083449e-8
+  pscbe1=8.091570768e+08 lpscbe1=-9.372451233e+0
+  pscbe2=9.340256864e-09 lpscbe2=-5.377386132e-17
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=8.432376873e+00 lbeta0=4.447171140e-7
* Gidl Induced Drain Leakage Model Parameters
+  agidl=1.232393706e-10 lagidl=-4.320315848e-17
+  bgidl=1.283381922e+09 lbgidl=-4.592904908e+1
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.527514144e-01 lkt1=-2.024377793e-8
+  kt2=-2.665978080e-02 lkt2=-1.096314708e-8
+  at=1.735027264e+05 lat=-7.250894732e-2
+  ute=2.094080000e-02 lute=-2.143332762e-8
+  ua1=2.668791712e-09 lua1=-2.709172611e-16
+  ub1=-1.027554176e-18 lub1=-3.382179098e-25
+  uc1=-1.237272963e-10 luc1=2.800585753e-17
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.75e-6
+  sbref=1.74e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.51 pmos
* Model Flag Parameters
+  lmin=2.5e-07 lmax=5.0e-07 wmin=1.65e-06 wmax=1.68e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.007126113e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-1.951671385e-8
+  k1=1.398369388e-01 lk1=2.247216569e-7
+  k2=1.465220025e-01 lk2=-8.438854283e-08 pk2=3.330669074e-28
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=1.478875091e+00 ldsub=-2.507006874e-07 wdsub=2.842170943e-20
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={2.083403189e-03+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-1.003097266e-7
+  nfactor={3.202647319e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.193559734e-7
+  eta0=-3.757605076e-01 leta0=2.368028140e-07 weta0=1.776356839e-21 peta0=1.332267630e-27
+  etab=-3.627991333e-04 letab=-7.171718105e-11
+  u0=7.680418113e-03 lu0=-1.074139862e-9
+  ua=-3.971058257e-10 lua=-4.656554257e-16
+  ub=1.846390384e-19 lub=4.587000370e-25
+  uc=-5.782776129e-11 luc=1.354011726e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=3.964825290e+04 lvsat=2.245154632e-2
+  a0=1.642639393e+00 la0=-2.419392149e-7
+  ags=1.256072862e+00 lags=-1.661056634e-9
+  a1=0.0
+  a2=1.368821359e+00 la2=-1.930905928e-7
+  b0=0.0
+  b1=0.0
+  keta=-1.841745284e-02 lketa=-1.494364133e-8
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=6.823070923e-01 lpclm=1.432788787e-8
+  pdiblc1=1.589122175e+00 lpdiblc1=-3.084172413e-7
+  pdiblc2=-8.678023286e-03 lpdiblc2=5.075830558e-09 ppdiblc2=6.938893904e-30
+  pdiblcb=2.450492987e-01 lpdiblcb=-1.284629422e-07 wpdiblcb=1.249000903e-22 ppdiblcb=7.077671782e-28
+  drout=1.285020706e+00 ldrout=-1.642780821e-7
+  pscbe1=7.816858459e+08 lpscbe1=5.009287583e+0
+  pscbe2=9.147344128e-09 lpscbe2=4.721981420e-17
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=9.648868735e+00 lbeta0=-1.921407060e-7
* Gidl Induced Drain Leakage Model Parameters
+  agidl=8.526043319e-11 lagidl=-2.332042518e-17
+  bgidl=1.409708245e+09 lbgidl=-1.120634058e+2
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.00074326333
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.5407449e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-6.305432205e-01 lkt1=7.283378841e-8
+  kt2=-4.629795127e-02 lkt2=-6.821720693e-10
+  at=6.249379701e+04 lat=-1.439355261e-2
+  ute=-2.000000091e-02 lute=4.782112484e-16
+  ua1=3.571328252e-09 lua1=-7.434131907e-16
+  ub1=-2.991364602e-18 lub1=6.898761243e-25
+  uc1=-1.183397965e-10 luc1=2.518539364e-17
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.1e-6
+  sbref=1.1e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.52 pmos
* Model Flag Parameters
+  lmin=1.8e-07 lmax=2.5e-07 wmin=1.65e-06 wmax=1.68e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.07847999562893+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+  k1=0.961428255393082
+  k2=-0.162005866831761
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.562303405039308
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-0.364652947389937+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={2.7662771322327+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+  eta0=0.49
+  etab=-0.000625
+  u0=0.0037533200490566
+  ua=-2.09956058459119e-9
+  ub=1.86166461966667e-18
+  uc=-8.324553995283e-12
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=121731.999327042
+  a0=0.758099999261006
+  ags=1.24999997272013
+  a1=0.0
+  a2=0.662874470440252
+  b0=0.0
+  b1=0.0
+  keta=-0.0730519999606918
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=0.734690420259434
+  pdiblc1=0.461536473183962
+  pdiblc2=0.00987941513820755
+  pdiblcb=-0.224616327814465
+  drout=0.684413503600629
+  pscbe1=800000000.518868
+  pscbe2=9.31998164677673e-9
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=8.94639467130503
* Gidl Induced Drain Leakage Model Parameters
+  agidl=3.10849060300319e-17
+  bgidl=999999975.393082
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.00074326333
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.5407449e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-0.364259992940252
+  kt2=-0.0487919994941038
+  at=9870.39612421382
+  ute=-0.0199999991650943
+  ua1=8.53380055896226e-10
+  ub1=-4.69150049528303e-19
+  uc1=-2.62609955581761e-11
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.1e-6
+  sbref=1.1e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.53 pmos
* Model Flag Parameters
+  lmin=1.5e-07 lmax=1.8e-07 wmin=1.65e-06 wmax=1.68e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-2.026e-8
+  vth0={-1.044505083e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-7.492147672e-09 wvth0=-8.586443073e-12 pvth0=1.893482420e-18
+  k1=1.524197065e-01 lk1=1.784025652e-07 wk1=-5.251349080e-12 pk1=1.158027487e-18
+  k2=1.952029349e-01 lk2=-7.877168496e-08 wk2=-8.716520838e-12 pk2=1.922167172e-18
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=2.254289871e+00 ldsub=-3.731168554e-07 wdsub=3.391698669e-11 pdsub=-7.479373906e-18
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-3.376856205e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-5.946834926e-09 wvoff=-8.936935103e-13 pvoff=1.970772914e-19
+  nfactor={4.195659245e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-3.152073436e-07 wnfactor=1.283810775e-11 pnfactor=-2.831059476e-18
+  eta0=2.635060538e+00 leta0=-4.730287498e-07 weta0=1.521567049e-11 peta0=-3.355359652e-18
+  etab=2.838279318e-01 letab=-6.272756051e-08 wetab=-3.395191542e-12 petab=7.487076384e-19
+  u0=8.930942449e-04 lu0=6.307369943e-10 wu0=2.136794119e-14 pu0=-4.712058299e-21
+  ua=-3.760773494e-09 lua=3.663306708e-16 wua=-2.125834015e-20 pua=4.687889182e-27
+  ub=3.656686821e-18 lub=-3.958382958e-25 wub=-2.919559084e-29 pub=6.438211660e-36
+  uc=1.394852754e-11 luc=-4.911659940e-18 wuc=5.612683334e-23 puc=-1.237708924e-29
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=3.853015113e+05 lvsat=-5.812234877e-02 wvsat=4.938202649e-07 pvsat=-1.088972464e-13
+  a0=1.422694474e+00 la0=-1.465563736e-07 wa0=4.629861508e-12 pa0=-1.020977066e-18
+  ags=1.249999799e+00 lags=3.820404970e-14
+  a1=0.0
+  a2=4.355362553e-01 la2=5.013262320e-08 wa2=1.841947699e-11 pa2=-4.061863066e-18
+  b0=-1.338267830e-23 lb0=2.951148219e-30 wb0=-1.354993220e-34 pb0=2.988031046e-41
+  b1=0.0
+  keta=-4.242675334e-01 lketa=7.745004943e-08 wketa=-2.883425651e-12 pketa=6.358530253e-19
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=1.167168806e+00 lpclm=-9.537013359e-08 wpclm=-3.402900120e-12 ppclm=7.504075370e-19
+  pdiblc1=2.337921697e+00 lpdiblc1=-4.137804696e-07 wpdiblc1=-1.680793832e-11 ppdiblc1=3.706486559e-18
+  pdiblc2=4.715932866e-02 lpdiblc2=-8.220966529e-09 wpdiblc2=2.048147554e-13 ppdiblc2=-4.516574958e-20
+  pdiblcb=-1.174780210e+00 lpdiblcb=2.095301394e-07 wpdiblcb=7.587962898e-13 ppdiblcb=-1.673297589e-19
+  drout=-1.319791092e+00 ldrout=4.419671974e-07 wdrout=3.314614605e-11 pdrout=-7.309388124e-18
+  pscbe1=8.023713568e+08 lpscbe1=-5.229314770e-01 wpscbe1=1.453757080e-03 ppscbe1=-3.205825195e-10
+  pscbe2=1.919566468e-08 lpscbe2=-2.177785623e-15 wpscbe2=1.322232474e-19 ppscbe2=-2.915787064e-26
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=1.333702501e+01 lbeta0=-9.682218024e-07 wbeta0=-2.630252402e-11 pbeta0=5.800232657e-18
* Gidl Induced Drain Leakage Model Parameters
+  agidl=-5.919330646e-14 lagidl=1.306016278e-20 wagidl=9.871577459e-20 pagidl=-2.176880261e-26
+  bgidl=9.999998191e+08 lbgidl=3.446073914e-5
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-1.106e-8
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.00074326333
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.5407449e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=1.864927527e+00 lkt1=-4.915804319e-07 wkt1=3.910329821e-11 pkt1=-8.623059315e-18
+  kt2=-2.117384306e-02 lkt2=-6.090355857e-09 wkt2=1.488685889e-12 pkt2=-3.282850116e-19
+  at=-1.133031594e+05 lat=2.716223247e-02 wat=-2.424534562e-06 pat=5.346583610e-13
+  ute=1.624827929e+00 lute=-3.627174547e-07 wute=-8.732179245e-12 pute=1.925620172e-18
+  ua1=3.237480574e-09 lua1=-5.257418462e-16 wua1=5.998103409e-21 pua1=-1.322701742e-27
+  ub1=-2.548349459e-18 lub1=4.585050539e-25 wub1=-1.523614605e-29 pub1=3.359874940e-36
+  uc1=1.396802315e-10 luc1=-3.659335939e-17 wuc1=2.859336849e-21 puc1=-6.305409626e-28
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.04e-6
+  sbref=1.04e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.54 pmos
* Model Flag Parameters
+  lmin=2.0e-05 lmax=0.0001 wmin=1.26e-06 wmax=1.65e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.259834082e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=4.924075150e-06 wvth0=2.406056551e-07 pvth0=-6.663978880e-12
+  k1=1.849382087e-01 lk1=8.470762697e-06 wk1=3.854695997e-07 pk1=-1.170666170e-11
+  k2=1.286259373e-01 lk2=-2.816583826e-06 wk2=-1.458642820e-07 pk2=3.741489562e-12
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-4.715644232e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=7.504810579e-06 wvoff=3.649205995e-07 pvoff=-1.017187089e-11
+  nfactor={-6.693837421e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=2.284627552e-04 wnfactor=1.163785812e-05 pnfactor=-3.051386441e-10
+  eta0=0.08
+  etab=-0.07
+  u0=1.370360267e-02 lu0=-1.630608552e-07 wu0=-7.098145722e-09 pu0=2.281011339e-13
+  ua=-3.475725128e-09 lua=9.221207121e-14 wua=4.100980059e-15 pua=-1.282506767e-19
+  ub=5.442539477e-18 lub=-1.551960419e-22 wub=-6.754663009e-24 pub=2.171088540e-28
+  uc=7.564781992e-11 luc=-6.086471515e-15 wuc=-2.410768480e-16 puc=8.717985972e-21
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=1.603105084e+05 lvsat=1.992025683e-04 wvsat=3.248771609e-06 pvsat=-3.249535720e-10
+  a0=1.326867898e+00 la0=3.309378006e-05 wa0=5.485627757e-07 pa0=-5.390948565e-11
+  ags=8.927781713e-01 lags=6.400225870e-07 wags=-5.558008100e-07 pags=-5.878209947e-12
+  a1=0.0
+  a2=0.8
+  b0=0.0
+  b1=0.0
+  keta=-1.064515478e-01 lketa=-3.653953997e-07 wketa=8.423953930e-08 pketa=1.366114176e-12
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=7.275754670e-01 lpclm=-1.851447115e-05 wpclm=-8.535684670e-07 ppclm=2.549280140e-11
+  pdiblc1=0.39
+  pdiblc2=-3.179819101e-04 lpdiblc2=1.005464475e-08 wpdiblc2=7.408964440e-10 ppdiblc2=-1.147654388e-14
+  pdiblcb=-1.319103139e-01 lpdiblcb=1.239888084e-05 wpdiblcb=2.095545781e-07 ppdiblcb=-2.016326049e-11
+  drout=0.56
+  pscbe1=4.239726518e+08 lpscbe1=6.716706801e+03 wpscbe1=4.516507025e+02 ppscbe1=-8.036086239e-3
+  pscbe2=7.503806773e-09 lpscbe2=2.879597693e-13 wpscbe2=3.527265313e-15 ppscbe2=-4.797211465e-19
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=2.058757924e-09 lalpha0=-3.922122847e-14 walpha0=-2.431351366e-15 palpha0=4.868421271e-20
+  alpha1=-4.215269960e-10 lalpha1=1.044280624e-14 walpha1=6.473568574e-16 palpha1=-1.296236298e-20
+  beta0=6.735038952e+00 lbeta0=-2.837325744e-04 wbeta0=-5.654801013e-06 pbeta0=4.540734320e-10
* Gidl Induced Drain Leakage Model Parameters
+  agidl=1.282878866e-08 lagidl=-1.084367098e-12 wagidl=-1.990776208e-14 pagidl=1.749919708e-18
+  bgidl=3.355490034e+09 lbgidl=-4.716520180e+04 wbgidl=-2.923803825e+03 pbgidl=5.854484437e-2
+  cgidl=300.0
+  egidl=7.257071840e-01 legidl=-6.258543503e-05 wegidl=-1.020698609e-06 pegidl=1.020938678e-10
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=2.039190131e-01 lkt1=-1.414588477e-05 wkt1=-8.231563291e-07 pkt1=1.801783069e-11
+  kt2=-4.943035601e-02 lkt2=1.147205360e-06 wkt2=1.870963931e-08 pkt2=-1.871403982e-12
+  at=0.0
+  ute=-2.824497794e-01 lute=-1.352770633e-05 wute=-1.199741933e-07 pute=2.292662874e-11
+  ua1=4.567547559e-10 lua1=8.400025098e-14 wua1=2.745244353e-15 pua1=-1.252859407e-19
+  ub1=3.063671297e-18 lub1=-1.564946401e-22 wub1=-6.188960794e-24 pub1=2.242376075e-28
+  uc1=-1.520799765e-09 luc1=6.667899670e-14 wuc1=2.551394711e-15 puc1=-9.627351018e-20
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.55 pmos
* Model Flag Parameters
+  lmin=8.0e-06 lmax=2.0e-05 wmin=1.26e-06 wmax=1.65e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.013919520e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} wvth0=-9.220190716e-8
+  k1=6.079788478e-01 wk1=-1.991759423e-7
+  k2=-1.203783334e-02 wk2=4.099045493e-8
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-9.676465875e-02+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} wvoff=-1.430755414e-7
+  nfactor={4.715882507e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} wnfactor=-3.601153013e-6
+  eta0=0.08
+  etab=-0.07
+  u0=5.560136630e-03 wu0=4.293514380e-9
+  ua=1.129462731e-09 wua=-2.304021494e-15
+  ub=-2.308147808e-18 wub=4.088028687e-24
+  uc=-2.283182917e-10 wuc=1.943104352e-16
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=1.603204569e+05 wvsat=-1.297982217e-5
+  a0=2.979613273e+00 wa0=-2.143745352e-6
+  ags=9.247417115e-01 wags=-8.493660746e-7
+  a1=0.0
+  a2=0.8
+  b0=0.0
+  b1=0.0
+  keta=-1.246998577e-01 wketa=1.524650149e-7
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-1.970607183e-01 wpclm=4.195743870e-7
+  pdiblc1=0.39
+  pdiblc2=1.841598085e-04 wpdiblc2=1.677432780e-10
+  pdiblcb=4.873055303e-01 wpdiblcb=-7.974242395e-7
+  drout=0.56
+  pscbe1=7.594135134e+08 wpscbe1=5.031835740e+1
+  pscbe2=2.188488309e-08 wpscbe2=-2.043061754e-14
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=-7.434925891e+00 wbeta0=1.702220243e-5
* Gidl Induced Drain Leakage Model Parameters
+  agidl=-4.132588037e-08 wagidl=6.748544891e-14
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=-2.399888867e+00 wegidl=4.077998711e-6
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-5.025444244e-01 wkt1=7.667700147e-8
+  kt2=7.862535550e-03 wkt2=-7.475065048e-8
+  at=0.0
+  ute=-9.580406010e-01 wute=1.025010742e-6
+  ua1=4.651833892e-09 wua1=-3.511694522e-15
+  ub1=-4.751869630e-18 wub1=5.009749898e-24
+  uc1=1.809233950e-09 wuc1=-2.256626565e-15
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.56 pmos
* Model Flag Parameters
+  lmin=4.0e-06 lmax=8.0e-06 wmin=1.26e-06 wmax=1.65e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.066103100e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=4.186959914e-07 wvth0=-3.017686951e-08 pvth0=-4.976591301e-13
+  k1=4.403333565e-01 lk1=1.345106952e-06 wk1=1.904052371e-08 pk1=-1.750864179e-12
+  k2=2.952911439e-02 lk2=-3.335132364e-07 wk2=-1.325073766e-08 pk2=4.352052936e-13
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-1.446182280e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=3.839540695e-07 wvoff=-7.585253962e-08 pvoff=-5.393650989e-13
+  nfactor={4.478956937e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.900977052e-06 wnfactor=-2.890579714e-06 pnfactor=-5.701299081e-12
+  eta0=0.08
+  etab=-0.07
+  u0=1.659636061e-02 lu0=-8.854936386e-08 wu0=-1.000562936e-08 pu0=1.147294658e-13
+  ua=4.201103791e-09 lua=-2.464537348e-14 wua=-6.237256800e-15 pua=3.155839214e-20
+  ub=-4.323937849e-18 lub=1.617373171e-23 wub=6.668679851e-24 pub=-2.070590623e-29
+  uc=-3.710778556e-10 luc=1.145434216e-15 wuc=3.726793004e-16 puc=-1.431146158e-21
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=7.530756142e+04 lvsat=6.821026669e-01 wvsat=2.389483926e-01 pvsat=-1.917311351e-6
+  a0=2.833037550e+00 la0=1.176053241e-06 wa0=-1.844533011e-06 pa0=-2.400736205e-12
+  ags=1.025174205e+00 lags=-8.058221213e-07 wags=-1.013719682e-06 pags=1.318694453e-12
+  a1=0.0
+  a2=0.8
+  b0=0.0
+  b1=0.0
+  keta=-1.541469495e-01 lketa=2.362693300e-07 wketa=1.903000215e-07 pketa=-3.035699324e-13
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-2.923957431e+00 lpclm=2.187931031e-05 wpclm=3.928217137e-06 ppclm=-2.815166528e-11
+  pdiblc1=0.39
+  pdiblc2=5.951723013e-03 lpdiblc2=-4.627615873e-08 wpdiblc2=-9.122596034e-09 ppdiblc2=7.454122328e-14
+  pdiblcb=7.919560869e-01 lpdiblcb=-2.444369834e-06 wpdiblcb=-1.292607878e-06 ppdiblcb=3.973115824e-12
+  drout=0.56
+  pscbe1=-6.414330815e+08 lpscbe1=1.123972067e+04 wpscbe1=2.319497513e+03 ppscbe1=-1.820680434e-2
+  pscbe2=9.275311625e-08 lpscbe2=-5.686126861e-13 wpscbe2=-1.363774569e-13 ppscbe2=9.303017846e-19
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=-1.390171428e+01 lbeta0=5.188640597e-05 wbeta0=2.151284576e-05 pbeta0=-3.603076657e-11
* Gidl Induced Drain Leakage Model Parameters
+  agidl=-8.320932716e-08 lagidl=3.360526730e-13 wagidl=1.357225873e-13 pagidl=-5.475020444e-19
+  bgidl=1.657082301e+08 lbgidl=6.693956702e+03 wbgidl=1.035583014e+03 pbgidl=-8.309021023e-3
+  cgidl=300.0
+  egidl=-4.914477080e+00 legidl=2.017584882e-05 wegidl=8.179976055e-06 pegidl=-3.291229726e-11
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-8.432140915e-01 lkt1=2.733369887e-06 wkt1=5.425645932e-07 pkt1=-3.738058410e-12
+  kt2=2.296706914e-02 lkt2=-1.211915274e-07 wkt2=-8.857696024e-08 pkt2=1.109356729e-13
+  at=-4.645435735e+05 lat=3.727274653e+00 wat=4.634095357e-01 pat=-3.718175678e-6
+  ute=1.218594893e+00 lute=-1.746427842e-05 wute=-1.717072482e-06 pute=2.200115959e-11
+  ua1=2.057366811e-08 lua1=-1.277491552e-13 wua1=-2.482958653e-14 pua1=1.710445329e-19
+  ub1=-2.038483853e-17 lub1=1.254314387e-22 wub1=2.632584235e-23 pub1=-1.710300941e-28
+  uc1=3.355113400e-09 luc1=-1.240339468e-14 wuc1=-4.179067303e-15 puc1=1.542474171e-20
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.57 pmos
* Model Flag Parameters
+  lmin=2.0e-06 lmax=4.0e-06 wmin=1.26e-06 wmax=1.65e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-8.533107440e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-4.374783072e-07 wvth0=-2.886360277e-07 pvth0=5.422564619e-13
+  k1=1.096616803e+00 lk1=-1.295462621e-06 wk1=-8.115554849e-07 pk1=1.591055473e-12
+  k2=-1.241603561e-01 lk2=2.848594217e-07 wk2=1.813421596e-07 pk2=-3.477431202e-13
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=-4.018703740e-01 ldsub=3.870104687e-06 wdsub=1.569072209e-06 pdsub=-6.313193414e-12
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={1.496189449e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-7.999150802e-07 wvoff=-4.759094893e-07 pvoff=1.070272039e-12
+  nfactor={1.083263857e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-2.366318805e-05 wnfactor=-1.246792077e-05 pnfactor=3.283332421e-11
+  eta0=-1.760041385e-01 leta0=1.030037771e-06 weta0=4.176123830e-07 peta0=-1.680271775e-12
+  etab=1.538063815e-01 letab=-9.004894520e-07 wetab=-3.650890835e-07 petab=1.468943229e-12
+  u0=-1.318046748e-02 lu0=3.125829952e-08 wu0=2.708388733e-08 pu0=-3.450094639e-14
+  ua=-3.490524632e-09 lua=6.302047316e-15 wua=3.312906421e-15 pua=-6.866880585e-21
+  ub=3.997342179e-19 lub=-2.832057322e-24 wub=7.593729165e-25 pub=3.070308410e-30
+  uc=-3.874751442e-11 luc=-1.917035581e-16 wuc=-4.574870161e-17 puc=2.524072769e-22
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=4.384856423e+05 lvsat=-7.791516052e-01 wvsat=-4.779488571e-01 pvsat=9.671390713e-7
+  a0=5.080434371e+00 la0=-7.866392817e-06 wa0=-4.873684545e-06 pa0=9.787115574e-12
+  ags=1.495274687e+00 lags=-2.697280814e-06 wags=-1.671991984e-06 pags=3.967266228e-12
+  a1=0.0
+  a2=0.8
+  b0=0.0
+  b1=0.0
+  keta=-1.943725976e-01 lketa=3.981180297e-07 wketa=2.494347789e-07 pketa=-5.414998112e-13
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=5.696546538e+00 lpclm=-1.280545982e-05 wpclm=-7.761076700e-06 ppclm=1.888044226e-11
+  pdiblc1=0.39
+  pdiblc2=-1.068983124e-02 lpdiblc2=2.068146763e-08 wpdiblc2=1.778874586e-08 ppdiblc2=-3.373709907e-14
+  pdiblcb=3.963346606e-01 lpdiblcb=-8.525791124e-07 wpdiblcb=-6.138589118e-07 ppdiblcb=1.242155785e-12
+  drout=0.56
+  pscbe1=3.495055853e+09 lpscbe1=-5.403525286e+03 wpscbe1=-4.396369151e+03 ppscbe1=8.814619501e-3
+  pscbe2=-7.766053239e-08 lpscbe2=1.170500375e-13 wpscbe2=1.541617985e-13 ppscbe2=-2.386887202e-19
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=-1.331867141e+01 lbeta0=4.954052131e-05 wbeta0=3.077394106e-05 pbeta0=-7.329296873e-11
* Gidl Induced Drain Leakage Model Parameters
+  agidl=3.115143511e-10 lagidl=4.896746241e-18 wagidl=-3.392371287e-16 pagidl=-5.457269101e-23
+  bgidl=1.594162233e+09 lbgidl=9.465434538e+02 wbgidl=-7.375169427e+02 pbgidl=-1.174917886e-3
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=1.003259608e-01 lkt1=-1.062982384e-06 wkt1=-7.223460343e-07 pkt1=1.351334798e-12
+  kt2=2.415912399e-02 lkt2=-1.259877839e-07 wkt2=-1.048197684e-07 pkt2=1.762889365e-13
+  at=8.299288720e+05 lat=-1.481061121e+00 wat=-9.031914872e-01 pat=1.780370870e-6
+  ute=-6.498441236e+00 lute=1.358537079e-05 wute=7.901569785e-06 pute=-1.669963995e-11
+  ua1=-2.448900850e-08 lua1=5.356142534e-14 wua1=3.452310417e-14 pua1=-6.776220517e-20
+  ub1=2.247396535e-17 lub1=-4.701181596e-23 wub1=-3.142440002e-23 pub1=6.132916104e-29
+  uc1=3.299196164e-10 luc1=-2.314669889e-16 wuc1=-3.869473985e-16 puc1=1.670714305e-22
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.58 pmos
* Model Flag Parameters
+  lmin=1.0e-06 lmax=2.0e-06 wmin=1.26e-06 wmax=1.65e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.042356151e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-5.494114484e-08 wvth0=-7.312103119e-08 pvth0=1.061575563e-13
+  k1=6.801276767e-01 lk1=-4.526885438e-07 wk1=-4.047725987e-07 pk1=7.679221676e-13
+  k2=-6.765553831e-02 lk2=1.705207929e-07 wk2=1.532139738e-07 pk2=-2.908251739e-13
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=2.461148824e+00 ldsub=-1.923271921e-06 wdsub=-3.385511527e-06 pdsub=3.712505867e-12
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.845563200e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=7.864725187e-08 wvoff=1.022560197e-07 pvoff=-9.965743154e-14
+  nfactor={-3.169956695e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=4.671343506e-06 wnfactor=6.951655680e-06 pnfactor=-6.462577132e-12
+  eta0=4.530157834e-01 leta0=-2.427966211e-07 weta0=-8.405626160e-07 peta0=8.656704987e-13
+  etab=2.855797071e-01 letab=-1.167135412e-06 wetab=6.935233330e-07 petab=-6.731801677e-13
+  u0=-4.775050666e-03 lu0=1.424977049e-08 wu0=2.144391609e-08 pu0=-2.308835179e-14
+  ua=-3.080356731e-10 lua=-1.377827427e-16 wua=4.150390420e-16 pua=-1.002987985e-21
+  ub=-2.518996187e-18 lub=3.074052027e-24 wub=3.868659247e-24 pub=-3.221394664e-30
+  uc=-2.743025600e-10 luc=2.849467878e-16 wuc=2.472748056e-16 puc=-3.405316504e-22
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=-2.282030237e+04 lvsat=1.543102000e-01 wvsat=1.023537829e-01 pvsat=-2.071149267e-7
+  a0=5.769601848e-01 la0=1.246477269e-06 wa0=9.842115152e-07 pa0=-2.066454261e-12
+  ags=-2.760982896e-01 lags=8.871278327e-07 wags=5.572039899e-07 pags=-5.435564095e-13
+  a1=0.0
+  a2=1.451488817e+00 la2=-1.318300652e-06 wa2=-1.062755466e-06 pa2=2.150506941e-12
+  b0=0.0
+  b1=0.0
+  keta=2.427245306e-02 lketa=-4.431460332e-08 wketa=-4.353363830e-08 pketa=5.132764029e-14
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-1.318774538e+00 lpclm=1.390182686e-06 wpclm=2.201764067e-06 ppclm=-1.279565286e-12
+  pdiblc1=-6.720091506e-01 lpdiblc1=2.148996756e-06 wpdiblc1=1.764176040e-06 ppdiblc1=-3.569845501e-12
+  pdiblc2=-1.389733272e-03 lpdiblc2=1.862533399e-09 wpdiblc2=2.258783959e-09 ppdiblc2=-2.311910557e-15
+  pdiblcb=-0.025
+  drout=1.508213853e-01 ldrout=8.279811105e-07 wdrout=-5.110339822e-08 pdrout=1.034087484e-13
+  pscbe1=8.053522799e+08 lpscbe1=3.914368776e+01 wpscbe1=-8.731024316e+00 ppscbe1=-6.385400181e-5
+  pscbe2=-4.996524305e-08 lpscbe2=6.100806558e-14 wpscbe2=7.385042494e-14 ppscbe2=-7.617704962e-20
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=9.609784573e+00 lbeta0=3.144332065e-06 wbeta0=-4.651630812e-06 pbeta0=-1.608615537e-12
* Gidl Induced Drain Leakage Model Parameters
+  agidl=3.364291395e-10 lagidl=-4.551882637e-17 wagidl=-3.888532269e-16 pagidl=4.582647600e-23
+  bgidl=2.127758299e+09 lbgidl=-1.331988595e+02 wbgidl=-1.399854800e+03 pbgidl=1.653360147e-4
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-3.976145051e-01 lkt1=-5.538989282e-08 wkt1=-7.562095979e-08 pkt1=4.267367519e-14
+  kt2=-7.529804378e-02 lkt2=7.526578424e-08 wkt2=2.363851397e-08 pkt2=-8.364896712e-14
+  at=-3.998846012e+04 lat=2.792339989e-01 wat=1.700799295e-01 pat=-3.914153071e-7
+  ute=-2.978847688e+00 lute=6.463402854e-06 wute=4.859310826e-06 pute=-1.054356810e-11
+  ua1=-7.686917526e-09 lua1=1.956205821e-14 wua1=1.715866275e-14 pua1=-3.262491068e-20
+  ub1=7.193658236e-18 lub1=-1.609180890e-23 wub1=-1.423067165e-23 pub1=2.653730781e-29
+  uc1=1.066677844e-09 luc1=-1.722311998e-15 wuc1=-1.483621414e-15 puc1=2.386213233e-21
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=2.75e-6
+  sbref=2.74e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.59 pmos
* Model Flag Parameters
+  lmin=5.0e-07 lmax=1.0e-06 wmin=1.26e-06 wmax=1.65e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.172676988e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=7.844483850e-08 wvth0=9.947525267e-08 pvth0=-7.049819220e-14
+  k1=-2.857882199e-01 lk1=5.359456947e-07 wk1=9.956699866e-07 pk1=-6.654588273e-13
+  k2=2.621139570e-01 lk2=-1.670048810e-07 wk2=-3.401227816e-07 pk2=2.141148621e-13
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=-2.313045093e+00 ldsub=2.963211037e-06 wdsub=4.503636282e-06 pdsub=-4.362194699e-12
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.890451615e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=8.324167092e-08 wvoff=1.116021737e-07 pvoff=-1.092234071e-13
+  nfactor={-3.468393155e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=4.976799192e-06 wnfactor=6.537409379e-06 pnfactor=-6.038587758e-12
+  eta0=1.739327914e+00 leta0=-1.559362813e-06 weta0=-2.236807786e-06 peta0=2.294755355e-12
+  etab=-1.749571700e+00 letab=9.158827566e-07 wetab=7.399033223e-08 petab=-3.907575079e-14
+  u0=1.633163951e-02 lu0=-7.353349044e-09 wu0=-7.989998817e-09 pu0=7.037848797e-15
+  ua=6.136633849e-10 lua=-1.081160163e-15 wua=-1.438084814e-15 pua=8.937213440e-22
+  ub=5.452654961e-19 lub=-6.228109086e-26 wub=3.927395695e-25 pub=3.362786436e-31
+  uc=4.930131410e-11 luc=-4.626824947e-17 wuc=-1.870320964e-16 puc=1.039901499e-22
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=2.283994792e+05 lvsat=-1.028182708e-01 wvsat=-2.910174336e-01 pvsat=1.955083808e-7
+  a0=8.916872087e-01 la0=9.243478653e-07 wa0=4.042431213e-07 pa0=-1.472845010e-12
+  ags=-1.124291425e-01 lags=7.196091872e-07 wags=6.927089238e-08 pags=-4.414712552e-14
+  a1=0.0
+  a2=-7.453673034e-01 la2=9.302255249e-07 wa2=2.179330085e-06 pa2=-1.167832462e-12
+  b0=0.0
+  b1=0.0
+  keta=4.103387664e-02 lketa=-6.147025557e-08 wketa=-3.671165551e-08 pketa=4.434520447e-14
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-2.934450675e+00 lpclm=3.043859526e-06 wpclm=5.654501100e-06 ppclm=-4.813510695e-12
+  pdiblc1=-1.420483243e+00 lpdiblc1=2.915074959e-06 wpdiblc1=1.848005831e-06 ppdiblc1=-3.655646968e-12
+  pdiblc2=-3.442422075e-03 lpdiblc2=3.963501442e-09 wpdiblc2=5.313421019e-09 ppdiblc2=-5.438392681e-15
+  pdiblcb=-1.147944754e-01 lpdiblcb=9.190644142e-08 wpdiblcb=1.043491127e-07 ppdiblcb=-1.068034038e-13
+  drout=1.043677834e+00 ldrout=-8.587532164e-08 wdrout=-5.421607201e-08 pdrout=1.065946322e-13
+  pscbe1=9.275454577e+08 lpscbe1=-8.592347362e+01 wpscbe1=-1.931236510e+02 ppscbe1=1.248755394e-4
+  pscbe2=1.036515687e-08 lpscbe2=-7.413053514e-16 wpscbe2=-1.671890688e-15 ppscbe2=1.121550869e-21
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=1.447467444e+01 lbeta0=-1.834980015e-06 wbeta0=-9.856630844e-06 pbeta0=3.718806096e-12
* Gidl Induced Drain Leakage Model Parameters
+  agidl=4.623564241e-10 lagidl=-1.744079207e-16 wagidl=-5.531921542e-16 pagidl=2.140306549e-22
+  bgidl=2.185315369e+09 lbgidl=-1.921096712e+02 wbgidl=-1.471298779e+03 pbgidl=2.384603557e-4
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-5.656356877e-01 lkt1=1.165831480e-07 wkt1=1.841449543e-07 pkt1=-2.232019332e-13
+  kt2=9.600731246e-02 lkt2=-1.000686740e-07 wkt2=-2.001033945e-07 pkt2=1.453553511e-13
+  at=4.402668747e+05 lat=-2.123169414e-01 wat=-4.351648857e-01 pat=2.280648661e-7
+  ute=6.254914471e+00 lute=-2.987537392e-06 wute=-1.016930670e-05 pute=4.838522509e-12
+  ua1=2.251983117e-08 lua1=-1.135515322e-14 wua1=-3.238244483e-14 pua1=1.808140375e-20
+  ub1=-1.825492140e-17 lub1=9.955321324e-24 wub1=2.810252178e-23 pub1=-1.679156233e-29
+  uc1=-1.604440802e-09 luc1=1.011631359e-15 wuc1=2.415446482e-15 puc1=-1.604560739e-21
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.75e-6
+  sbref=1.74e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.60 pmos
* Model Flag Parameters
+  lmin=2.5e-07 lmax=5.0e-07 wmin=1.26e-06 wmax=1.65e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-8.662531095e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-8.197419055e-08 wvth0=-2.298021868e-07 pvth0=1.018851329e-13
+  k1=-9.867398537e-01 lk1=9.029078940e-07 wk1=1.837753177e-06 pk1=-1.106306219e-12
+  k2=6.162966578e-01 lk2=-3.524266085e-07 wk2=-7.663302415e-07 pk2=4.372429915e-13
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=7.270601689e+00 ldsub=-2.054019726e-06 wdsub=-9.447881432e-06 pdsub=2.941703855e-12
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={2.527106899e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-2.003783524e-07 wvoff=-4.088412753e-07 pvoff=1.632391474e-13
+  nfactor={9.788494842e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.963446812e-06 wnfactor=-1.074330866e-05 pnfactor=3.008213750e-12
+  eta0=-3.131258653e+00 leta0=9.904866669e-07 weta0=4.494966971e-06 peta0=-1.229463366e-12
+  etab=2.626320276e-03 letab=-1.427951106e-09 wetab=-4.876066798e-09 petab=2.212386428e-15
+  u0=8.556312568e-03 lu0=-3.282809883e-09 wu0=-1.428822100e-09 pu0=3.602941562e-15
+  ua=2.257937692e-09 lua=-1.941970648e-15 wua=-4.331098149e-15 pua=2.408271685e-21
+  ub=-3.256487204e-18 lub=1.928012482e-24 wub=5.613412887e-24 pub=-2.396848252e-30
+  uc=-4.357090571e-11 luc=2.352215043e-18 wuc=-2.325680932e-17 puc=1.825051162e-23
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=-1.421258041e+05 lvsat=9.115912551e-02 wvsat=2.965229295e-01 pvsat=-1.120807501e-7
+  a0=4.160673783e+00 la0=-7.870319862e-07 wa0=-4.107598996e-06 pa0=8.891945752e-13
+  ags=2.242054900e+00 lags=-5.130102986e-07 wags=-1.608404891e-06 pags=8.341497006e-13
+  a1=0.0
+  a2=1.912301648e+00 la2=-4.611173247e-07 wa2=-8.865641790e-07 pa2=4.372245029e-13
+  b0=0.0
+  b1=0.0
+  keta=5.835383152e-02 lketa=-7.053759835e-08 wketa=-1.252348466e-07 pketa=9.068886547e-14
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=4.891986972e+00 lpclm=-1.053437111e-06 wpclm=-6.867132917e-06 ppclm=1.741815146e-12
+  pdiblc1=7.997081835e+00 lpdiblc1=-2.015208711e-06 wpdiblc1=-1.045312517e-05 ppdiblc1=2.784241134e-12
+  pdiblc2=-4.552373478e-03 lpdiblc2=4.544583201e-09 wpdiblc2=-6.730057013e-09 ppdiblc2=8.666089381e-16
+  pdiblcb=4.012918651e-01 lpdiblcb=-1.782750795e-07 wpdiblcb=-2.548741237e-07 ppdiblcb=8.125714492e-14
+  drout=4.130032884e-01 ldrout=2.442954163e-07 wdrout=1.422497597e-06 pdrout=-6.664945078e-13
+  pscbe1=7.232956861e+08 lpscbe1=2.100536683e+01 wpscbe1=9.525023272e+01 ppscbe1=-2.609395618e-5
+  pscbe2=7.968550522e-09 lpscbe2=5.133660054e-16 wpscbe2=1.922933002e-15 ppscbe2=-7.604112296e-22
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=1.321894906e+01 lbeta0=-1.177582660e-06 wbeta0=-5.823772064e-06 pbeta0=1.607523867e-12
* Gidl Induced Drain Leakage Model Parameters
+  agidl=5.639846648e-10 lagidl=-2.276123373e-16 wagidl=-7.809294348e-16 pagidl=3.332556760e-22
+  bgidl=3.620354977e+09 lbgidl=-9.433816067e+02 wbgidl=-3.606166116e+03 pbgidl=1.356106104e-3
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-8.529053273e-01 lkt1=2.669745497e-07 wkt1=3.627330786e-07 pkt1=-3.166963880e-13
+  kt2=-1.604411764e-01 lkt2=3.418723889e-08 wkt2=1.861986471e-07 pkt2=-5.688149375e-14
+  at=2.784336040e+05 lat=-1.275939875e-01 wat=-3.522565608e-01 pat=1.846606999e-7
+  ute=-1.769354095e+00 lute=1.213327688e-06 wute=2.853672352e-06 pute=-1.979267484e-12
+  ua1=-1.156287008e-09 lua1=1.039768171e-15 wua1=7.712026401e-15 pua1=-2.908853827e-21
+  ub1=3.135134957e-18 lub1=-1.242800979e-24 wub1=-9.993987188e-24 pub1=3.152722044e-30
+  uc1=4.459443786e-10 luc1=-6.178629081e-17 wuc1=-9.205009749e-16 puc1=1.418744736e-22
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.25e-6
+  sbref=1.24e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.61 pmos
* Model Flag Parameters
+  lmin=1.8e-07 lmax=2.5e-07 wmin=1.26e-06 wmax=1.65e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-2.026e-8
+  vth0={-1.382375472e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=6.287476286e-08 wvth0=4.957361815e-07 pvth0=-1.025658402e-13
+  k1=7.758209005e+00 lk1=-1.581556506e-06 wk1=-1.108739813e-05 pk1=2.579948845e-12
+  k2=-2.749211087e+00 lk2=6.034164447e-07 wk2=4.220435434e-06 pk2=-9.843363506e-13
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=-4.809873132e+00 ldsub=1.327936996e-06 wdsub=8.763481164e-06 pdsub=-2.166226439e-12
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-9.922236141e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=1.488459107e-07 wvoff=1.023738457e-06 pvoff=-2.428081665e-13
+  nfactor={-2.565182849e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.503510157e-06 wnfactor=8.697061387e-06 pnfactor=-2.452634021e-12
+  eta0=-2.788042768e+00 leta0=9.523369849e-07 weta0=5.347379382e-06 peta0=-1.553520658e-12
+  etab=-2.698658865e-01 letab=7.764773381e-08 wetab=4.392051193e-07 petab=-1.266645740e-13
+  u0=-3.047078025e-02 lu0=7.851305703e-09 wu0=5.582881654e-08 pu0=-1.280761516e-14
+  ua=-1.398218141e-08 lua=2.655410080e-15 wua=1.938378664e-14 pua=-4.331696113e-21
+  ub=9.897371716e-18 lub=-1.773615475e-24 wub=-1.310842399e-23 pub=2.893249264e-30
+  uc=-2.000594219e-10 luc=4.796145522e-17 wuc=3.127717214e-16 puc=-7.823817898e-23
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=-4.540862225e+04 lvsat=6.872663345e-02 wvsat=2.726518160e-01 pvsat=-1.121118328e-7
+  a0=1.942801166e+00 la0=-1.916117778e-07 wa0=-1.932569842e-06 pa0=3.125709280e-13
+  ags=-2.416906385e+00 lags=8.086261708e-07 wags=5.981721667e-06 pags=-1.319089231e-12
+  a1=0.0
+  a2=-1.267091402e+00 la2=4.339002684e-07 wa2=3.148299288e-06 pa2=-7.078093586e-13
+  b0=0.0
+  b1=0.0
+  keta=-3.420721220e-01 lketa=4.141004915e-08 wketa=4.388449925e-07 pketa=-6.755105369e-14
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=1.877288253e+00 lpclm=-2.430807753e-07 wpclm=-1.863887852e-06 ppclm=3.965308625e-13
+  pdiblc1=3.849592278e-01 lpdiblc1=7.101453488e-08 wpdiblc1=1.249183163e-07 ppdiblc1=-1.158440223e-13
+  pdiblc2=-1.332163730e-03 lpdiblc2=3.891505873e-09 wpdiblc2=1.828913468e-08 ppdiblc2=-6.348104569e-15
+  pdiblcb=-3.358418803e-01 lpdiblcb=2.479674291e-08 wpdiblcb=1.814391295e-07 ppdiblcb=-4.045023240e-14
+  drout=2.732866059e+00 ldrout=-4.144875018e-07 wdrout=-3.341583297e-06 pdrout=6.761418561e-13
+  pscbe1=8.003824119e+08 lpscbe1=-8.432899007e-02 wpscbe1=-6.238169524e-01 ppscbe1=1.375635203e-7
+  pscbe2=1.061108282e-08 lpscbe2=-2.224354073e-16 wpscbe2=-2.106137197e-15 ppscbe2=3.628526517e-22
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=3.676687383e+00 lbeta0=1.521445287e-06 wbeta0=8.596325948e-06 pbeta0=-2.481891097e-12
* Gidl Induced Drain Leakage Model Parameters
+  agidl=-1.113003672e-09 lagidl=2.454395984e-16 wagidl=1.815611777e-15 pagidl=-4.003787446e-22
+  bgidl=-2.439282110e+09 lbgidl=7.584304682e+02 wbgidl=5.610404566e+03 pbgidl=-1.237206387e-3
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-1.106e-8
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-1.842988752e+00 lkt1=5.712067691e-07 wkt1=2.412208820e-06 pkt1=-9.317936086e-13
+  kt2=-3.702971357e-02 lkt2=4.585691050e-10 wkt2=-1.918748768e-08 pkt2=-7.480509411e-16
+  at=-6.171055829e+05 lat=1.246477493e-01 wat=1.022768359e+00 pat=-2.033343832e-7
+  ute=8.533360344e+00 lute=-1.704405348e-06 wute=-1.395285723e-05 pute=2.780348721e-12
+  ua1=4.050390218e-09 lua1=-4.082513220e-16 wua1=-5.215193162e-15 pua1=6.659689506e-22
+  ub1=-1.085415616e-18 lub1=-9.389003328e-26 wub1=1.005296763e-24 pub1=1.531601824e-31
+  uc1=7.340109022e-10 luc1=-1.493155606e-16 wuc1=-1.240210259e-15 puc1=2.435742931e-22
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.04e-6
+  sbref=1.04e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.62 pmos
* Model Flag Parameters
+  lmin=1.5e-07 lmax=1.8e-07 wmin=1.26e-06 wmax=1.65e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-2.026e-8
+  vth0={-9.551685118e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-3.133291599e-08 wvth0=-1.457408340e-07 pvth0=3.889267129e-14
+  k1=-2.797625280e+00 lk1=7.462160702e-07 wk1=4.812320534e-06 pk1=-9.262571139e-13
+  k2=1.481215542e+00 lk2=-3.294772357e-07 wk2=-2.097845075e-06 pk2=4.089708673e-13
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=8.289211859e+00 ldsub=-1.560673226e-06 wdsub=-9.844565345e-06 pdsub=1.937219977e-12
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.044514321e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-2.487361084e-08 wvoff=-2.173420946e-07 pvoff=3.087491667e-14
+  nfactor={1.023161802e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.318440371e-06 wnfactor=-9.846277711e-06 pnfactor=1.636543117e-12
+  eta0=1.050284235e+01 leta0=-1.978569000e-06 weta0=-1.283447695e-05 peta0=2.455942300e-12
+  etab=1.272032523e+00 letab=-2.623717035e-07 wetab=-1.612033876e-06 petab=3.256746492e-13
+  u0=-6.830732044e-03 lu0=2.638202272e-09 wu0=1.259968293e-08 pu0=-3.274726611e-15
+  ua=-8.889088190e-09 lua=1.532281164e-15 wua=8.365654912e-15 pua=-1.901977705e-21
+  ub=9.362545582e-18 lub=-1.655675616e-24 wub=-9.307836828e-24 pub=2.055143783e-30
+  uc=1.105959666e-10 luc=-2.054427105e-17 wuc=-1.576582051e-16 puc=2.550102842e-23
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=1.368694826e+06 lvsat=-2.431114590e-01 wvsat=-1.604181486e+00 pvsat=3.017674470e-7
+  a0=3.853735885e+00 la0=-6.130111018e-07 wa0=-3.965685154e-06 pa0=7.609135164e-13
+  ags=1.249999161e+00 lags=1.597980122e-13 wags=1.041112732e-12 pags=-1.983527973e-19
+  a1=0.0
+  a2=-2.503195986e-01 la2=2.096817504e-07 wa2=1.118835870e-06 pa2=-2.602720857e-13
+  b0=-5.597672795e-23 lb0=1.234398805e-29 wb0=6.948234505e-29 pb0=-1.532224673e-35
+  b1=0.0
+  keta=-1.623342194e+00 lketa=3.239557253e-07 wketa=1.956014036e-06 pketa=-4.021171711e-13
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=2.583920779e+00 lpclm=-3.989073799e-07 wpclm=-2.311111228e-06 ppclm=4.951525612e-13
+  pdiblc1=8.555396193e+00 lpdiblc1=-1.730730225e-06 wpdiblc1=-1.014240886e-05 ppdiblc1=2.148306968e-12
+  pdiblc2=1.722478240e-01 lpdiblc2=-3.438635302e-08 wpdiblc2=-2.040531551e-07 ppdiblc2=4.268281719e-14
+  pdiblcb=-4.197690012e+00 lpdiblcb=8.764114929e-07 wpdiblcb=4.931188876e-06 ppdiblcb=-1.087865047e-12
+  drout=-7.529724582e+00 ldrout=1.848618986e-06 wdrout=1.013012377e-05 pdrout=-2.294638986e-12
+  pscbe1=8.099225170e+08 lpscbe1=-2.188112971e+00 wpscbe1=-1.231654253e+01 ppscbe1=2.716043364e-6
+  pscbe2=5.091023655e-08 lpscbe2=-9.109204788e-15 wpscbe2=-5.173496086e-14 ppscbe2=1.130700085e-20
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=2.894087620e+01 lbeta0=-4.049813630e-06 wbeta0=-2.545415184e-05 pbeta0=5.026920264e-12
* Gidl Induced Drain Leakage Model Parameters
+  agidl=5.526644047e-15 lagidl=-1.190063457e-21 wagidl=-6.860068509e-21 pagidl=1.477192448e-27
+  bgidl=9.999992434e+08 lbgidl=1.441405916e-04 wbgidl=9.391018295e-04 pbgidl=-1.789176798e-10
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-1.106e-8
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=1.007151470e+01 lkt1=-2.056179532e-06 wkt1=-1.338713676e-05 pkt1=2.552278080e-12
+  kt2=8.057340185e-02 lkt2=-2.547526991e-08 wkt2=-1.659759430e-07 pkt2=3.162173923e-14
+  at=-5.670711856e+05 lat=1.136141640e-01 wat=7.402166511e-01 pat=-1.410260805e-7
+  ute=7.684211440e+00 lute=-1.517151031e-06 wute=-9.884511390e-06 pute=1.883197095e-12
+  ua1=1.217118698e-08 lua1=-2.199049425e-15 wua1=-1.457329912e-14 pua1=2.729618477e-21
+  ub1=-1.020798987e-17 lub1=1.917820041e-24 wub1=1.249494170e-23 pub1=-2.380536318e-30
+  uc1=7.510020288e-10 luc1=-1.530624438e-16 wuc1=-9.972292717e-16 puc1=1.899921258e-22
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.04e-6
+  sbref=1.04e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.63 pmos
* Model Flag Parameters
+  lmin=2.0e-05 lmax=0.0001 wmin=1.12e-06 wmax=1.26e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-5.165091571e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-1.144725702e-05 wvth0=-6.820627614e-07 pvth0=1.365729734e-11
+  k1=1.028787392e+00 lk1=-1.163906551e-05 wk1=-6.619767639e-07 pk1=1.325510497e-11
+  k2=-1.254950285e-01 lk2=2.933047982e-06 wk2=1.695689575e-07 pk2=-3.395367411e-12
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.051579485e-04 lcit=-1.905397086e-09 wcit=-1.181168971e-10 pcit=2.365116052e-15
+  voff={2.752828955e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-9.757717908e-06 wvoff=-5.621200654e-07 pvoff=1.125562237e-11
+  nfactor={8.891969522e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.417117898e-04 wnfactor=-7.708367640e-06 pnfactor=1.543486536e-10
+  eta0=0.08
+  etab=-0.07
+  u0=-5.727520750e-03 lu0=2.952792555e-07 wu0=1.702116371e-08 pu0=-3.408236120e-13
+  ua=4.397848549e-09 lua=-1.026118015e-13 wua=-5.672266487e-15 pua=1.135787414e-19
+  ub=-7.400829821e-18 lub=1.679192597e-22 wub=9.187451686e-24 pub=-1.839651226e-28
+  uc=-1.533801106e-10 luc=1.633983339e-15 wuc=4.320910932e-17 puc=-8.651984647e-22
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=9.486601895e+05 lvsat=-1.578554579e+01 wvsat=-9.785531365e-01 pvsat=1.959407830e-5
+  a0=3.750159209e+00 la0=-5.001076776e-05 wa0=-2.459400876e-06 pa0=4.924586264e-11
+  ags=3.304807341e+00 lags=-6.135880002e-05 wags=-3.549785082e-06 pags=7.107919258e-11
+  a1=0.0
+  a2=-8.719667255e-01 la2=3.347865917e-05 wa2=2.075365481e-06 pa2=-4.155612222e-11
+  b0=8.839097972e-07 lb0=-1.769898550e-11 wb0=-1.097172482e-12 pb0=2.196925513e-17
+  b1=-3.330065962e-08 lb1=6.667964240e-13 wb1=4.133517637e-14 pb1=-8.276757308e-19
+  keta=-5.755552203e-01 lketa=1.148719348e-05 wketa=6.665247931e-07 pketa=-1.334617252e-11
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=4.839361768e-01 lpclm=-6.867610759e-06 wpclm=-5.511458380e-07 ppclm=1.103587971e-11
+  pdiblc1=0.39
+  pdiblc2=-9.459509058e-03 lpdiblc2=1.958061391e-07 wpdiblc2=1.208801813e-08 ppdiblc2=-2.420446728e-13
+  pdiblcb=2.234758398e+00 lpdiblcb=-4.785376849e-05 wpdiblcb=-2.728125027e-06 ppdiblcb=5.462666604e-11
+  drout=0.56
+  pscbe1=6.920360458e+08 lpscbe1=2.160842249e+03 wpscbe1=1.189111173e+02 ppscbe1=-2.381019135e-3
+  pscbe2=3.460011475e-09 lpscbe2=3.935525391e-14 wpscbe2=8.546715189e-15 ppscbe2=-1.711353225e-19
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.083509839e-09 lalpha0=-1.969332892e-14 walpha0=-1.220803224e-15 palpha0=2.444477778e-20
+  alpha1=1.083509839e-09 lalpha1=-1.969332892e-14 walpha1=-1.220803224e-15 palpha1=2.444477778e-20
+  beta0=-2.633682676e+02 lbeta0=5.399279233e-03 wbeta0=3.296168706e-04 pbeta0=-6.600090000e-9
* Gidl Induced Drain Leakage Model Parameters
+  agidl=-3.705149840e-09 lagidl=3.353388467e-13 wagidl=6.153528238e-16 pagidl=-1.232152957e-20
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=-9.659333470e-02 legidl=1.966395734e-5
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-6.292853180e-01 lkt1=3.774710205e-06 wkt1=2.110768775e-07 pkt1=-4.226502078e-12
+  kt2=1.680981011e-01 lkt2=-4.414316601e-06 wkt2=-2.513023437e-07 pkt2=5.031957506e-12
+  at=-6.981936344e+05 lat=1.398029420e+01 wat=8.666482089e-01 pat=-1.735334774e-5
+  ute=-2.805521135e+00 lute=5.352797526e-05 wute=3.011843635e-06 pute=-6.030771126e-11
+  ua1=6.689964509e-09 lua1=-9.745928168e-14 wua1=-4.991864384e-15 pua1=9.995469633e-20
+  ub1=-6.366792424e-18 lub1=1.131509801e-22 wub1=5.516809771e-24 pub1=-1.104659508e-28
+  uc1=5.016217549e-09 luc1=-1.006177639e-13 wuc1=-5.562821844e-15 puc1=1.113872745e-19
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.64 pmos
* Model Flag Parameters
+  lmin=8.0e-06 lmax=2.0e-05 wmin=1.12e-06 wmax=1.26e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.0881997+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+  k1=0.44751769
+  k2=0.02098511
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-0.21202992+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.8147029+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+  eta0=0.08
+  etab=-0.07
+  u0=0.0090191
+  ua=-7.2671504e-10
+  ub=9.8527111e-19
+  uc=-7.1776909e-11
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=160310.0
+  a0=1.252558
+  ags=0.240471
+  a1=0.0
+  a2=0.8
+  b0=0.0
+  b1=0.0
+  keta=-0.0018702
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=0.14095898
+  pdiblc1=0.39
+  pdiblc2=0.00031929802
+  pdiblcb=-0.15511953
+  drout=0.56
+  pscbe1=799951250.0
+  pscbe2=5.4254628e-9
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=6.2785893
* Gidl Induced Drain Leakage Model Parameters
+  agidl=1.304209773e-8
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.88544965
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-0.4407715
+  kt2=-0.052358472
+  at=0.0
+  ute=-0.13226612
+  ua1=1.8227243e-9
+  ub1=-7.1588888e-19
+  uc1=-8.7612717e-12
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.65 pmos
* Model Flag Parameters
+  lmin=4.0e-06 lmax=8.0e-06 wmin=1.12e-06 wmax=1.26e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.090414346e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=1.776925644e-8
+  k1=4.556728822e-01 lk1=-6.543334786e-8
+  k2=1.885398624e-02 lk2=1.709911408e-8
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.057269452e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-5.057204472e-8
+  nfactor={2.150233085e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-2.692133146e-6
+  eta0=0.08
+  etab=-0.07
+  u0=8.535573484e-03 lu0=3.879584672e-9
+  ua=-8.237874492e-10 lua=7.788624164e-16 wua=1.654361225e-30
+  ub=1.048518672e-18 lub=-5.074680762e-25
+  uc=-7.083802061e-11 luc=-7.533189791e-18
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=2.678104074e+05 lvsat=-8.625316685e-1
+  a0=1.347035279e+00 la0=-7.580403376e-7
+  ags=2.084960866e-01 lags=2.565513575e-7
+  a1=0.0
+  a2=0.8
+  b0=0.0
+  b1=0.0
+  keta=-8.364571240e-04 lketa=-8.294256640e-9
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=2.407132755e-01 lpclm=-8.003805848e-7
+  pdiblc1=0.39
+  pdiblc2=-1.397670217e-03 lpdiblc2=1.377612899e-08 wpdiblc2=8.673617380e-25 ppdiblc2=-1.387778781e-29
+  pdiblcb=-2.494013897e-01 lpdiblcb=7.564723865e-7
+  drout=0.56
+  pscbe1=1.227212561e+09 lpscbe1=-3.428139670e+3
+  pscbe2=-1.711599940e-08 lpscbe2=1.808618728e-13
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=3.429576331e+00 lbeta0=2.285911254e-5
* Gidl Induced Drain Leakage Model Parameters
+  agidl=2.613220901e-08 lagidl=-1.050287696e-13
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=1.675517744e+00 legidl=-6.339127153e-6
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.061103840e-01 lkt1=-2.781041573e-7
+  kt2=-4.839276194e-02 lkt2=-3.181895402e-8
+  at=-9.120917488e+04 lat=7.318186388e-1
+  ute=-1.647219648e-01 lute=2.604101198e-7
+  ua1=5.703275549e-10 lua1=1.004863033e-14
+  ub1=8.239234094e-19 lub1=-1.235471470e-23 pub1=1.232595164e-44
+  uc1=-1.164852119e-11 luc1=2.316590399e-17
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.66 pmos
* Model Flag Parameters
+  lmin=2.0e-06 lmax=4.0e-06 wmin=1.12e-06 wmax=1.26e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.085843201e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-6.228379991e-10
+  k1=4.428072554e-01 lk1=-1.366824095e-8
+  k2=2.193345702e-02 lk2=4.708801823e-9
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=8.622137339e-01 ldsub=-1.215963003e-6
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.337857314e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=6.232304277e-8
+  nfactor={7.881674337e-01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=2.788165241e-6
+  eta0=1.604349200e-01 leta0=-3.236315093e-7
+  etab=-1.403185835e-01 letab=2.829282271e-7
+  u0=8.638994592e-03 lu0=3.463467775e-9
+  ua=-8.215637429e-10 lua=7.699152898e-16 wua=-1.654361225e-30
+  ub=1.011504174e-18 lub=-3.585395030e-25
+  uc=-7.560382119e-11 luc=1.164210416e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=53438.0
+  a0=1.154071298e+00 la0=1.835409954e-8
+  ags=1.482758150e-01 lags=4.988488244e-7
+  a1=0.0
+  a2=0.8
+  b0=0.0
+  b1=0.0
+  keta=6.578345336e-03 lketa=-3.812786263e-08 wketa=6.938893904e-24
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-5.559724103e-01 lpclm=2.405100206e-06 wpclm=-1.110223025e-22
+  pdiblc1=0.39
+  pdiblc2=3.641230659e-03 lpdiblc2=-6.497989463e-9
+  pdiblcb=-9.820554637e-02 lpdiblcb=1.481328872e-7
+  drout=0.56
+  pscbe1=-4.676991234e+07 lpscbe1=1.697754289e+3
+  pscbe2=4.653609693e-08 lpscbe2=-7.524360986e-14
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=1.147359093e+01 lbeta0=-9.506141085e-6
* Gidl Induced Drain Leakage Model Parameters
+  agidl=3.821637237e-11 lagidl=-3.906838872e-17
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.816142056e-01 lkt1=2.568697892e-8
+  kt2=-6.028632264e-02 lkt2=1.603502535e-8
+  at=1.022950518e+05 lat=-4.674948746e-2
+  ute=-1.327375183e-01 lute=1.317200597e-7
+  ua1=3.323674104e-09 lua1=-1.029514575e-15
+  ub1=-2.842323112e-18 lub1=2.396501504e-24
+  uc1=1.818504214e-11 luc1=-9.687003470e-17 puc1=5.169878828e-38
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.67 pmos
* Model Flag Parameters
+  lmin=1.0e-06 lmax=2.0e-06 wmin=1.12e-06 wmax=1.26e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.101264296e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=3.058205737e-8
+  k1=3.540326720e-01 lk1=1.659689040e-7
+  k2=5.577749960e-02 lk2=-6.377529522e-08 pk2=5.551115123e-29
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=-2.663045674e-01 ldsub=1.067616350e-6
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.021762939e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-1.639286090e-9
+  nfactor={2.430472285e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-5.350714714e-7
+  eta0=-2.241626400e-01 leta0=4.546093453e-07 weta0=8.500145032e-23 peta0=-2.116362641e-28
+  etab=8.442995791e-01 letab=-1.709466317e-06 wetab=3.608224830e-22 petab=7.546047120e-28
+  u0=1.250070846e-02 lu0=-4.350787479e-9
+  ua=2.633023699e-11 lua=-9.458151364e-16
+  ub=5.976931819e-19 lub=4.788153150e-25
+  uc=-7.509174596e-11 luc=1.060590969e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=5.963848416e+04 lvsat=-1.254680371e-2
+  a0=1.369865781e+00 la0=-4.183103528e-7
+  ags=1.727992847e-01 lags=4.492250930e-7
+  a1=0.0
+  a2=5.953062352e-01 la2=4.142019269e-7
+  b0=0.0
+  b1=0.0
+  keta=-1.079934288e-02 lketa=-2.963762975e-9
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=4.550220723e-01 lpclm=3.593326501e-7
+  pdiblc1=7.492555200e-01 lpdiblc1=-7.269607298e-7
+  pdiblc2=0.00043
+  pdiblcb=-0.025
+  drout=1.096512000e-01 ldrout=9.112898038e-7
+  pscbe1=7.983183467e+08 lpscbe1=-1.229870506e+1
+  pscbe2=9.530520115e-09 lpscbe2=-3.620850560e-16
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=5.862313582e+00 lbeta0=1.848390856e-6
* Gidl Induced Drain Leakage Model Parameters
+  agidl=2.315918186e-11 lagidl=-8.599862589e-18
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.585366557e-01 lkt1=-2.101090483e-8
+  kt2=-5.625426130e-02 lkt2=7.876068592e-9
+  at=9.703221664e+04 lat=-3.610003518e-2
+  ute=9.359355551e-01 lute=-2.030761278e-06 wute=4.440892099e-22 pute=1.110223025e-27
+  ua1=6.136533540e-09 lua1=-6.721391901e-15
+  ub1=-4.270929418e-18 lub1=5.287314936e-24
+  uc1=-1.285649500e-10 luc1=2.000815094e-16 wuc1=1.033975766e-31 puc1=-1.033975766e-37
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=2.75e-6
+  sbref=2.74e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.68 pmos
* Model Flag Parameters
+  lmin=5.0e-07 lmax=1.0e-06 wmin=1.12e-06 wmax=1.26e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.092537218e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=2.164971849e-8
+  k1=5.163486096e-01 lk1=-1.647044061e-10
+  k2=-1.189752607e-02 lk2=5.491447057e-9
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=1.315197776e+00 ldsub=-5.510829280e-7
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-1.991356383e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-4.751457949e-9
+  nfactor={1.798308567e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.119607376e-7
+  eta0=-6.270080000e-02 leta0=2.893499228e-7
+  etab=-1.689963224e+00 letab=8.844023472e-7
+  u0=9.894695136e-03 lu0=-1.683480718e-9
+  ua=-5.448939775e-10 lua=-3.611557284e-16
+  ub=8.616663893e-19 lub=2.086334578e-25
+  uc=-1.013764555e-10 luc=3.750883558e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=-6.051498240e+03 lvsat=5.468820708e-2
+  a0=1.217355653e+00 la0=-2.622131867e-7
+  ags=-5.662276614e-02 lags=6.840431505e-7
+  a1=0.0
+  a2=1.010355926e+00 la2=-1.060973294e-8
+  b0=0.0
+  b1=0.0
+  keta=1.145804192e-02 lketa=-2.574464147e-8
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=1.620957890e+00 lpclm=-8.340259780e-7
+  pdiblc1=6.831681950e-02 lpdiblc1=-3.000635109e-8
+  pdiblc2=8.382037816e-04 lpdiblc2=-4.178047345e-10
+  pdiblcb=-3.072820088e-02 lpdiblcb=5.862928163e-09 wpdiblcb=5.551115123e-23
+  drout=1.0
+  pscbe1=7.719601783e+08 lpscbe1=1.467940745e+1
+  pscbe2=9.018239607e-09 lpscbe2=1.622442887e-16
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=6.533924275e+00 lbeta0=1.160983879e-6
* Gidl Induced Drain Leakage Model Parameters
+  agidl=1.669088570e-11 lagidl=-1.979432105e-18
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.172838726e-01 lkt1=-6.323395343e-8
+  kt2=-6.520102427e-02 lkt2=1.703325943e-8
+  at=8.968707775e+04 lat=-2.858213862e-2
+  ute=-1.937735245e+00 lute=9.104982595e-7
+  ua1=-3.568282344e-09 lua1=3.211681253e-15 pua1=1.654361225e-36
+  ub1=4.385178260e-18 lub1=-3.572384395e-24 pub1=1.540743956e-45
+  uc1=3.415037467e-10 luc1=-2.810432031e-16 wuc1=2.067951531e-31 puc1=-2.067951531e-37
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.75e-6
+  sbref=1.74e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.69 pmos
* Model Flag Parameters
+  lmin=2.5e-07 lmax=5.0e-07 wmin=1.12e-06 wmax=1.26e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.051387542e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=1.070397737e-10
+  k1=4.938004126e-01 lk1=1.163972768e-8
+  k2=-1.078294214e-03 lk2=-1.726372043e-10
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=-3.408496543e-01 ldsub=3.158910227e-07 pdsub=-2.220446049e-28
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-7.666214318e-02+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-6.886878211e-8
+  nfactor={1.133414681e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=4.600459844e-7
+  eta0=0.49
+  etab=-1.301962000e-03 letab=3.544031462e-10
+  u0=7.405217482e-03 lu0=-3.801893760e-10
+  ua=-1.231304109e-09 lua=-1.806296181e-18
+  ub=1.265819661e-18 lub=-2.948863286e-27
+  uc=-6.230717731e-11 luc=1.705528707e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=9.676053951e+04 lvsat=8.640490753e-4
+  a0=8.514885312e-01 la0=-7.067443105e-8
+  ags=9.462833920e-01 lags=1.590017186e-7
+  a1=0.0
+  a2=1.198063207e+00 la2=-1.088782482e-7
+  b0=0.0
+  b1=0.0
+  keta=-4.253851648e-02 lketa=2.523636788e-9
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-6.403483396e-01 lpclm=3.498130593e-07 wpclm=-1.110223025e-22 ppclm=1.387778781e-28
+  pdiblc1=-4.242191933e-01 lpdiblc1=2.278461023e-07 wpdiblc1=-3.053113318e-22 ppdiblc1=-9.020562075e-29
+  pdiblc2=-9.974276988e-03 lpdiblc2=5.242745198e-09 wpdiblc2=-4.336808690e-24 ppdiblc2=1.355252716e-30
+  pdiblcb=1.959588488e-01 lpdiblcb=-1.128122761e-07 wpdiblcb=-1.110223025e-22 ppdiblcb=6.938893904e-29
+  drout=1.559003196e+00 ldrout=-2.926493531e-7
+  pscbe1=8.000316736e+08 lpscbe1=-1.658177145e-2
+  pscbe2=9.517713802e-09 lpscbe2=-9.924044155e-17
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=8.527171537e+00 lbeta0=1.174790728e-7
* Gidl Induced Drain Leakage Model Parameters
+  agidl=-6.515176521e-11 lagidl=4.086683250e-17 wagidl=5.169878828e-32 pagidl=1.292469707e-38
+  bgidl=7.151366880e+08 lbgidl=1.491316411e+2
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-5.606784192e-01 lkt1=1.183595963e-8
+  kt2=-1.043485456e-02 lkt2=-1.163792574e-8
+  at=-5.353157337e+03 lat=2.117332525e-2
+  ute=5.296362567e-01 lute=-3.812200691e-7
+  ua1=5.056715784e-09 lua1=-1.303677767e-15
+  ub1=-4.916272944e-18 lub1=1.297111340e-24
+  uc1=-2.956344010e-10 luc1=5.251136002e-17
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.25e-6
+  sbref=1.24e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.70 pmos
* Model Flag Parameters
+  lmin=1.8e-07 lmax=2.5e-07 wmin=1.12e-06 wmax=1.26e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-7.194201058e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-9.069269328e-08 wvth0=-3.336785280e-07 pvth0=9.126775097e-14
+  k1=-4.134836916e+00 lk1=1.277664610e-06 wk1=3.838778706e-06 pk1=-1.049982752e-12
+  k2=2.031590043e+00 lk2=-5.561480807e-07 wk2=-1.776285437e-06 pk2=4.858495928e-13
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=1.681819276e+01 ldsub=-4.377450258e-06 wdsub=-1.822025683e-05 pdsub=4.983604649e-12
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-7.968354126e-02+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-6.804236930e-08 wvoff=-1.243757331e-07 pvoff=3.401925051e-14
+  nfactor={1.088584881e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-2.207439799e-06 wnfactor=-8.154922672e-06 pnfactor=2.230534449e-12
+  eta0=7.035815116e+00 leta0=-1.790411351e-06 weta0=-6.945255682e-06 peta0=1.899666334e-12
+  etab=6.871388140e-01 letab=-1.879479179e-07 wetab=-7.567336189e-07 petab=2.069817795e-13
+  u0=-5.930098458e-03 lu0=3.267286240e-09 wu0=2.455464036e-08 pu0=-6.716185230e-15
+  ua=-5.894820924e-09 lua=1.273758823e-15 wua=9.070369742e-15 pua=-2.480927532e-21
+  ub=6.179859204e-18 lub=-1.347036959e-24 wub=-8.310432082e-24 pub=2.273069383e-30
+  uc=1.985696149e-10 luc=-5.429973314e-17 wuc=-1.869987699e-16 puc=5.114790355e-23
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=2.146865009e+06 lvsat=-5.598805255e-01 wvsat=-2.455668433e+00 pvsat=6.716744298e-7
+  a0=6.272934813e+00 la0=-1.553548418e-06 wa0=-7.287613996e-06 pa0=1.993308180e-12
+  ags=2.334702171e+00 lags=-2.207585859e-7
+  a1=0.0
+  a2=-6.312122885e-01 la2=3.914651851e-07 wa2=2.314096929e-06 pa2=-6.329517919e-13
+  b0=0.0
+  b1=0.0
+  keta=-6.907644317e-02 lketa=9.782290495e-09 wketa=9.569766188e-08 pketa=-2.617522448e-14
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-4.822239554e-01 lpclm=3.065628778e-07 wpclm=1.090064501e-06 ppclm=-2.981544424e-13
+  pdiblc1=7.971008132e-01 lpdiblc1=-1.062093458e-07 wpdiblc1=-3.940106377e-07 ppdiblc1=1.077697896e-13
+  pdiblc2=6.066557585e-02 lpdiblc2=-1.407866735e-08 wpdiblc2=-5.906964723e-08 ppdiblc2=1.615672991e-14
+  pdiblcb=1.897581226e+00 lpdiblcb=-5.782400286e-07 wpdiblcb=-2.593412599e-06 ppdiblcb=7.093502139e-13
+  drout=-3.167474748e+00 ldrout=1.000136894e-06 wdrout=4.025238972e-06 pdrout=-1.100983364e-12
+  pscbe1=7.998868799e+08 lpscbe1=2.302219403e-2
+  pscbe2=-4.994530916e-08 lpscbe2=1.616508560e-14 wpscbe2=7.308383597e-14 ppscbe2=-1.998989081e-20
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=2.927294729e+01 lbeta0=-5.556905511e-06 wbeta0=-2.333304593e-05 pbeta0=6.382054724e-12
* Gidl Induced Drain Leakage Model Parameters
+  agidl=3.292360240e-10 lagidl=-6.700611560e-17
+  bgidl=2.017368972e+09 lbgidl=-2.070549331e+2
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=5.125995571e+00 lkt1=-1.543583110e-06 wkt1=-6.297309268e-06 pkt1=1.722440031e-12
+  kt2=1.792894955e-01 lkt2=-6.353132997e-08 wkt2=-2.877459213e-07 pkt2=7.870426440e-14
+  at=6.977915000e+05 lat=-1.711508014e-01 wat=-6.222761045e-01 pat=1.702049601e-7
+  ute=-1.849465996e+00 lute=2.695119790e-07 wute=-8.885603135e-07 pute=2.430390169e-13
+  ua1=-5.513586527e-09 lua1=1.587511321e-15 wua1=6.698552446e-15 pua1=-1.832188065e-21
+  ub1=1.139923162e-17 lub1=-3.165505469e-24 wub1=-1.448182980e-23 pub1=3.961070087e-30
+  uc1=1.415567104e-10 luc1=-6.706915277e-17 wuc1=-4.893611081e-16 puc1=1.338500503e-22
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.1e-6
+  sbref=1.1e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.71 pmos
* Model Flag Parameters
+  lmin=1.5e-07 lmax=1.8e-07 wmin=1.12e-06 wmax=1.26e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-2.026e-8
+  vth0={-2.012588297e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=1.869012070e-07 wvth0=1.166804738e-06 pvth0=-2.319952351e-13
+  k1=8.834020042e+00 lk1=-1.475504562e-06 wk1=-9.625715118e-06 pk1=1.831502499e-12
+  k2=-4.002296001e+00 lk2=7.279894905e-07 wk2=4.708684266e-06 pk2=-9.036329708e-13
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=-3.953171858e+01 ldsub=7.683184320e-06 wdsub=4.951421662e-05 pdsub=-9.536921568e-12
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-1.468678060e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=2.325751313e-07 wvoff=1.351907020e-06 pvoff=-2.886889984e-13
+  nfactor={-2.856058106e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=6.306899747e-06 wnfactor=3.830539283e-05 pnfactor=-7.828578063e-12
+  eta0=-1.204350685e+01 leta0=2.267407894e-06 weta0=1.515167501e-05 peta0=-2.814469932e-12
+  etab=-8.140433274e-01 letab=1.273935020e-07 wetab=9.773536676e-07 petab=-1.581299870e-13
+  u0=6.770584239e-02 lu0=-1.269799543e-08 wu0=-7.992047989e-08 pu0=1.576166618e-14
+  ua=2.271061593e-08 lua=-4.927915198e-15 wua=-3.085817302e-14 pua=6.116883154e-21
+  ub=-2.153527282e-17 lub=4.652186127e-24 wub=2.904476001e-23 pub=-5.774628378e-30
+  uc=4.236636355e-10 luc=-1.084731164e-16 wuc=-5.462603366e-16 puc=1.346446422e-22
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=-4.819179497e+06 lvsat=9.295048592e-01 wvsat=6.076653651e+00 pvsat=-1.153768356e-6
+  a0=-1.299502796e+00 la0=-1.344218042e-08 wa0=2.430885730e-06 pa0=1.668540217e-14
+  ags=1.25
+  a1=0.0
+  a2=1.313083672e+01 la2=-2.610642825e-06 wa2=-1.549081880e-05 pa2=3.240517840e-12
+  b0=0.0
+  b1=0.0
+  keta=2.495586571e+00 lketa=-5.549600838e-07 wketa=-3.156696909e-06 pketa=6.888564132e-13
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-2.043510685e+00 lpclm=6.764649860e-07 wpclm=3.432789881e-06 ppclm=-8.396770461e-13
+  pdiblc1=-1.197285950e+01 lpdiblc1=2.700950650e-06 wpdiblc1=1.533874014e-05 ppdiblc1=-3.352614415e-12
+  pdiblc2=-3.633859218e-01 lpdiblc2=7.825717961e-08 wpdiblc2=4.608140158e-07 ppdiblc2=-9.713844585e-14
+  pdiblcb=-1.112727668e+01 lpdiblcb=2.245701320e-06 wpdiblcb=1.353269078e-05 ppdiblcb=-2.787526168e-12
+  drout=2.724583443e+01 ldrout=-5.623064737e-06 wdrout=-3.303580392e-05 pdrout=6.979752813e-12
+  pscbe1=800000000.0
+  pscbe2=1.134508762e-07 lpscbe2=-1.851677362e-14 wpscbe2=-1.293649057e-13 ppscbe2=2.298435263e-20
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=-4.932709054e+01 lbeta0=1.131180721e-05 wbeta0=7.169768377e-05 pbeta0=-1.404102956e-11
* Gidl Induced Drain Leakage Model Parameters
+  agidl=8.654312399e-15 lagidl=-1.908448970e-21 wagidl=-1.074235566e-20 pagidl=2.368904270e-27
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-1.106e-8
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.00074326333
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.5407449e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-1.381618242e+01 lkt1=2.504610677e-06 wkt1=1.626399281e-05 pkt1=-3.108903104e-12
+  kt2=-2.793217387e+00 lkt2=5.866591238e-07 wkt2=3.401180098e-06 pkt2=-7.282035440e-13
+  at=-1.588233631e+06 lat=3.186672556e-01 wat=2.007757002e+00 pat=-3.955527417e-7
+  ute=1.159905489e+01 lute=-2.673643544e-06 wute=-1.474389694e-05 pute=3.318718869e-12
+  ua1=2.971089011e-08 lua1=-6.047585647e-15 wua1=-3.634484151e-14 pua1=7.506698731e-21
+  ub1=-4.616634170e-17 lub1=9.264440486e-24 wub1=5.712903699e-23 pub1=-1.149969057e-29
+  uc1=4.721291063e-10 luc1=-1.455692554e-16 wuc1=-6.510721214e-16 puc1=1.806910408e-22
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.04e-6
+  sbref=1.04e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.72 pmos
* Model Flag Parameters
+  lmin=2.0e-05 lmax=0.0001 wmin=1.0e-06 wmax=1.12e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.135850030e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=9.541273302e-7
+  k1=4.276854265e-01 lk1=3.971117239e-7
+  k2=2.848051751e-02 lk2=-1.500844421e-7
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=-2.097023076e-06 lcit=2.422249835e-10 wcit=8.470329473e-28 pcit=-1.490777987e-31
+  voff={-2.351451054e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=4.628473774e-7
+  nfactor={1.892456558e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.556901933e-6
+  eta0=0.08
+  etab=-0.07
+  u0=9.728391786e-03 lu0=-1.420251827e-8
+  ua=-7.528013241e-10 lua=5.223392304e-16
+  ub=9.417519267e-19 lub=8.714072373e-25
+  uc=-1.141444728e-10 luc=8.483477603e-16
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=6.009393472e+04 lvsat=2.006678387e+0
+  a0=1.516922664e+00 la0=-5.293511136e-6
+  ags=8.145735879e-02 lags=3.184012825e-6
+  a1=0.0
+  a2=1.012549980e+00 la2=-4.255998776e-6
+  b0=-1.123676727e-07 lb0=2.249996341e-12
+  b1=4.233370455e-09 lb1=-8.476697797e-14
+  keta=2.967654180e-02 lketa=-6.316768153e-7
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-1.652677694e-02 lpclm=3.153419204e-06 ppclm=4.440892099e-28
+  pdiblc1=0.39
+  pdiblc2=1.516905606e-03 lpdiblc2=-2.398031945e-8
+  pdiblcb=-2.424906624e-01 lpdiblcb=1.749477616e-6
+  drout=0.56
+  pscbe1=8.000122018e+08 lpscbe1=-1.220470237e+0
+  pscbe2=1.122077829e-08 lpscbe2=-1.160426156e-13
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=-2.502940000e-11 lalpha0=2.503528691e-15
+  alpha1=-2.502940000e-11 lalpha1=2.503528691e-15
+  beta0=3.593732677e+01 lbeta0=-5.938723229e-04 pbeta0=9.094947018e-25
* Gidl Induced Drain Leakage Model Parameters
+  agidl=-3.146384318e-09 lagidl=3.241503941e-13 wagidl=1.654361225e-30 pagidl=-8.271806126e-35
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=-9.659333470e-02 legidl=1.966395734e-05 pegidl=-3.552713679e-27
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.376188837e-01 lkt1=-6.312647596e-8
+  kt2=-6.009470113e-02 lkt2=1.549065388e-7
+  at=8.875837106e+04 lat=-1.777255018e+0
+  ute=-7.064397988e-02 lute=-1.233892155e-6
+  ua1=2.157147563e-09 lua1=-6.696330892e-15
+  ub1=-1.357303605e-18 lub1=1.284338058e-23
+  uc1=-3.505211423e-11 luc1=5.264352112e-16 puc1=8.271806126e-37
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.73 pmos
* Model Flag Parameters
+  lmin=8.0e-06 lmax=2.0e-05 wmin=1.0e-06 wmax=1.12e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.0881997+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+  k1=0.44751769
+  k2=0.02098511
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-0.21202992+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.8147029+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+  eta0=0.08
+  etab=-0.07
+  u0=0.0090191
+  ua=-7.2671504e-10
+  ub=9.8527111e-19
+  uc=-7.1776909e-11
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=160310.0
+  a0=1.252558
+  ags=0.240471
+  a1=0.0
+  a2=0.8
+  b0=0.0
+  b1=0.0
+  keta=-0.0018702
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=0.14095898
+  pdiblc1=0.39
+  pdiblc2=0.00031929802
+  pdiblcb=-0.15511953
+  drout=0.56
+  pscbe1=799951250.0
+  pscbe2=5.4254628e-9
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=6.2785893
* Gidl Induced Drain Leakage Model Parameters
+  agidl=1.304209773e-8
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.88544965
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-0.4407715
+  kt2=-0.052358472
+  at=0.0
+  ute=-0.13226612
+  ua1=1.8227243e-9
+  ub1=-7.1588888e-19
+  uc1=-8.7612717e-12
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.74 pmos
* Model Flag Parameters
+  lmin=4.0e-06 lmax=8.0e-06 wmin=1.0e-06 wmax=1.12e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.090414346e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=1.776925644e-8
+  k1=4.556728822e-01 lk1=-6.543334786e-8
+  k2=1.885398624e-02 lk2=1.709911408e-8
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.057269452e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-5.057204472e-8
+  nfactor={2.150233085e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-2.692133146e-6
+  eta0=0.08
+  etab=-0.07
+  u0=8.535573484e-03 lu0=3.879584672e-9
+  ua=-8.237874492e-10 lua=7.788624164e-16
+  ub=1.048518672e-18 lub=-5.074680762e-25
+  uc=-7.083802061e-11 luc=-7.533189791e-18
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=2.678104074e+05 lvsat=-8.625316685e-01 wvsat=-4.656612873e-16
+  a0=1.347035279e+00 la0=-7.580403376e-7
+  ags=2.084960866e-01 lags=2.565513575e-7
+  a1=0.0
+  a2=0.8
+  b0=0.0
+  b1=0.0
+  keta=-8.364571240e-04 lketa=-8.294256640e-9
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=2.407132755e-01 lpclm=-8.003805848e-7
+  pdiblc1=0.39
+  pdiblc2=-1.397670217e-03 lpdiblc2=1.377612899e-08 wpdiblc2=-8.673617380e-25 ppdiblc2=-3.469446952e-30
+  pdiblcb=-2.494013897e-01 lpdiblcb=7.564723865e-7
+  drout=0.56
+  pscbe1=1.227212561e+09 lpscbe1=-3.428139670e+3
+  pscbe2=-1.711599940e-08 lpscbe2=1.808618728e-13 wpscbe2=-1.323488980e-29 ppscbe2=-1.058791184e-34
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=3.429576331e+00 lbeta0=2.285911254e-5
* Gidl Induced Drain Leakage Model Parameters
+  agidl=2.613220901e-08 lagidl=-1.050287696e-13
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=1.675517744e+00 legidl=-6.339127153e-6
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.061103840e-01 lkt1=-2.781041573e-7
+  kt2=-4.839276194e-02 lkt2=-3.181895402e-8
+  at=-9.120917488e+04 lat=7.318186388e-1
+  ute=-1.647219648e-01 lute=2.604101198e-7
+  ua1=5.703275549e-10 lua1=1.004863033e-14
+  ub1=8.239234094e-19 lub1=-1.235471470e-23 pub1=6.162975822e-45
+  uc1=-1.164852119e-11 luc1=2.316590399e-17
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.75 pmos
* Model Flag Parameters
+  lmin=2.0e-06 lmax=4.0e-06 wmin=1.0e-06 wmax=1.12e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.085843201e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-6.228379991e-10
+  k1=4.428072554e-01 lk1=-1.366824095e-8
+  k2=2.193345702e-02 lk2=4.708801823e-9
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=8.622137339e-01 ldsub=-1.215963003e-6
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.337857314e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=6.232304277e-8
+  nfactor={7.881674337e-01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=2.788165241e-6
+  eta0=1.604349200e-01 leta0=-3.236315093e-7
+  etab=-1.403185835e-01 letab=2.829282271e-7
+  u0=8.638994592e-03 lu0=3.463467775e-9
+  ua=-8.215637429e-10 lua=7.699152898e-16
+  ub=1.011504174e-18 lub=-3.585395030e-25
+  uc=-7.560382119e-11 luc=1.164210416e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=53438.0
+  a0=1.154071298e+00 la0=1.835409954e-8
+  ags=1.482758150e-01 lags=4.988488244e-7
+  a1=0.0
+  a2=0.8
+  b0=0.0
+  b1=0.0
+  keta=6.578345336e-03 lketa=-3.812786263e-08 pketa=-1.387778781e-29
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-5.559724103e-01 lpclm=2.405100206e-06 ppclm=-1.110223025e-27
+  pdiblc1=0.39
+  pdiblc2=3.641230659e-03 lpdiblc2=-6.497989463e-9
+  pdiblcb=-9.820554637e-02 lpdiblcb=1.481328872e-7
+  drout=0.56
+  pscbe1=-4.676991234e+07 lpscbe1=1.697754289e+3
+  pscbe2=4.653609693e-08 lpscbe2=-7.524360986e-14
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=1.147359093e+01 lbeta0=-9.506141085e-6
* Gidl Induced Drain Leakage Model Parameters
+  agidl=3.821637237e-11 lagidl=-3.906838872e-17
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.816142056e-01 lkt1=2.568697892e-8
+  kt2=-6.028632264e-02 lkt2=1.603502535e-8
+  at=1.022950518e+05 lat=-4.674948746e-2
+  ute=-1.327375183e-01 lute=1.317200597e-7
+  ua1=3.323674104e-09 lua1=-1.029514575e-15
+  ub1=-2.842323112e-18 lub1=2.396501504e-24
+  uc1=1.818504214e-11 luc1=-9.687003470e-17 puc1=-5.169878828e-38
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.76 pmos
* Model Flag Parameters
+  lmin=1.0e-06 lmax=2.0e-06 wmin=1.0e-06 wmax=1.12e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.101264296e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=3.058205737e-8
+  k1=3.540326720e-01 lk1=1.659689040e-7
+  k2=5.577749960e-02 lk2=-6.377529522e-08 pk2=-5.551115123e-29
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=-2.663045674e-01 ldsub=1.067616350e-6
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.021762939e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-1.639286090e-9
+  nfactor={2.430472285e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-5.350714714e-7
+  eta0=-2.241626400e-01 leta0=4.546093453e-07 weta0=-2.046973702e-22 peta0=2.237793284e-28
+  etab=8.442995791e-01 letab=-1.709466317e-06 wetab=1.908195824e-23 petab=-7.459310947e-28
+  u0=1.250070846e-02 lu0=-4.350787479e-9
+  ua=2.633023699e-11 lua=-9.458151364e-16
+  ub=5.976931819e-19 lub=4.788153150e-25
+  uc=-7.509174596e-11 luc=1.060590969e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=5.963848416e+04 lvsat=-1.254680371e-02 wvsat=1.164153218e-16
+  a0=1.369865781e+00 la0=-4.183103528e-7
+  ags=1.727992847e-01 lags=4.492250930e-7
+  a1=0.0
+  a2=5.953062352e-01 la2=4.142019269e-7
+  b0=0.0
+  b1=0.0
+  keta=-1.079934288e-02 lketa=-2.963762975e-9
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=4.550220723e-01 lpclm=3.593326501e-7
+  pdiblc1=7.492555200e-01 lpdiblc1=-7.269607298e-7
+  pdiblc2=0.00043
+  pdiblcb=-0.025
+  drout=1.096512000e-01 ldrout=9.112898038e-7
+  pscbe1=7.983183467e+08 lpscbe1=-1.229870506e+1
+  pscbe2=9.530520115e-09 lpscbe2=-3.620850560e-16
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=5.862313582e+00 lbeta0=1.848390856e-6
* Gidl Induced Drain Leakage Model Parameters
+  agidl=2.315918186e-11 lagidl=-8.599862589e-18
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.585366557e-01 lkt1=-2.101090483e-8
+  kt2=-5.625426130e-02 lkt2=7.876068592e-9
+  at=9.703221664e+04 lat=-3.610003518e-2
+  ute=9.359355551e-01 lute=-2.030761278e-06 wute=-4.440892099e-22 pute=1.110223025e-27
+  ua1=6.136533540e-09 lua1=-6.721391901e-15
+  ub1=-4.270929418e-18 lub1=5.287314936e-24
+  uc1=-1.285649500e-10 luc1=2.000815094e-16
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=2.75e-6
+  sbref=2.74e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.77 pmos
* Model Flag Parameters
+  lmin=5.0e-07 lmax=1.0e-06 wmin=1.0e-06 wmax=1.12e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.092537218e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=2.164971849e-8
+  k1=5.163486096e-01 lk1=-1.647044061e-10
+  k2=-1.189752607e-02 lk2=5.491447057e-9
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=1.315197776e+00 ldsub=-5.510829280e-7
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-1.991356383e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-4.751457949e-9
+  nfactor={1.798308567e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.119607376e-7
+  eta0=-6.270080000e-02 leta0=2.893499228e-7
+  etab=-1.689963224e+00 letab=8.844023472e-7
+  u0=9.894695136e-03 lu0=-1.683480718e-9
+  ua=-5.448939775e-10 lua=-3.611557284e-16
+  ub=8.616663893e-19 lub=2.086334578e-25
+  uc=-1.013764555e-10 luc=3.750883558e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=-6.051498240e+03 lvsat=5.468820708e-2
+  a0=1.217355653e+00 la0=-2.622131867e-7
+  ags=-5.662276614e-02 lags=6.840431505e-7
+  a1=0.0
+  a2=1.010355926e+00 la2=-1.060973294e-8
+  b0=0.0
+  b1=0.0
+  keta=1.145804192e-02 lketa=-2.574464147e-8
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=1.620957890e+00 lpclm=-8.340259780e-7
+  pdiblc1=6.831681950e-02 lpdiblc1=-3.000635109e-08 ppdiblc1=-5.551115123e-29
+  pdiblc2=8.382037816e-04 lpdiblc2=-4.178047345e-10
+  pdiblcb=-3.072820088e-02 lpdiblcb=5.862928163e-9
+  drout=1.0
+  pscbe1=7.719601783e+08 lpscbe1=1.467940745e+1
+  pscbe2=9.018239607e-09 lpscbe2=1.622442887e-16
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=6.533924275e+00 lbeta0=1.160983879e-6
* Gidl Induced Drain Leakage Model Parameters
+  agidl=1.669088570e-11 lagidl=-1.979432105e-18
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.172838726e-01 lkt1=-6.323395343e-8
+  kt2=-6.520102427e-02 lkt2=1.703325943e-8
+  at=8.968707775e+04 lat=-2.858213862e-2
+  ute=-1.937735245e+00 lute=9.104982595e-7
+  ua1=-3.568282344e-09 lua1=3.211681253e-15 pua1=-1.654361225e-36
+  ub1=4.385178260e-18 lub1=-3.572384395e-24 wub1=3.081487911e-39 pub1=3.081487911e-45
+  uc1=3.415037467e-10 luc1=-2.810432031e-16 wuc1=2.067951531e-31
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.75e-6
+  sbref=1.74e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.78 pmos
* Model Flag Parameters
+  lmin=2.5e-07 lmax=5.0e-07 wmin=1.0e-06 wmax=1.12e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.051387542e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=1.070397737e-10
+  k1=4.938004126e-01 lk1=1.163972768e-8
+  k2=-1.078294214e-03 lk2=-1.726372043e-10
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=-3.408496543e-01 ldsub=3.158910227e-07 pdsub=2.220446049e-28
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-7.666214318e-02+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-6.886878211e-8
+  nfactor={1.133414681e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=4.600459844e-7
+  eta0=0.49
+  etab=-1.301962000e-03 letab=3.544031462e-10
+  u0=7.405217482e-03 lu0=-3.801893760e-10
+  ua=-1.231304109e-09 lua=-1.806296181e-18
+  ub=1.265819661e-18 lub=-2.948863286e-27
+  uc=-6.230717731e-11 luc=1.705528707e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=9.676053951e+04 lvsat=8.640490753e-4
+  a0=8.514885312e-01 la0=-7.067443105e-8
+  ags=9.462833920e-01 lags=1.590017186e-7
+  a1=0.0
+  a2=1.198063207e+00 la2=-1.088782482e-7
+  b0=0.0
+  b1=0.0
+  keta=-4.253851648e-02 lketa=2.523636788e-9
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-6.403483396e-01 lpclm=3.498130593e-07 wpclm=-2.220446049e-22 ppclm=1.942890293e-28
+  pdiblc1=-4.242191933e-01 lpdiblc1=2.278461023e-07 wpdiblc1=2.220446049e-22 ppdiblc1=-3.469446952e-29
+  pdiblc2=-9.974276988e-03 lpdiblc2=5.242745198e-09 wpdiblc2=-5.312590645e-24 ppdiblc2=2.168404345e-30
+  pdiblcb=1.959588488e-01 lpdiblcb=-1.128122761e-07 ppdiblcb=-1.110223025e-28
+  drout=1.559003196e+00 ldrout=-2.926493531e-7
+  pscbe1=8.000316736e+08 lpscbe1=-1.658177145e-2
+  pscbe2=9.517713802e-09 lpscbe2=-9.924044155e-17
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=8.527171537e+00 lbeta0=1.174790728e-7
* Gidl Induced Drain Leakage Model Parameters
+  agidl=-6.515176521e-11 lagidl=4.086683250e-17 wagidl=-5.169878828e-32 pagidl=-2.584939414e-38
+  bgidl=7.151366880e+08 lbgidl=1.491316411e+2
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-5.606784192e-01 lkt1=1.183595963e-8
+  kt2=-1.043485456e-02 lkt2=-1.163792574e-8
+  at=-5.353157337e+03 lat=2.117332525e-2
+  ute=5.296362567e-01 lute=-3.812200691e-07 wute=4.440892099e-22
+  ua1=5.056715784e-09 lua1=-1.303677767e-15
+  ub1=-4.916272944e-18 lub1=1.297111340e-24
+  uc1=-2.956344010e-10 luc1=5.251136002e-17
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.25e-6
+  sbref=1.24e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.79 pmos
* Model Flag Parameters
+  lmin=1.8e-07 lmax=2.5e-07 wmin=1.0e-06 wmax=1.12e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.022413851e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-7.817844044e-9
+  k1=-6.490689072e-01 lk1=3.242373440e-7
+  k2=4.186502447e-01 lk2=-1.149767872e-07 wk2=-9.020562075e-23 pk2=6.765421556e-29
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=2.734546461e-01 ldsub=1.478665104e-7
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-1.926217918e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-3.715149901e-8
+  nfactor={3.480845624e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.820233270e-7
+  eta0=7.292390102e-01 leta0=-6.543665407e-8
+  etab=-6.25e-6
+  u0=1.636651887e-02 lu0=-2.831284531e-9
+  ua=2.341445631e-09 lua=-9.790248052e-16
+  ub=-1.366352887e-18 lub=7.170029723e-25
+  uc=2.876708666e-11 luc=-7.855345608e-18 wuc=1.494418099e-32 puc=3.029225876e-40
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=-8.298232454e+04 lvsat=5.002731725e-2
+  a0=-3.445166400e-01 la0=2.564569034e-7
+  ags=2.334702171e+00 lags=-2.207585859e-7
+  a1=0.0
+  a2=1.470082331e+00 la2=-1.832809193e-7
+  b0=0.0
+  b1=0.0
+  keta=1.782094629e-02 lketa=-1.398588347e-8
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=5.075991775e-01 lpclm=3.582645444e-8
+  pdiblc1=4.393230456e-01 lpdiblc1=-8.349970846e-9
+  pdiblc2=7.027921183e-03 lpdiblc2=5.923039542e-10
+  pdiblcb=-4.573434420e-01 lpdiblcb=6.587896648e-08 wpdiblcb=8.881784197e-22
+  drout=4.876068049e-01 ldrout=3.989877440e-10
+  pscbe1=7.998868799e+08 lpscbe1=2.302219403e-2
+  pscbe2=1.641780183e-08 lpscbe2=-1.986552518e-15
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=8.085587642e+00 lbeta0=2.382610996e-7
* Gidl Induced Drain Leakage Model Parameters
+  agidl=3.292360240e-10 lagidl=-6.700611560e-17
+  bgidl=2.017368972e+09 lbgidl=-2.070549331e+2
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-5.922187016e-01 lkt1=2.046285767e-8
+  kt2=-8.199556515e-02 lkt2=7.935359819e-9
+  at=1.327393562e+05 lat=-1.659773905e-2
+  ute=-2.656315088e+00 lute=4.902013427e-7
+  ua1=5.689729556e-10 lua1=-7.619034873e-17
+  ub1=-1.750861908e-18 lub1=4.313081131e-25 pub1=1.925929944e-46
+  uc1=-3.028031827e-10 luc1=5.447216517e-17
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.1e-6
+  sbref=1.1e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.80 pmos
* Model Flag Parameters
+  lmin=1.5e-07 lmax=1.8e-07 wmin=1.0e-06 wmax=1.12e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-2.026e-8
+  vth0={-9.530807322e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-2.376020697e-08 wvth0=-1.277295297e-12 pvth0=2.816691573e-19
+  k1=9.347669910e-02 lk1=1.875746915e-07 wk1=5.301943204e-13 pk1=-1.169184518e-19
+  k2=2.733816934e-01 lk2=-9.254616282e-08 wk2=1.398770824e-13 pk2=-3.084569400e-20
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=5.429215060e+00 ldsub=-9.767305050e-07 wdsub=-6.886389059e-13 pdsub=1.518586519e-19
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.410911288e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-2.956630085e-08 wvoff=-9.469666651e-14 pvoff=2.088250906e-20
+  nfactor={6.222243513e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-8.017607750e-07 wnfactor=4.204775175e-11 pnfactor=-9.272370221e-18
+  eta0=1.714843079e+00 leta0=-2.882479788e-07 weta0=-1.053348785e-11 peta0=2.322844741e-18
+  etab=7.343266554e-02 letab=-1.619474965e-08 wetab=1.205938537e-12 petab=-2.659335662e-19
+  u0=-4.865231863e-03 lu0=1.614244299e-09 wu0=1.219036599e-14 pu0=-2.688219508e-21
+  ua=-5.309870781e-09 lua=6.264656711e-16 wua=4.420573260e-21 pua=-9.748248146e-28
+  ub=4.838586734e-18 lub=-5.914191449e-25 wub=-3.304376911e-29 pub=7.286811969e-36
+  uc=-7.236340326e-11 luc=1.378979400e-17 wuc=3.524264629e-22 puc=-7.771708358e-29
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=6.986694175e+05 lvsat=-1.181637494e-01 wvsat=1.141271023e-06 pvsat=-2.516730856e-13
+  a0=9.078297385e-01 la0=1.711292876e-09 wa0=1.221508191e-11 pa0=-2.693669861e-18
+  ags=1.25
+  a1=0.0
+  a2=-9.354572783e-01 la2=3.318792433e-07 wa2=-3.071957693e-12 pa2=6.774281101e-19
+  b0=0.0
+  b1=0.0
+  keta=-3.708236724e-01 lketa=7.054978877e-08 wketa=4.318858799e-13 pketa=-9.523947420e-20
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=1.073601416e+00 lpclm=-8.599577991e-08 wpclm=1.603066288e-12 ppclm=-3.535081756e-19
+  pdiblc1=1.955357505e+00 lpdiblc1=-3.433633618e-07 wpdiblc1=-1.526007091e-11 ppdiblc1=3.365150837e-18
+  pdiblc2=5.505184156e-02 lpdiblc2=-9.948455892e-09 wpdiblc2=2.232371950e-13 ppdiblc2=-4.922826624e-20
+  pdiblcb=1.160916731e+00 lpdiblcb=-2.854769051e-07 wpdiblcb=4.744476804e-11 ppdiblcb=-1.046252025e-17
+  drout=-2.752067647e+00 ldrout=7.148453254e-07 wdrout=4.570065610e-11 pdrout=-1.007790868e-17
+  pscbe1=800000000.0
+  pscbe2=-4.017537105e-09 lpscbe2=2.353911941e-15 wpscbe2=-2.312525422e-19 ppscbe2=5.099581060e-26
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=1.577731231e+01 lbeta0=-1.438016104e-06 wbeta0=2.784057813e-11 pbeta0=-6.139404277e-18
* Gidl Induced Drain Leakage Model Parameters
+  agidl=-1.009669780e-14 lagidl=2.226523799e-21 wagidl=9.907606842e-21 pagidl=-2.184825461e-27
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-1.106e-8
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=9.521864647e-01 lkt1=-3.184001097e-07 wkt1=1.673981799e-12 pkt1=-3.691464681e-19
+  kt2=2.951914855e-01 lkt2=-7.457908898e-08 wkt2=1.881265177e-12 pkt2=-4.148565971e-19
+  at=2.348924372e+05 lat=-4.051094353e-02 wat=-6.893663919e-07 pat=1.520190769e-13
+  ute=-1.789002428e+00 lute=3.398880113e-07 wute=-4.290497671e-12 pute=9.461405459e-19
+  ua1=-3.291682485e-09 lua1=7.687972189e-16 wua1=-3.237671200e-20 pua1=7.139712529e-27
+  ub1=5.709125795e-18 lub1=-1.177741263e-24 wub1=3.714888582e-29 pub1=-8.192072300e-36
+  uc1=-1.190733596e-10 luc1=1.850611769e-17 wuc1=2.600610619e-21 puc1=-5.734866538e-28
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.04e-6
+  sbref=1.04e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.81 pmos
* Model Flag Parameters
+  lmin=2.0e-05 lmax=0.0001 wmin=9.4e-07 wmax=1.0e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.135850030e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=9.541273302e-7
+  k1=4.276854265e-01 lk1=3.971117239e-7
+  k2=2.848051751e-02 lk2=-1.500844421e-7
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=-2.097023076e-06 lcit=2.422249835e-10 wcit=-2.541098842e-27 pcit=-8.131516294e-32
+  voff={-2.351451054e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=4.628473774e-7
+  nfactor={1.892456558e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.556901933e-6
+  eta0=0.08
+  etab=-0.07
+  u0=9.728391786e-03 lu0=-1.420251827e-8
+  ua=-7.528013241e-10 lua=5.223392304e-16
+  ub=9.417519267e-19 lub=8.714072373e-25
+  uc=-1.141444728e-10 luc=8.483477603e-16
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=6.009393472e+04 lvsat=2.006678387e+0
+  a0=1.516922664e+00 la0=-5.293511136e-06 wa0=3.552713679e-21
+  ags=8.145735879e-02 lags=3.184012825e-6
+  a1=0.0
+  a2=1.012549980e+00 la2=-4.255998776e-6
+  b0=-1.123676727e-07 lb0=2.249996341e-12
+  b1=4.233370455e-09 lb1=-8.476697797e-14
+  keta=2.967654180e-02 lketa=-6.316768153e-7
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-1.652677694e-02 lpclm=3.153419204e-06 ppclm=1.776356839e-27
+  pdiblc1=0.39
+  pdiblc2=1.516905606e-03 lpdiblc2=-2.398031945e-8
+  pdiblcb=-2.424906624e-01 lpdiblcb=1.749477616e-6
+  drout=0.56
+  pscbe1=8.000122018e+08 lpscbe1=-1.220470237e+0
+  pscbe2=1.122077829e-08 lpscbe2=-1.160426156e-13
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=-2.502940000e-11 lalpha0=2.503528691e-15
+  alpha1=-2.502940000e-11 lalpha1=2.503528691e-15
+  beta0=3.593732677e+01 lbeta0=-5.938723229e-4
* Gidl Induced Drain Leakage Model Parameters
+  agidl=-3.146384318e-09 lagidl=3.241503941e-13 wagidl=-8.271806126e-31 pagidl=-1.323488980e-34
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=-9.659333470e-02 legidl=1.966395734e-05 pegidl=1.421085472e-26
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.376188837e-01 lkt1=-6.312647596e-8
+  kt2=-6.009470113e-02 lkt2=1.549065388e-7
+  at=8.875837106e+04 lat=-1.777255018e+0
+  ute=-7.064397988e-02 lute=-1.233892155e-06 wute=-2.220446049e-22
+  ua1=2.157147563e-09 lua1=-6.696330892e-15
+  ub1=-1.357303605e-18 lub1=1.284338058e-23
+  uc1=-3.505211423e-11 luc1=5.264352112e-16
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.82 pmos
* Model Flag Parameters
+  lmin=8.0e-06 lmax=2.0e-05 wmin=9.4e-07 wmax=1.0e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.0881997+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+  k1=0.44751769
+  k2=0.02098511
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-0.21202992+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.8147029+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+  eta0=0.08
+  etab=-0.07
+  u0=0.0090191
+  ua=-7.2671504e-10
+  ub=9.8527111e-19
+  uc=-7.1776909e-11
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=160310.0
+  a0=1.252558
+  ags=0.240471
+  a1=0.0
+  a2=0.8
+  b0=0.0
+  b1=0.0
+  keta=-0.0018702
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=0.14095898
+  pdiblc1=0.39
+  pdiblc2=0.00031929802
+  pdiblcb=-0.15511953
+  drout=0.56
+  pscbe1=799951250.0
+  pscbe2=5.4254628e-9
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=6.2785893
* Gidl Induced Drain Leakage Model Parameters
+  agidl=1.304209773e-8
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.88544965
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-0.4407715
+  kt2=-0.052358472
+  at=0.0
+  ute=-0.13226612
+  ua1=1.8227243e-9
+  ub1=-7.1588888e-19
+  uc1=-8.7612717e-12
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.83 pmos
* Model Flag Parameters
+  lmin=4.0e-06 lmax=8.0e-06 wmin=9.4e-07 wmax=1.0e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.090414346e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=1.776925644e-8
+  k1=4.556728822e-01 lk1=-6.543334786e-8
+  k2=1.885398624e-02 lk2=1.709911408e-8
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.057269452e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-5.057204472e-8
+  nfactor={2.150233085e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-2.692133146e-6
+  eta0=0.08
+  etab=-0.07
+  u0=8.535573484e-03 lu0=3.879584672e-9
+  ua=-8.237874492e-10 lua=7.788624164e-16
+  ub=1.048518672e-18 lub=-5.074680762e-25
+  uc=-7.083802061e-11 luc=-7.533189791e-18
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=2.678104074e+05 lvsat=-8.625316685e-1
+  a0=1.347035279e+00 la0=-7.580403376e-7
+  ags=2.084960866e-01 lags=2.565513575e-7
+  a1=0.0
+  a2=0.8
+  b0=0.0
+  b1=0.0
+  keta=-8.364571240e-04 lketa=-8.294256640e-9
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=2.407132755e-01 lpclm=-8.003805848e-7
+  pdiblc1=0.39
+  pdiblc2=-1.397670217e-03 lpdiblc2=1.377612899e-8
+  pdiblcb=-2.494013897e-01 lpdiblcb=7.564723865e-7
+  drout=0.56
+  pscbe1=1.227212561e+09 lpscbe1=-3.428139670e+03 wpscbe1=-3.814697266e-12
+  pscbe2=-1.711599940e-08 lpscbe2=1.808618728e-13 wpscbe2=2.646977960e-29 ppscbe2=-1.058791184e-34
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=3.429576331e+00 lbeta0=2.285911254e-5
* Gidl Induced Drain Leakage Model Parameters
+  agidl=2.613220901e-08 lagidl=-1.050287696e-13
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=1.675517744e+00 legidl=-6.339127153e-06 pegidl=-1.421085472e-26
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.061103840e-01 lkt1=-2.781041573e-7
+  kt2=-4.839276194e-02 lkt2=-3.181895402e-8
+  at=-9.120917488e+04 lat=7.318186388e-1
+  ute=-1.647219648e-01 lute=2.604101198e-7
+  ua1=5.703275549e-10 lua1=1.004863033e-14
+  ub1=8.239234094e-19 lub1=-1.235471470e-23 pub1=1.232595164e-44
+  uc1=-1.164852119e-11 luc1=2.316590399e-17
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.84 pmos
* Model Flag Parameters
+  lmin=2.0e-06 lmax=4.0e-06 wmin=9.4e-07 wmax=1.0e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.085843201e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-6.228379991e-10
+  k1=4.428072554e-01 lk1=-1.366824095e-8
+  k2=2.193345702e-02 lk2=4.708801823e-9
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=8.622137339e-01 ldsub=-1.215963003e-6
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.337857314e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=6.232304277e-8
+  nfactor={7.881674337e-01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=2.788165241e-6
+  eta0=1.604349200e-01 leta0=-3.236315093e-7
+  etab=-1.403185835e-01 letab=2.829282271e-7
+  u0=8.638994592e-03 lu0=3.463467775e-9
+  ua=-8.215637429e-10 lua=7.699152898e-16
+  ub=1.011504174e-18 lub=-3.585395030e-25
+  uc=-7.560382119e-11 luc=1.164210416e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=53438.0
+  a0=1.154071298e+00 la0=1.835409954e-8
+  ags=1.482758150e-01 lags=4.988488244e-7
+  a1=0.0
+  a2=0.8
+  b0=0.0
+  b1=0.0
+  keta=6.578345336e-03 lketa=-3.812786263e-08 pketa=-2.775557562e-29
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-5.559724103e-01 lpclm=2.405100206e-06 wpclm=-4.440892099e-22 ppclm=2.220446049e-27
+  pdiblc1=0.39
+  pdiblc2=3.641230659e-03 lpdiblc2=-6.497989463e-9
+  pdiblcb=-9.820554637e-02 lpdiblcb=1.481328872e-7
+  drout=0.56
+  pscbe1=-4.676991234e+07 lpscbe1=1.697754289e+3
+  pscbe2=4.653609693e-08 lpscbe2=-7.524360986e-14 ppscbe2=-2.117582368e-34
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=1.147359093e+01 lbeta0=-9.506141085e-6
* Gidl Induced Drain Leakage Model Parameters
+  agidl=3.821637237e-11 lagidl=-3.906838872e-17
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.816142056e-01 lkt1=2.568697892e-8
+  kt2=-6.028632264e-02 lkt2=1.603502535e-8
+  at=1.022950518e+05 lat=-4.674948746e-2
+  ute=-1.327375183e-01 lute=1.317200597e-7
+  ua1=3.323674104e-09 lua1=-1.029514575e-15
+  ub1=-2.842323112e-18 lub1=2.396501504e-24
+  uc1=1.818504214e-11 luc1=-9.687003470e-17 wuc1=2.584939414e-32
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.85 pmos
* Model Flag Parameters
+  lmin=1.0e-06 lmax=2.0e-06 wmin=9.4e-07 wmax=1.0e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.101264296e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=3.058205737e-8
+  k1=3.540326720e-01 lk1=1.659689040e-7
+  k2=5.577749960e-02 lk2=-6.377529522e-8
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=-2.663045674e-01 ldsub=1.067616350e-06 pdsub=-1.776356839e-27
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.021762939e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-1.639286090e-9
+  nfactor={2.430472285e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-5.350714714e-7
+  eta0=-2.241626400e-01 leta0=4.546093453e-07 weta0=-1.249000903e-22 peta0=-8.673617380e-30
+  etab=8.442995791e-01 letab=-1.709466317e-06 wetab=-8.569533971e-22 petab=-9.540979118e-28
+  u0=1.250070846e-02 lu0=-4.350787479e-9
+  ua=2.633023699e-11 lua=-9.458151364e-16
+  ub=5.976931819e-19 lub=4.788153150e-25
+  uc=-7.509174596e-11 luc=1.060590969e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=5.963848416e+04 lvsat=-1.254680371e-2
+  a0=1.369865781e+00 la0=-4.183103528e-7
+  ags=1.727992847e-01 lags=4.492250930e-7
+  a1=0.0
+  a2=5.953062352e-01 la2=4.142019269e-7
+  b0=0.0
+  b1=0.0
+  keta=-1.079934288e-02 lketa=-2.963762975e-9
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=4.550220723e-01 lpclm=3.593326501e-7
+  pdiblc1=7.492555200e-01 lpdiblc1=-7.269607298e-7
+  pdiblc2=0.00043
+  pdiblcb=-0.025
+  drout=1.096512000e-01 ldrout=9.112898038e-7
+  pscbe1=7.983183467e+08 lpscbe1=-1.229870506e+1
+  pscbe2=9.530520115e-09 lpscbe2=-3.620850560e-16
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=5.862313582e+00 lbeta0=1.848390856e-6
* Gidl Induced Drain Leakage Model Parameters
+  agidl=2.315918186e-11 lagidl=-8.599862589e-18
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.585366557e-01 lkt1=-2.101090483e-8
+  kt2=-5.625426130e-02 lkt2=7.876068592e-9
+  at=9.703221664e+04 lat=-3.610003518e-2
+  ute=9.359355551e-01 lute=-2.030761278e-06 wute=-8.881784197e-22
+  ua1=6.136533540e-09 lua1=-6.721391901e-15
+  ub1=-4.270929418e-18 lub1=5.287314936e-24 wub1=-6.162975822e-39 pub1=-6.162975822e-45
+  uc1=-1.285649500e-10 luc1=2.000815094e-16 puc1=1.033975766e-37
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=2.75e-6
+  sbref=2.74e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.86 pmos
* Model Flag Parameters
+  lmin=5.0e-07 lmax=1.0e-06 wmin=9.4e-07 wmax=1.0e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.092537218e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=2.164971849e-8
+  k1=5.163486096e-01 lk1=-1.647044061e-10
+  k2=-1.189752607e-02 lk2=5.491447057e-9
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=1.315197776e+00 ldsub=-5.510829280e-07 pdsub=-1.776356839e-27
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-1.991356383e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-4.751457949e-9
+  nfactor={1.798308567e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.119607376e-7
+  eta0=-6.270080000e-02 leta0=2.893499228e-07 peta0=4.440892099e-28
+  etab=-1.689963224e+00 letab=8.844023472e-7
+  u0=9.894695136e-03 lu0=-1.683480718e-9
+  ua=-5.448939775e-10 lua=-3.611557284e-16
+  ub=8.616663893e-19 lub=2.086334578e-25
+  uc=-1.013764555e-10 luc=3.750883558e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=-6.051498240e+03 lvsat=5.468820708e-2
+  a0=1.217355653e+00 la0=-2.622131867e-7
+  ags=-5.662276614e-02 lags=6.840431505e-7
+  a1=0.0
+  a2=1.010355926e+00 la2=-1.060973294e-8
+  b0=0.0
+  b1=0.0
+  keta=1.145804192e-02 lketa=-2.574464147e-8
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=1.620957890e+00 lpclm=-8.340259780e-7
+  pdiblc1=6.831681950e-02 lpdiblc1=-3.000635109e-8
+  pdiblc2=8.382037816e-04 lpdiblc2=-4.178047345e-10
+  pdiblcb=-3.072820088e-02 lpdiblcb=5.862928163e-9
+  drout=1.0
+  pscbe1=7.719601783e+08 lpscbe1=1.467940745e+1
+  pscbe2=9.018239607e-09 lpscbe2=1.622442887e-16
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=6.533924275e+00 lbeta0=1.160983879e-6
* Gidl Induced Drain Leakage Model Parameters
+  agidl=1.669088570e-11 lagidl=-1.979432105e-18
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.172838726e-01 lkt1=-6.323395343e-8
+  kt2=-6.520102427e-02 lkt2=1.703325943e-8
+  at=8.968707775e+04 lat=-2.858213862e-02 wat=-2.328306437e-16
+  ute=-1.937735245e+00 lute=9.104982595e-7
+  ua1=-3.568282344e-09 lua1=3.211681253e-15 wua1=-1.654361225e-30
+  ub1=4.385178260e-18 lub1=-3.572384395e-24 wub1=-3.081487911e-39 pub1=-3.081487911e-45
+  uc1=3.415037467e-10 luc1=-2.810432031e-16 puc1=2.067951531e-37
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.75e-6
+  sbref=1.74e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.87 pmos
* Model Flag Parameters
+  lmin=2.5e-07 lmax=5.0e-07 wmin=9.4e-07 wmax=1.0e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.051387542e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=1.070397737e-10
+  k1=4.938004126e-01 lk1=1.163972768e-8
+  k2=-1.078294214e-03 lk2=-1.726372043e-10
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=-3.408496543e-01 ldsub=3.158910227e-07 pdsub=4.440892099e-28
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-7.666214318e-02+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-6.886878211e-8
+  nfactor={1.133414681e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=4.600459844e-7
+  eta0=0.49
+  etab=-1.301962000e-03 letab=3.544031462e-10
+  u0=7.405217482e-03 lu0=-3.801893760e-10
+  ua=-1.231304109e-09 lua=-1.806296181e-18
+  ub=1.265819661e-18 lub=-2.948863286e-27
+  uc=-6.230717731e-11 luc=1.705528707e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=9.676053951e+04 lvsat=8.640490753e-4
+  a0=8.514885312e-01 la0=-7.067443105e-8
+  ags=9.462833920e-01 lags=1.590017186e-7
+  a1=0.0
+  a2=1.198063207e+00 la2=-1.088782482e-7
+  b0=0.0
+  b1=0.0
+  keta=-4.253851648e-02 lketa=2.523636788e-9
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-6.403483396e-01 lpclm=3.498130593e-07 wpclm=2.220446049e-22 ppclm=-1.387778781e-28
+  pdiblc1=-4.242191933e-01 lpdiblc1=2.278461023e-07 wpdiblc1=-5.551115123e-23 ppdiblc1=1.387778781e-29
+  pdiblc2=-9.974276988e-03 lpdiblc2=5.242745198e-09 wpdiblc2=-9.974659987e-24 ppdiblc2=-6.884683795e-30
+  pdiblcb=1.959588488e-01 lpdiblcb=-1.128122761e-07 wpdiblcb=-1.110223025e-22 ppdiblcb=-5.551115123e-29
+  drout=1.559003196e+00 ldrout=-2.926493531e-7
+  pscbe1=8.000316736e+08 lpscbe1=-1.658177145e-2
+  pscbe2=9.517713802e-09 lpscbe2=-9.924044155e-17
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=8.527171537e+00 lbeta0=1.174790728e-7
* Gidl Induced Drain Leakage Model Parameters
+  agidl=-6.515176521e-11 lagidl=4.086683250e-17 pagidl=2.584939414e-38
+  bgidl=7.151366880e+08 lbgidl=1.491316411e+2
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-5.606784192e-01 lkt1=1.183595963e-8
+  kt2=-1.043485456e-02 lkt2=-1.163792574e-8
+  at=-5.353157337e+03 lat=2.117332525e-2
+  ute=5.296362567e-01 lute=-3.812200691e-07 pute=2.220446049e-28
+  ua1=5.056715784e-09 lua1=-1.303677767e-15 wua1=1.323488980e-29
+  ub1=-4.916272944e-18 lub1=1.297111340e-24
+  uc1=-2.956344010e-10 luc1=5.251136002e-17
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.25e-6
+  sbref=1.24e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.88 pmos
* Model Flag Parameters
+  lmin=1.8e-07 lmax=2.5e-07 wmin=9.4e-07 wmax=1.0e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.022413851e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-7.817844044e-9
+  k1=-6.490689072e-01 lk1=3.242373440e-7
+  k2=4.186502447e-01 lk2=-1.149767872e-07 wk2=-2.359223927e-22 pk2=-3.122502257e-29
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=2.734546461e-01 ldsub=1.478665104e-7
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-1.926217918e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-3.715149901e-8
+  nfactor={3.480845624e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.820233270e-7
+  eta0=7.292390102e-01 leta0=-6.543665407e-8
+  etab=-6.25e-6
+  u0=1.636651887e-02 lu0=-2.831284531e-9
+  ua=2.341445631e-09 lua=-9.790248052e-16
+  ub=-1.366352887e-18 lub=7.170029723e-25
+  uc=2.876708666e-11 luc=-7.855345608e-18 wuc=-1.332859385e-32 puc=4.038967835e-40
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=-8.298232454e+04 lvsat=5.002731725e-2
+  a0=-3.445166400e-01 la0=2.564569034e-7
+  ags=2.334702171e+00 lags=-2.207585859e-7
+  a1=0.0
+  a2=1.470082331e+00 la2=-1.832809193e-7
+  b0=0.0
+  b1=0.0
+  keta=1.782094629e-02 lketa=-1.398588347e-8
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=5.075991775e-01 lpclm=3.582645444e-8
+  pdiblc1=4.393230456e-01 lpdiblc1=-8.349970846e-9
+  pdiblc2=7.027921183e-03 lpdiblc2=5.923039542e-10
+  pdiblcb=-4.573434420e-01 lpdiblcb=6.587896648e-8
+  drout=4.876068049e-01 ldrout=3.989877440e-10
+  pscbe1=7.998868799e+08 lpscbe1=2.302219403e-2
+  pscbe2=1.641780183e-08 lpscbe2=-1.986552518e-15
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=8.085587642e+00 lbeta0=2.382610996e-7
* Gidl Induced Drain Leakage Model Parameters
+  agidl=3.292360240e-10 lagidl=-6.700611560e-17
+  bgidl=2.017368972e+09 lbgidl=-2.070549331e+2
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-5.922187016e-01 lkt1=2.046285767e-8
+  kt2=-8.199556515e-02 lkt2=7.935359819e-9
+  at=1.327393562e+05 lat=-1.659773905e-2
+  ute=-2.656315088e+00 lute=4.902013427e-7
+  ua1=5.689729556e-10 lua1=-7.619034873e-17
+  ub1=-1.750861908e-18 lub1=4.313081131e-25 wub1=-1.540743956e-39
+  uc1=-3.028031827e-10 luc1=5.447216517e-17
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.1e-6
+  sbref=1.1e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.89 pmos
* Model Flag Parameters
+  lmin=1.5e-07 lmax=1.8e-07 wmin=9.4e-07 wmax=1.0e-6
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-2.026e-8
+  vth0={-1.854947105e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-1.930282765e-07 wvth0=-7.532119480e-07 pvth0=1.660982988e-13
+  k1=1.159348757e+00 lk1=-4.747141476e-08 wk1=-1.045909876e-06 pk1=2.306440459e-13
+  k2=-1.263501225e+00 lk2=2.463672584e-07 wk2=1.508100315e-06 pk2=-3.325662815e-13
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=5.663696152e+00 ldsub=-1.028438276e-06 wdsub=-2.300904192e-07 pdsub=5.073953924e-14
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={1.086694184e+01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-2.479109731e-06 wvoff=-1.090000182e-05 pvoff=2.403668401e-12
+  nfactor={1.329749387e+02+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-2.875326513e-05 wnfactor=-1.243788287e-04 pnfactor=2.742801931e-11
+  eta0=2.288232837e+00 leta0=-4.146918883e-07 weta0=-5.626618484e-07 peta0=1.240781908e-13
+  etab=-4.415447927e-01 letab=9.736807943e-08 wetab=5.053341663e-07 petab=-1.114362904e-13
+  u0=-5.925721101e-02 lu0=1.360876354e-08 wu0=5.337333835e-08 pu0=-1.176988857e-14
+  ua=-1.563364139e-08 lua=2.903063565e-15 wua=1.013043145e-14 pua=-2.233962743e-21
+  ub=1.489481188e-17 lub=-2.809017914e-24 wub=-9.867925205e-24 pub=2.176074866e-30
+  uc=-7.009672971e-11 luc=1.328994715e-17 wuc=-2.223870863e-18 puc=4.904080028e-25
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=7.111518667e+06 lvsat=-1.532325266e+00 wvsat=-6.292748268e+00 pvsat=1.387676848e-6
+  a0=7.964908362e+00 la0=-1.554515685e-06 wa0=-6.924901440e-06 pa0=1.527079266e-12
+  ags=1.250000031e+00 lags=-6.888562609e-15 wags=-3.065278520e-14 pags=6.759552917e-21
+  a1=0.0
+  a2=-6.193528785e+00 la2=1.491389172e-06 wa2=5.159595272e-06 pa2=-1.137793949e-12
+  b0=0.0
+  b1=0.0
+  keta=-3.285561737e-01 lketa=6.122895995e-08 wketa=-4.147548110e-08 pketa=9.146173093e-15
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=1.068705626e+00 lpclm=-8.491616029e-08 wpclm=4.805704761e-09 ppclm=-1.059754014e-15
+  pdiblc1=2.431710580e+00 lpdiblc1=-4.484087421e-07 wpdiblc1=-4.674471955e-07 ppdiblc1=1.030814556e-13
+  pdiblc2=8.845274624e-02 lpdiblc2=-1.731402339e-08 wpdiblc2=-3.277514930e-08 ppdiblc2=7.227575924e-15
+  pdiblcb=-2.142488265e-01 lpdiblcb=1.777460366e-08 wpdiblcb=1.349458902e-06 ppdiblcb=-2.975826770e-13
+  drout=-2.752021545e+00 ldrout=7.148351589e-07 wdrout=4.616423723e-13 pdrout=-1.018013762e-19
+  pscbe1=7.999999952e+08 lpscbe1=1.063938141e-06 wpscbe1=4.734329224e-06 ppscbe1=-1.044012070e-12
+  pscbe2=-3.529479812e-08 lpscbe2=9.251173540e-15 wpscbe2=3.069126922e-14 ppscbe2=-6.768038688e-21
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=1.975419248e+01 lbeta0=-2.314997720e-06 wbeta0=-3.902373325e-06 pbeta0=8.605513655e-13
* Gidl Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=9.999999966e+08 lbgidl=7.578430176e-07 wbgidl=3.372238159e-06 pbgidl=-7.436447144e-13
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-1.106e-8
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=1.682597805e+01 lkt1=-3.818888630e-06 wkt1=-1.557650554e-05 pkt1=3.434931003e-12
+  kt2=2.951933965e-01 lkt2=-7.457951039e-08 wkt2=6.077740977e-15 pkt2=-1.340263456e-21
+  at=8.542471780e+05 lat=-1.770910510e-01 wat=-6.077561546e-01 pat=1.340223872e-7
+  ute=-3.255901161e+00 lute=6.633685200e-07 wute=1.439422363e-06 pute=-3.174214196e-13
+  ua1=-3.291715626e-09 lua1=7.688045271e-16 wua1=1.437063525e-22 pua1=-3.169012555e-29
+  ub1=5.709164458e-18 lub1=-1.177749789e-24 wub1=-7.894836554e-31 pub1=1.740969349e-37
+  uc1=-1.190706991e-10 luc1=1.850553099e-17 wuc1=-1.008935768e-23 puc1=2.224905020e-30
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.04e-6
+  sbref=1.04e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.90 pmos
* Model Flag Parameters
+  lmin=2.0e-05 lmax=0.0001 wmin=8.6e-07 wmax=9.4e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.236161512e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=1.098763492e-05 wvth0=9.241416025e-08 pvth0=-9.243589606e-12
+  k1=3.859353744e-01 lk1=4.573098901e-06 wk1=3.846315405e-08 pk1=-3.847220059e-12
+  k2=4.425953613e-02 lk2=-1.728357427e-06 wk2=-1.453676804e-08 pk2=1.454018709e-12
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=-2.756317048e-05 lcit=2.789438687e-09 wcit=2.346124855e-11 pcit=-2.346676663e-15
+  voff={-2.838062277e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=5.330104114e-06 wvoff=4.483012943e-08 pvoff=-4.484067348e-12
+  nfactor={2.056140310e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.792912697e-05 wnfactor=-1.507972576e-07 pnfactor=1.508327251e-11
+  eta0=0.08
+  etab=-0.07
+  u0=1.122156321e-02 lu0=-1.635547801e-07 wu0=-1.375617025e-09 pu0=1.375940570e-13
+  ua=-8.077170790e-10 lua=6.015206344e-15 wua=5.059234739e-17 pua=-5.060424671e-21
+  ub=8.501371608e-19 lub=1.003503860e-23 wub=8.440211859e-26 pub=-8.442196996e-30
+  uc=-2.033348973e-10 luc=9.769487972e-15 wuc=8.216864079e-17 puc=-8.218796685e-21
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=-1.508767375e+05 lvsat=2.310870764e+01 wvsat=1.943613732e-01 pvsat=-1.944070869e-5
+  a0=2.073452106e+00 la0=-6.095954489e-05 wa0=-5.127149919e-07 pa0=5.128355825e-11
+  ags=-2.532915130e-01 lags=3.666677329e-05 wags=3.083947626e-07 pags=-3.084672970e-11
+  a1=0.0
+  a2=1.460001315e+00 la2=-4.901165630e-05 wa2=-4.122243860e-07 pa2=4.123213412e-11
+  b0=-3.489194009e-07 lb0=2.591073286e-11 wb0=2.179284838e-13 pb0=-2.179797406e-17
+  b1=1.314528501e-08 lb1=-9.761680415e-13 wb1=-8.210297345e-15 pb1=8.212228406e-19
+  keta=9.608742418e-02 lketa=-7.274327038e-06 wketa=-6.118248644e-08 pketa=6.119687656e-12
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-3.480592106e-01 lpclm=3.631446021e-05 wpclm=3.054315482e-07 ppclm=-3.055033857e-11
+  pdiblc1=0.39
+  pdiblc2=4.038059044e-03 lpdiblc2=-2.761549608e-07 wpdiblc2=-2.322668070e-09 ppdiblc2=2.323214362e-13
+  pdiblcb=-4.264207187e-01 lpdiblcb=2.014680928e-05 wpdiblcb=1.694496108e-07 ppdiblcb=-1.694894654e-11
+  drout=0.56
+  pscbe1=8.001405151e+08 lpscbe1=-1.405481320e+01 wpscbe1=-1.182114048e-01 ppscbe1=1.182392081e-5
+  pscbe2=2.342083425e-08 lpscbe2=-1.336335157e-12 wpscbe2=-1.123956995e-14 ppscbe2=1.124221350e-18
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=-2.882360675e-10 lalpha0=2.883038606e-14 walpha0=2.424849329e-16 palpha0=-2.425419654e-20
+  alpha1=-2.882360675e-10 lalpha1=2.883038606e-14 walpha1=2.424849329e-16 palpha1=-2.425419654e-20
+  beta0=9.837366135e+01 lbeta0=-6.838974283e-03 wbeta0=-5.752084683e-05 pbeta0=5.753437573e-9
* Gidl Induced Drain Leakage Model Parameters
+  agidl=-3.722570015e-08 lagidl=3.732883523e-12 wagidl=3.139631946e-14 pagidl=-3.140370387e-18
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=-2.163949183e+00 legidl=2.264481664e-04 wegidl=1.904597057e-06 pegidl=-1.905045018e-10
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.309821276e-01 lkt1=-7.269581845e-07 wkt1=-6.114257584e-09 pkt1=6.115695658e-13
+  kt2=-7.638068738e-02 lkt2=1.783888210e-06 wkt2=1.500382312e-08 pkt2=-1.500735202e-12
+  at=2.756087843e+05 lat=-2.046669106e+01 wat=-1.721400539e-01 pat=1.721805412e-5
+  ute=5.908037409e-02 lute=-1.420937867e-05 wute=-1.195114150e-07 pute=1.195395241e-11
+  ua1=2.861161439e-09 lua1=-7.711427692e-14 wua1=-6.485882718e-16 pua1=6.487408197e-20
+  ub1=-2.707583078e-18 lub1=1.479030864e-22 wub1=1.243974670e-24 pub1=-1.244267253e-28
+  uc1=-9.039849713e-11 luc1=6.062375248e-15 wuc1=5.098907287e-17 puc1=-5.100106550e-21
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.91 pmos
* Model Flag Parameters
+  lmin=8.0e-06 lmax=2.0e-05 wmin=8.6e-07 wmax=9.4e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-4.194564823e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-5.365674582e-06 wvth0=-6.160944017e-07 pvth0=4.943245754e-12
+  k1=7.258513711e-01 lk1=-2.233215857e-06 wk1=-2.564210270e-07 pk1=2.057399239e-12
+  k2=-8.420834747e-02 lk2=8.440218099e-07 wk2=9.691178695e-08 pk2=-7.775736608e-13
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.797743160e-04 lcit=-1.362187620e-09 wcit=-1.564083237e-10 pcit=1.254945313e-15
+  voff={1.123775618e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-2.602889918e-06 wvoff=-2.988675296e-07 pvoff=2.397969601e-12
+  nfactor={7.234778868e-01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=8.755465718e-06 wnfactor=1.005315050e-06 pnfactor=-8.066165413e-12
+  eta0=0.08
+  etab=-0.07
+  u0=-9.353761633e-04 lu0=7.986993859e-08 wu0=9.170780164e-09 pu0=-7.358193806e-14
+  ua=-3.606100070e-10 lua=-2.937451054e-15 wua=-3.372823159e-16 pua=2.706191408e-21
+  ub=1.596036216e-18 lub=-4.900486042e-24 wub=-5.626807906e-25 pub=4.514680577e-30
+  uc=5.228259212e-10 luc=-4.770807700e-15 wuc=-5.477909386e-16 puc=4.395211552e-21
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=1.566781148e+06 lvsat=-1.128484939e+01 wvsat=-1.295742488e+00 pvsat=1.039641576e-5
+  a0=-2.457638279e+00 la0=2.976883405e-05 wa0=3.418099946e-06 pa0=-2.742519328e-11
+  ags=2.472130145e+00 lags=-1.790576178e-05 wags=-2.055965084e-06 pags=1.649607697e-11
+  a1=0.0
+  a2=-2.183008898e+00 la2=2.393423155e-05 wa2=2.748162573e-06 pa2=-2.204993737e-11
+  b0=1.577011522e-06 lb0=-1.265318348e-11 wb0=-1.452856559e-12 pb0=1.165702365e-17
+  b1=-5.941276369e-08 lb1=4.766994977e-13 wb1=5.473531563e-14 pb1=-4.391698997e-19
+  keta=-4.446094159e-01 lketa=3.552326954e-06 wketa=4.078832429e-07 pketa=-3.272659357e-12
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=2.351175204e+00 lpclm=-1.773371408e-05 wpclm=-2.036210321e-06 ppclm=1.633757424e-11
+  pdiblc1=0.39
+  pdiblc2=-1.648839157e-02 lpdiblc2=1.348568335e-07 wpdiblc2=1.548445380e-08 ppdiblc2=-1.242398248e-13
+  pdiblcb=1.071080845e+00 lpdiblcb=-9.838443235e-06 wpdiblcb=-1.129664072e-06 ppdiblcb=9.063882276e-12
+  drout=0.56
+  pscbe1=7.990958283e+08 lpscbe1=6.863492872e+00 wpscbe1=7.880760321e-01 ppscbe1=-6.323143805e-6
+  pscbe2=-7.590824359e-08 lpscbe2=6.525826199e-13 wpscbe2=7.493046635e-14 ppscbe2=-6.012060954e-19
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.854711116e-09 lalpha0=-1.407895974e-14 walpha0=-1.616566220e-15 palpha0=1.297055139e-20
+  alpha1=1.854711116e-09 lalpha1=-1.407895974e-14 walpha1=-1.616566220e-15 palpha1=1.297055139e-20
+  beta0=-4.099636412e+02 lbeta0=3.339727861e-03 wbeta0=3.834723122e-04 pbeta0=-3.076797766e-9
* Gidl Induced Drain Leakage Model Parameters
+  agidl=2.402375366e-07 lagidl=-1.822907148e-12 wagidl=-2.093087964e-13 pagidl=1.679393314e-18
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=1.466782197e+01 legidl=-1.105831400e-04 wegidl=-1.269731371e-05 pegidl=1.018771505e-10
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.850165408e-01 lkt1=3.550009698e-07 wkt1=4.076171723e-08 pkt1=-3.270524534e-13
+  kt2=5.621476965e-02 lkt2=-8.711395758e-07 wkt2=-1.000254875e-07 pkt2=8.025564993e-13
+  at=-1.245669422e+06 lat=9.994653517e+00 wat=1.147600359e+00 pat=-9.207794435e-6
+  ute=-9.970951465e-01 lute=6.938972991e-06 wute=7.967427669e-07 pute=-6.392681525e-12
+  ua1=-2.870701542e-09 lua1=3.765779611e-14 wua1=4.323921812e-15 pua1=-3.469307314e-20
+  ub1=8.285974271e-18 lub1=-7.222662903e-23 wub1=-8.293164469e-24 pub1=6.654037098e-29
+  uc1=3.602146143e-10 luc1=-2.960485401e-15 wuc1=-3.399271525e-16 puc1=2.727412306e-21
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.92 pmos
* Model Flag Parameters
+  lmin=4.0e-06 lmax=8.0e-06 wmin=8.6e-07 wmax=9.4e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.090414346e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=1.776925644e-8
+  k1=4.556728822e-01 lk1=-6.543334786e-8
+  k2=1.885398624e-02 lk2=1.709911408e-8
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.057269452e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-5.057204472e-8
+  nfactor={2.150233085e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-2.692133146e-6
+  eta0=0.08
+  etab=-0.07
+  u0=8.535573484e-03 lu0=3.879584672e-9
+  ua=-8.237874492e-10 lua=7.788624164e-16
+  ub=1.048518672e-18 lub=-5.074680762e-25
+  uc=-7.083802061e-11 luc=-7.533189791e-18
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=2.678104074e+05 lvsat=-8.625316685e-1
+  a0=1.347035279e+00 la0=-7.580403376e-7
+  ags=2.084960866e-01 lags=2.565513575e-7
+  a1=0.0
+  a2=0.8
+  b0=0.0
+  b1=0.0
+  keta=-8.364571240e-04 lketa=-8.294256640e-9
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=2.407132755e-01 lpclm=-8.003805848e-7
+  pdiblc1=0.39
+  pdiblc2=-1.397670217e-03 lpdiblc2=1.377612899e-08 ppdiblc2=1.387778781e-29
+  pdiblcb=-2.494013897e-01 lpdiblcb=7.564723865e-7
+  drout=0.56
+  pscbe1=1.227212561e+09 lpscbe1=-3.428139670e+3
+  pscbe2=-1.711599940e-08 lpscbe2=1.808618728e-13 ppscbe2=5.293955920e-35
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=3.429576331e+00 lbeta0=2.285911254e-5
* Gidl Induced Drain Leakage Model Parameters
+  agidl=2.613220901e-08 lagidl=-1.050287696e-13
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=1.675517744e+00 legidl=-6.339127153e-6
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.061103840e-01 lkt1=-2.781041573e-7
+  kt2=-4.839276194e-02 lkt2=-3.181895402e-8
+  at=-9.120917488e+04 lat=7.318186388e-1
+  ute=-1.647219648e-01 lute=2.604101198e-7
+  ua1=5.703275549e-10 lua1=1.004863033e-14
+  ub1=8.239234094e-19 lub1=-1.235471470e-23
+  uc1=-1.164852119e-11 luc1=2.316590399e-17
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.93 pmos
* Model Flag Parameters
+  lmin=2.0e-06 lmax=4.0e-06 wmin=8.6e-07 wmax=9.4e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.085843201e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-6.228379991e-10
+  k1=4.428072554e-01 lk1=-1.366824095e-8
+  k2=2.193345702e-02 lk2=4.708801823e-9
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=8.622137339e-01 ldsub=-1.215963003e-6
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.337857314e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=6.232304277e-8
+  nfactor={7.881674337e-01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=2.788165241e-6
+  eta0=1.604349200e-01 leta0=-3.236315093e-7
+  etab=-1.403185835e-01 letab=2.829282271e-7
+  u0=8.638994592e-03 lu0=3.463467775e-9
+  ua=-8.215637429e-10 lua=7.699152898e-16
+  ub=1.011504174e-18 lub=-3.585395030e-25
+  uc=-7.560382119e-11 luc=1.164210416e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=53438.0
+  a0=1.154071298e+00 la0=1.835409954e-8
+  ags=1.482758150e-01 lags=4.988488244e-7
+  a1=0.0
+  a2=0.8
+  b0=0.0
+  b1=0.0
+  keta=6.578345336e-03 lketa=-3.812786263e-08 wketa=-6.938893904e-24 pketa=1.387778781e-29
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-5.559724103e-01 lpclm=2.405100206e-06 wpclm=-4.440892099e-22 ppclm=-4.440892099e-28
+  pdiblc1=0.39
+  pdiblc2=3.641230659e-03 lpdiblc2=-6.497989463e-9
+  pdiblcb=-9.820554637e-02 lpdiblcb=1.481328872e-7
+  drout=0.56
+  pscbe1=-4.676991234e+07 lpscbe1=1.697754289e+3
+  pscbe2=4.653609693e-08 lpscbe2=-7.524360986e-14
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=1.147359093e+01 lbeta0=-9.506141085e-6
* Gidl Induced Drain Leakage Model Parameters
+  agidl=3.821637237e-11 lagidl=-3.906838872e-17
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.816142056e-01 lkt1=2.568697892e-8
+  kt2=-6.028632264e-02 lkt2=1.603502535e-8
+  at=1.022950518e+05 lat=-4.674948746e-2
+  ute=-1.327375183e-01 lute=1.317200597e-7
+  ua1=3.323674104e-09 lua1=-1.029514575e-15
+  ub1=-2.842323112e-18 lub1=2.396501504e-24
+  uc1=1.818504214e-11 luc1=-9.687003470e-17 puc1=-2.584939414e-38
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.94 pmos
* Model Flag Parameters
+  lmin=1.0e-06 lmax=2.0e-06 wmin=8.6e-07 wmax=9.4e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.101264296e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=3.058205737e-8
+  k1=3.540326720e-01 lk1=1.659689040e-7
+  k2=5.577749960e-02 lk2=-6.377529522e-08 wk2=-5.551115123e-23 pk2=-5.551115123e-29
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=-2.663045674e-01 ldsub=1.067616350e-6
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.021762939e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-1.639286090e-9
+  nfactor={2.430472285e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-5.350714714e-7
+  eta0=-2.241626400e-01 leta0=4.546093453e-07 weta0=-4.857225733e-23 peta0=-9.020562075e-29
+  etab=8.442995791e-01 letab=-1.709466317e-06 wetab=1.994931997e-22 petab=-5.204170428e-29
+  u0=1.250070846e-02 lu0=-4.350787479e-9
+  ua=2.633023699e-11 lua=-9.458151364e-16
+  ub=5.976931819e-19 lub=4.788153150e-25
+  uc=-7.509174596e-11 luc=1.060590969e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=5.963848416e+04 lvsat=-1.254680371e-2
+  a0=1.369865781e+00 la0=-4.183103528e-7
+  ags=1.727992847e-01 lags=4.492250930e-7
+  a1=0.0
+  a2=5.953062352e-01 la2=4.142019269e-7
+  b0=0.0
+  b1=0.0
+  keta=-1.079934288e-02 lketa=-2.963762975e-9
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=4.550220723e-01 lpclm=3.593326501e-7
+  pdiblc1=7.492555200e-01 lpdiblc1=-7.269607298e-7
+  pdiblc2=0.00043
+  pdiblcb=-0.025
+  drout=1.096512000e-01 ldrout=9.112898038e-7
+  pscbe1=7.983183467e+08 lpscbe1=-1.229870506e+1
+  pscbe2=9.530520115e-09 lpscbe2=-3.620850560e-16
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=5.862313582e+00 lbeta0=1.848390856e-6
* Gidl Induced Drain Leakage Model Parameters
+  agidl=2.315918186e-11 lagidl=-8.599862589e-18
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.585366557e-01 lkt1=-2.101090483e-8
+  kt2=-5.625426130e-02 lkt2=7.876068592e-9
+  at=9.703221664e+04 lat=-3.610003518e-2
+  ute=9.359355551e-01 lute=-2.030761278e-06 wute=-4.440892099e-22 pute=-1.110223025e-27
+  ua1=6.136533540e-09 lua1=-6.721391901e-15 pua1=-6.617444900e-36
+  ub1=-4.270929418e-18 lub1=5.287314936e-24
+  uc1=-1.285649500e-10 luc1=2.000815094e-16 puc1=2.067951531e-37
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=2.75e-6
+  sbref=2.74e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.95 pmos
* Model Flag Parameters
+  lmin=5.0e-07 lmax=1.0e-06 wmin=8.6e-07 wmax=9.4e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.092061262e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=2.116256770e-08 wvth0=-4.384852127e-10 pvth0=4.487983849e-16
+  k1=4.471235566e-01 lk1=7.068852186e-08 wk1=6.377510305e-08 pk1=-6.527509347e-14
+  k2=-6.518873286e-02 lk2=6.003606303e-08 wk2=4.909569666e-08 pk2=-5.025042745e-14
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=1.944769162e+00 ldsub=-1.195461833e-06 wdsub=-5.800064896e-07 pdsub=5.936482422e-13
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-5.101041279e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=5.012447003e-06 wvoff=4.515988413e-06 pvoff=-4.622204461e-12
+  nfactor={2.536604250e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-6.436996599e-07 wnfactor=-6.801711405e-07 pnfactor=6.961687658e-13
+  eta0=-4.740445288e-01 leta0=7.103684561e-07 weta0=3.789594597e-07 peta0=-3.878725862e-13
+  etab=-1.690283377e+00 letab=8.847300294e-07 wetab=2.949472572e-10 petab=-3.018844167e-16
+  u0=8.057717978e-03 lu0=1.967021435e-10 wu0=1.692355621e-09 pu0=-1.732159825e-15
+  ua=-1.689296881e-10 lua=-7.459626979e-16 wua=-3.463653728e-16 pua=3.545118864e-22
+  ub=5.972194891e-19 lub=4.793001491e-25 wub=2.436275246e-25 pub=-2.493576440e-31
+  uc=-1.172584348e-10 luc=5.376435909e-17 wuc=1.463162288e-17 puc=-1.497575865e-23
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=5.536765674e+05 lvsat=-5.182046627e-01 wvsat=-5.156617945e-01 pvsat=5.277901599e-7
+  a0=1.556970942e+00 la0=-6.098162269e-07 wa0=-3.128780561e-07 pa0=3.202369480e-13
+  ags=-5.662276679e-02 lags=6.840431512e-07 wags=5.991918073e-16 pags=-6.132836461e-22
+  a1=0.0
+  a2=5.852637642e-01 la2=4.244805969e-07 wa2=3.916255064e-07 pa2=-4.008365384e-13
+  b0=9.657083187e-16 lb0=-9.884217783e-22 wb0=-8.896800342e-22 pb0=9.106053086e-28
+  b1=4.014891572e-19 lb1=-4.109321821e-25 wb1=-3.698807188e-25 pb1=3.785803133e-31
+  keta=6.495412389e-03 lketa=-2.066529089e-08 wketa=4.571931633e-09 pketa=-4.679463465e-15
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=1.966421532e+00 lpclm=-1.187614925e-06 wpclm=-3.182659801e-07 ppclm=3.257515960e-13
+  pdiblc1=1.185765774e-01 lpdiblc1=-8.144821854e-08 wpdiblc1=-4.630290772e-08 ppdiblc1=4.739195211e-14
+  pdiblc2=1.490008763e-03 lpdiblc2=-1.084940169e-09 wpdiblc2=-6.004896790e-10 ppdiblc2=6.146131962e-16
+  pdiblcb=-2.061411941e-01 lpdiblcb=1.854016350e-07 wpdiblcb=1.616030791e-07 ppdiblcb=-1.654039835e-13
+  drout=5.833670991e-01 ldrout=4.264321067e-07 wdrout=3.838322259e-07 pdrout=-3.928599598e-13
+  pscbe1=2.070457412e+08 lpscbe1=5.928806321e+02 wpscbe1=5.204398533e+02 ppscbe1=-5.326805987e-4
+  pscbe2=6.779351986e-08 lpscbe2=-5.999543056e-14 wpscbe2=-5.414801999e-14 ppscbe2=5.542158142e-20
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=6.269740331e+00 lbeta0=1.431381430e-06 wbeta0=2.433852705e-07 pbeta0=-2.491096921e-13
* Gidl Induced Drain Leakage Model Parameters
+  agidl=-1.254542251e-10 lagidl=1.435089317e-16 wagidl=1.309543105e-16 pagidl=-1.340343559e-22
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-3.710212029e-01 lkt1=-1.105847211e-07 wkt1=-4.262050217e-08 pkt1=4.362293639e-14
+  kt2=-8.814795627e-02 lkt2=4.051990327e-08 wkt2=2.114036593e-08 pkt2=-2.163758734e-14
+  at=1.280264439e+05 lat=-6.782324670e-02 wat=-3.532098456e-02 pat=3.615173412e-8
+  ute=-1.971926414e+00 lute=9.454936047e-07 wute=3.149936657e-08 pute=-3.224023167e-14
+  ua1=-4.337391766e-09 lua1=3.998880129e-15 wua1=7.085589762e-16 pua1=-7.252242833e-22
+  ub1=5.727350586e-18 lub1=-4.946124613e-24 wub1=-1.236505782e-24 pub1=1.265588398e-30
+  uc1=4.507626996e-10 luc1=-3.928719265e-16 wuc1=-1.006572140e-16 puc1=1.030246717e-22
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.75e-6
+  sbref=1.74e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.96 pmos
* Model Flag Parameters
+  lmin=2.5e-07 lmax=5.0e-07 wmin=8.6e-07 wmax=9.4e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.109173714e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=3.012127881e-08 wvth0=5.323678299e-08 pvth0=-2.765127802e-14
+  k1=1.109811951e+00 lk1=-2.762421066e-07 wk1=-5.675141823e-07 pk1=2.652174732e-13
+  k2=-1.605798384e-01 lk2=1.099752146e-07 wk2=1.469443066e-07 pk2=-1.014761317e-13
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=-1.939047575e+00 ldsub=8.377939055e-07 wdsub=1.472374995e-06 pdsub=-4.808145127e-13
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={8.123588622e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-1.910911242e-06 wvoff=-7.554661423e-06 pvoff=1.697022141e-12
+  nfactor={-4.930806507e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=3.265639219e-06 wnfactor=5.586797182e-06 pnfactor=-2.584714491e-12
+  eta0=1.312687464e+00 leta0=-2.250214766e-07 weta0=-7.579189251e-07 peta0=2.073059858e-13
+  etab=-1.415877886e-03 letab=5.741164906e-10 wetab=1.049475160e-10 petab=-2.024157522e-16
+  u0=6.564068158e-03 lu0=9.786576973e-10 wu0=7.749273201e-10 pu0=-1.251867761e-15
+  ua=-2.996744630e-09 lua=7.344549806e-16 wua=1.626450919e-15 pua=-6.782968990e-22
+  ub=2.503952912e-18 lub=-5.189129324e-25 wub=-1.140657496e-24 pub=4.753432499e-31
+  uc=-4.247910009e-11 luc=1.461588176e-17 wuc=-1.826705235e-17 puc=2.247355810e-24
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=-3.848712483e+05 lvsat=-2.685611021e-02 wvsat=4.437138804e-01 pvsat=2.553780658e-8
+  a0=4.256318575e-01 la0=-1.753758954e-08 wa0=3.923298295e-07 pa0=-4.895348425e-14
+  ags=6.986456739e-01 lags=2.886450171e-07 wags=2.281416958e-07 pags=-1.194367409e-13
+  a1=0.0
+  a2=2.002479027e+00 la2=-3.174599373e-07 wa2=-7.410857714e-07 pa2=1.921604698e-13
+  b0=-1.931416637e-15 lb0=5.282810787e-22 wb0=1.779360068e-21 pb0=-4.866905659e-28
+  b1=-8.029783143e-19 lb1=2.196306285e-25 wb1=7.397614376e-25 pb1=-2.023395484e-31
+  keta=-1.409751721e-02 lketa=-9.884480386e-09 wketa=-2.620189628e-08 pketa=1.143125093e-14
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-1.347163432e+00 lpclm=5.471130757e-07 wpclm=6.511689539e-07 ppclm=-1.817669807e-13
+  pdiblc1=-5.726628509e-01 lpdiblc1=2.804294470e-07 wpdiblc1=1.367569853e-07 ppdiblc1=-4.844356308e-14
+  pdiblc2=-1.837542311e-02 lpdiblc2=9.315010725e-09 wpdiblc2=7.739740690e-09 ppdiblc2=-3.751664206e-15
+  pdiblcb=-2.762138169e-01 lpdiblcb=2.220860544e-07 wpdiblcb=4.349994561e-07 ppdiblcb=-3.085324548e-13
+  drout=2.848056641e+00 ldrout=-7.591781623e-07 wdrout=-1.187568846e-06 pdrout=4.297999291e-13
+  pscbe1=1.929886384e+09 lpscbe1=-3.090609010e+02 wpscbe1=-1.040903508e+03 ppscbe1=2.847138781e-4
+  pscbe2=-1.116014043e-07 lpscbe2=3.392140013e-14 wpscbe2=1.115836522e-13 ppscbe2=-3.134226358e-20
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=8.517860617e+00 lbeta0=2.544454975e-07 wbeta0=8.577889655e-09 pbeta0=-1.261833320e-13
* Gidl Induced Drain Leakage Model Parameters
+  agidl=-7.502812130e-10 lagidl=4.706183564e-16 wagidl=6.311905766e-16 pagidl=-3.959180459e-22
+  bgidl=4.828711902e+08 lbgidl=2.707272745e+02 wbgidl=2.139796996e+02 pbgidl=-1.120226523e-4
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.00074326333
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.5407449e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-7.150100359e-01 lkt1=6.950031279e-08 wkt1=1.421813972e-07 pkt1=-5.312455396e-14
+  kt2=3.741936112e-02 lkt2=-2.521709874e-08 wkt2=-4.408674899e-08 pkt2=1.251011186e-14
+  at=-1.300048782e+05 lat=6.726131105e-02 wat=1.148381402e-01 pat=-4.245957086e-8
+  ute=9.377795349e-01 lute=-5.777956537e-07 wute=-3.760109742e-07 pute=1.810995819e-13
+  ua1=6.648068028e-09 lua1=-1.752227783e-15 wua1=-1.466068265e-15 pua1=4.132365700e-22
+  ub1=-7.546993544e-18 lub1=2.003260026e-24 wub1=2.423609229e-24 pub1=-6.505550122e-31
+  uc1=-4.478273428e-10 luc1=7.755793247e-17 wuc1=1.402110959e-16 puc1=-2.307470589e-23
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.1e-6
+  sbref=1.1e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.97 pmos
* Model Flag Parameters
+  lmin=1.8e-07 lmax=2.5e-07 wmin=8.6e-07 wmax=9.4e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.056751455e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=1.578274251e-08 wvth0=3.163427332e-08 pvth0=-2.174255958e-14
+  k1=2.740141511e+00 lk1=-7.221698477e-07 wk1=-3.122384660e-06 pk1=9.640256464e-13
+  k2=-9.232216845e-01 lk2=3.185730123e-07 wk2=1.236229036e-06 pk2=-3.994172909e-13
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=-1.961943366e+01 ldsub=5.673733106e-06 wdsub=1.832676099e-05 pdsub=-5.090826170e-12
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={7.254636573e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-1.673235478e-06 wvoff=-6.860950608e-06 pvoff=1.507278359e-12
+  nfactor={1.544191267e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-2.306706931e-06 wnfactor=-1.101939616e-05 pnfactor=1.957411513e-12
+  eta0=-5.025852912e+00 leta0=1.508696087e-06 weta0=5.302005046e-06 peta0=-1.450204419e-12
+  etab=-8.338919171e-01 letab=2.282729627e-07 wetab=7.682355163e-07 petab=-2.103014889e-13
+  u0=4.357750687e-02 lu0=-9.145258059e-09 wu0=-2.506872134e-08 pu0=5.816887020e-15
+  ua=9.954991835e-09 lua=-2.808103977e-15 wua=-7.014146939e-15 pua=1.685079427e-21
+  ub=-7.378858977e-18 lub=2.184233775e-24 wub=5.539153510e-24 pub=-1.351718657e-30
+  uc=3.745742757e-10 luc=-9.945655758e-17 wuc=-3.185824807e-16 puc=8.438963176e-23
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=-4.854511133e+06 lvsat=1.195679791e+00 wvsat=4.395875889e+00 pvsat=-1.055457546e-6
+  a0=5.406891204e+00 la0=-1.380011646e-06 wa0=-5.298611007e-06 pa0=1.507632653e-12
+  ags=3.219122860e+00 lags=-4.007559028e-07 wags=-8.147920164e-07 pags=1.658264881e-13
+  a1=0.0
+  a2=3.947369826e+00 la2=-8.494264687e-07 wa2=-2.282255605e-06 pa2=6.137012426e-13
+  b0=0.0
+  b1=0.0
+  keta=1.531559476e+00 lketa=-4.326525812e-07 wketa=-1.394564923e-06 pketa=3.857059059e-13
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-1.317697242e+00 lpclm=5.390534834e-07 wpclm=1.681594483e-06 ppclm=-4.636089714e-13
+  pdiblc1=-6.438863031e+00 lpdiblc1=1.884952520e-06 wpdiblc1=6.336680243e-06 ppdiblc1=-1.744246572e-12
+  pdiblc2=-1.534895234e-01 lpdiblc2=4.627141944e-08 wpdiblc2=1.478802272e-07 ppdiblc2=-4.208289008e-14
+  pdiblcb=-5.040604436e+00 lpdiblcb=1.525242177e-06 wpdiblcb=4.222430023e-06 ppdiblcb=-1.344470463e-12
+  drout=1.446588620e+01 ldrout=-3.936886904e-06 wdrout=-1.287779742e-05 pdrout=3.627311248e-12
+  pscbe1=7.997946110e+08 lpscbe1=4.180064201e-02 wpscbe1=8.500476963e-02 ppscbe1=-1.730005833e-8
+  pscbe2=5.121817788e-08 lpscbe2=-1.061301198e-14 wpscbe2=-3.206061204e-14 ppscbe2=7.947315563e-21
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=-1.765866458e+01 lbeta0=7.414248670e-06 wbeta0=2.371745873e-05 pbeta0=-6.611036421e-12
* Gidl Induced Drain Leakage Model Parameters
+  agidl=1.080202923e-08 lagidl=-2.689169595e-15 wagidl=-9.648291139e-15 pagidl=2.415725793e-21
+  bgidl=2.846889940e+09 lbgidl=-3.758791340e+02 wbgidl=-7.642144419e+02 pbgidl=1.555330093e-4
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.00074326333
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.5407449e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-1.094728920e+01 lkt1=2.868233310e-06 wkt1=9.539836508e-06 pkt1=-2.623571180e-12
+  kt2=-1.717196849e+00 lkt2=4.547055269e-07 wkt2=1.506465157e-06 pkt2=-4.115968454e-13
+  at=5.611303158e+02 lat=3.154889641e-02 wat=1.217720985e-01 pat=-4.435614715e-8
+  ute=2.174776622e+00 lute=-9.161390968e-07 wute=-4.450749522e-06 pute=1.295622069e-12
+  ua1=1.716354095e-08 lua1=-4.628419937e-15 wua1=-1.528811085e-14 pua1=4.193841657e-21
+  ub1=-2.765469405e-17 lub1=7.503118269e-24 wub1=2.386447525e-23 pub1=-6.515060686e-30
+  uc1=-1.356702599e-10 luc1=-7.823272837e-18 wuc1=-1.539748820e-16 puc1=5.739104277e-23
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.1e-6
+  sbref=1.1e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.98 pmos
* Model Flag Parameters
+  lmin=1.5e-07 lmax=1.8e-07 wmin=8.6e-07 wmax=9.4e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-2.026e-8
+  vth0={-3.264087566e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-1.439540989e-07 wvth0=-6.233917829e-07 pvth0=1.208876331e-13
+  k1=-1.172147688e+01 lk1=2.406583484e-06 wk1=1.082083412e-05 pk1=-2.030208019e-12
+  k2=5.875207988e+00 lk2=-1.154006335e-06 wk2=-5.068592599e-06 pk2=9.575586999e-13
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=5.901908945e+01 ldsub=-1.119370780e-05 wdsub=-4.938492031e-05 pdsub=9.415717721e-12
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-3.662014214e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=5.943392047e-07 wvoff=2.485118580e-06 pvoff=-4.278140462e-13
+  nfactor={4.187705455e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-8.328863356e-06 wnfactor=-4.045289874e-05 pnfactor=8.611589838e-12
+  eta0=1.683846524e+01 leta0=-3.186802158e-06 weta0=-1.396738356e-05 peta0=2.677945764e-12
+  etab=1.673525447e+00 letab=-3.055951025e-07 wetab=-1.443220823e-06 petab=2.598024062e-13
+  u0=-5.302491152e-02 lu0=1.139360499e-08 wu0=4.763169534e-08 pu0=-9.729125024e-15
+  ua=-2.573106509e-08 lua=4.826824724e-15 wua=1.943290518e-14 pua=-4.006270034e-21
+  ub=2.369183097e-17 lub=-4.485025999e-24 wub=-1.797237258e-23 pub=3.720134187e-30
+  uc=-8.366050051e-10 luc=1.593251037e-16 wuc=7.039387410e-16 puc=-1.340476927e-22
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=5.907639769e+06 lvsat=-1.077714743e+00 wvsat=-5.183648347e+00 pvsat=9.688569025e-7
+  a0=-8.863828386e+00 la0=1.651695239e-06 wa0=8.578942522e-06 pa0=-1.426713085e-12
+  ags=1.249999336e+00 lags=1.266467891e-13 wags=6.102395105e-13 pags=-1.162628287e-19
+  a1=0.0
+  a2=-1.204343407e+01 la2=2.605913121e-06 wa2=1.054894922e-05 pa2=-2.164573657e-12
+  b0=0.0
+  b1=0.0
+  keta=-4.322831259e+00 lketa=8.222182479e-07 wketa=3.638338315e-06 pketa=-6.919319502e-13
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=5.826944007e+00 lpclm=-9.914557353e-07 wpclm=-4.378826086e-06 ppclm=8.341097733e-13
+  pdiblc1=2.025411758e+01 lpdiblc1=-3.843933717e-06 wpdiblc1=-1.688673174e-05 ppdiblc1=3.231283541e-12
+  pdiblc2=5.583653931e-01 lpdiblc2=-1.068417809e-07 wpdiblc2=-4.656925133e-07 ppdiblc2=8.970699215e-14
+  pdiblcb=1.880451558e+01 lpdiblcb=-3.605680402e-06 wpdiblcb=-1.617199622e-05 ppdiblcb=3.040604963e-12
+  drout=-4.220791155e+01 ldrout=8.231971310e-06 wdrout=3.634960716e-05 pdrout=-6.925327158e-12
+  pscbe1=7.999999959e+08 lpscbe1=7.700996399e-07 wpscbe1=4.058937073e-06 ppscbe1=-7.733097076e-13
+  pscbe2=-9.105638215e-08 lpscbe2=1.987487044e-14 wpscbe2=8.206285526e-14 ppscbe2=-1.655535318e-20
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=8.969667289e+01 lbeta0=-1.564043909e-05 wbeta0=-6.833842214e-05 pbeta0=1.313690739e-11
* Gidl Induced Drain Leakage Model Parameters
+  agidl=-1.772440360e-08 lagidl=3.376853374e-15 wagidl=1.632899675e-14 pagidl=-3.111000461e-21
+  bgidl=9.999966275e+08 lbgidl=6.425194740e-04 wbgidl=3.107183899e-03 pbgidl=-5.919806728e-10
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-1.106e-8
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=2.769813041e+01 lkt1=-5.414271456e-06 wkt1=-2.559271509e-05 pkt1=4.904712529e-12
+  kt2=4.411667933e+00 lkt2=-8.588502391e-07 wkt2=-3.792392723e-06 pkt2=7.225266615e-13
+  at=1.621593020e+06 lat=-3.232857805e-01 wat=-1.314690393e+00 pat=2.687074981e-7
+  ute=-1.853788579e+01 lute=3.574892236e-06 wute=1.551828691e-05 pute=-2.999726696e-12
+  ua1=-4.572646945e-08 lua1=8.853473822e-15 wua1=3.909395067e-14 pua1=-7.448179483e-21
+  ub1=7.071598043e-17 lub1=-1.356284834e-23 wub1=-5.988896015e-23 pub1=1.141004469e-29
+  uc1=-1.140497910e-09 luc1=2.131078435e-16 wuc1=9.410122790e-16 puc1=-1.792816594e-22
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.04e-6
+  sbref=1.04e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.99 pmos
* Model Flag Parameters
+  lmin=2.0e-05 lmax=0.0001 wmin=8.4e-07 wmax=8.6e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.126311+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+  k1=0.43165561
+  k2=0.026980026
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=3.2465718e-7
+  voff={-0.23051772+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.8768912+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+  eta0=0.08
+  etab=-0.07
+  u0=0.0095864
+  ua=-7.4757916e-10
+  ub=9.5046395e-19
+  uc=-1.0566299e-10
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=80156.0
+  a0=1.464
+  ags=0.11329
+  a1=0.0
+  a2=0.97
+  b0=-8.9873e-8
+  b1=3.3859e-9
+  keta=0.023361259
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=0.015
+  pdiblc1=0.39
+  pdiblc2=0.0012771588
+  pdiblcb=-0.225
+  drout=0.56
+  pscbe1=800000000.0
+  pscbe2=1.0060625e-8
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=0.0
+  alpha1=0.0
+  beta0=30.0
* Gidl Induced Drain Leakage Model Parameters
+  agidl=9.43573999999999e-11
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-0.43825
+  kt2=-0.058546
+  at=70990.0
+  ute=-0.08298
+  ua1=2.0902e-9
+  ub1=-1.2289e-18
+  uc1=-2.9789e-11
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.100 pmos
* Model Flag Parameters
+  lmin=8.0e-06 lmax=2.0e-05 wmin=8.4e-07 wmax=8.6e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.151793231e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=5.102439717e-7
+  k1=4.210498003e-01 lk1=2.123656422e-7
+  k2=3.098838670e-02 lk2=-8.026149068e-8
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=-6.144535039e-06 lcit=1.295359998e-10 wcit=3.388131789e-27 pcit=-5.421010862e-32
+  voff={-2.428791561e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=2.475194627e-7
+  nfactor={1.918471956e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-8.325930941e-7
+  eta0=0.08
+  etab=-0.07
+  u0=9.965711908e-03 lu0=-7.595159576e-9
+  ua=-7.615294670e-10 lua=2.793342514e-16
+  ub=9.271909546e-19 lub=4.660072882e-25 wub=6.162975822e-39
+  uc=-1.283201274e-10 luc=4.536756436e-16
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=2.656289816e+04 lvsat=1.073122547e+0
+  a0=1.605375760e+00 la0=-2.830840351e-6
+  ags=2.825339191e-02 lags=1.702732223e-6
+  a1=0.0
+  a2=1.083666533e+00 la2=-2.276004104e-6
+  b0=-1.499644844e-07 lb0=1.203243040e-12
+  b1=5.649803031e-09 lb1=-4.533130761e-14
+  keta=4.023168533e-02 lketa=-3.378053190e-7
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-6.921953293e-02 lpclm=1.686371502e-06 ppclm=1.776356839e-27
+  pdiblc1=0.39
+  pdiblc2=1.917610060e-03 lpdiblc2=-1.282408862e-8
+  pdiblcb=-2.717239457e-01 lpdiblcb=9.355778616e-07 wpdiblcb=-1.776356839e-21
+  drout=0.56
+  pscbe1=8.000325956e+08 lpscbe1=-6.526776473e-1
+  pscbe2=1.315981805e-08 lpscbe2=-6.205675405e-14
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=-6.686266667e-11 lalpha0=1.338825943e-15
+  alpha1=-6.686266667e-11 lalpha1=1.338825943e-15
+  beta0=4.586076776e+01 lbeta0=-3.175884006e-4
* Gidl Induced Drain Leakage Model Parameters
+  agidl=-8.562847058e-09 lagidl=1.733477066e-13 wagidl=2.481541838e-29 pagidl=-3.705769144e-34
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=-4.251725813e-01 legidl=1.051580369e-05 pegidl=-1.421085472e-26
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.365640579e-01 lkt1=-3.375849616e-8
+  kt2=-6.268314622e-02 lkt2=8.284023011e-8
+  at=1.184558071e+05 lat=-9.504325371e-1
+  ute=-5.002598587e-02 lute=-6.598553610e-7
+  ua1=2.269041386e-09 lua1=-3.581034063e-15
+  ub1=-1.571912915e-18 lub1=6.868325966e-24
+  uc1=-4.384869988e-11 luc1=2.815246818e-16
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.101 pmos
* Model Flag Parameters
+  lmin=4.0e-06 lmax=8.0e-06 wmin=8.4e-07 wmax=8.6e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.090414346e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=1.776925644e-8
+  k1=4.556728822e-01 lk1=-6.543334786e-8
+  k2=1.885398624e-02 lk2=1.709911408e-8
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.057269452e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-5.057204472e-8
+  nfactor={2.150233085e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-2.692133146e-06 wnfactor=1.421085472e-20
+  eta0=0.08
+  etab=-0.07
+  u0=8.535573484e-03 lu0=3.879584672e-9
+  ua=-8.237874492e-10 lua=7.788624164e-16
+  ub=1.048518672e-18 lub=-5.074680762e-25
+  uc=-7.083802061e-11 luc=-7.533189791e-18
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=2.678104074e+05 lvsat=-8.625316685e-1
+  a0=1.347035279e+00 la0=-7.580403376e-7
+  ags=2.084960866e-01 lags=2.565513575e-7
+  a1=0.0
+  a2=0.8
+  b0=0.0
+  b1=0.0
+  keta=-8.364571240e-04 lketa=-8.294256640e-9
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=2.407132755e-01 lpclm=-8.003805848e-7
+  pdiblc1=0.39
+  pdiblc2=-1.397670217e-03 lpdiblc2=1.377612899e-08 wpdiblc2=-3.469446952e-24 ppdiblc2=2.775557562e-29
+  pdiblcb=-2.494013897e-01 lpdiblcb=7.564723865e-07 wpdiblcb=1.776356839e-21
+  drout=0.56
+  pscbe1=1.227212561e+09 lpscbe1=-3.428139670e+3
+  pscbe2=-1.711599940e-08 lpscbe2=1.808618728e-13 wpscbe2=5.293955920e-29 ppscbe2=-4.235164736e-34
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=3.429576331e+00 lbeta0=2.285911254e-5
* Gidl Induced Drain Leakage Model Parameters
+  agidl=2.613220901e-08 lagidl=-1.050287696e-13
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=1.675517744e+00 legidl=-6.339127153e-6
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.061103840e-01 lkt1=-2.781041573e-7
+  kt2=-4.839276194e-02 lkt2=-3.181895402e-8
+  at=-9.120917488e+04 lat=7.318186388e-1
+  ute=-1.647219648e-01 lute=2.604101198e-7
+  ua1=5.703275549e-10 lua1=1.004863033e-14
+  ub1=8.239234094e-19 lub1=-1.235471470e-23 pub1=2.465190329e-44
+  uc1=-1.164852119e-11 luc1=2.316590399e-17
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.102 pmos
* Model Flag Parameters
+  lmin=2.0e-06 lmax=4.0e-06 wmin=8.4e-07 wmax=8.6e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.085843201e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-6.228379991e-10
+  k1=4.428072554e-01 lk1=-1.366824095e-8
+  k2=2.193345702e-02 lk2=4.708801823e-9
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=8.622137339e-01 ldsub=-1.215963003e-6
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.337857314e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=6.232304277e-8
+  nfactor={7.881674337e-01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=2.788165241e-6
+  eta0=1.604349200e-01 leta0=-3.236315093e-7
+  etab=-1.403185835e-01 letab=2.829282271e-7
+  u0=8.638994592e-03 lu0=3.463467775e-9
+  ua=-8.215637429e-10 lua=7.699152898e-16
+  ub=1.011504174e-18 lub=-3.585395030e-25
+  uc=-7.560382119e-11 luc=1.164210416e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=53438.0
+  a0=1.154071298e+00 la0=1.835409954e-8
+  ags=1.482758150e-01 lags=4.988488244e-7
+  a1=0.0
+  a2=0.8
+  b0=0.0
+  b1=0.0
+  keta=6.578345336e-03 lketa=-3.812786263e-08 pketa=-5.551115123e-29
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-5.559724103e-01 lpclm=2.405100206e-06 wpclm=4.440892099e-22 ppclm=-8.881784197e-28
+  pdiblc1=0.39
+  pdiblc2=3.641230659e-03 lpdiblc2=-6.497989463e-9
+  pdiblcb=-9.820554637e-02 lpdiblcb=1.481328872e-7
+  drout=0.56
+  pscbe1=-4.676991234e+07 lpscbe1=1.697754289e+3
+  pscbe2=4.653609693e-08 lpscbe2=-7.524360986e-14
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=1.147359093e+01 lbeta0=-9.506141085e-6
* Gidl Induced Drain Leakage Model Parameters
+  agidl=3.821637237e-11 lagidl=-3.906838872e-17
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.816142056e-01 lkt1=2.568697892e-8
+  kt2=-6.028632264e-02 lkt2=1.603502535e-8
+  at=1.022950518e+05 lat=-4.674948746e-2
+  ute=-1.327375183e-01 lute=1.317200597e-07 wute=-8.881784197e-22
+  ua1=3.323674104e-09 lua1=-1.029514575e-15
+  ub1=-2.842323112e-18 lub1=2.396501504e-24
+  uc1=1.818504214e-11 luc1=-9.687003470e-17
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.103 pmos
* Model Flag Parameters
+  lmin=1.0e-06 lmax=2.0e-06 wmin=8.4e-07 wmax=8.6e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.101264296e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=3.058205737e-8
+  k1=3.540326720e-01 lk1=1.659689040e-7
+  k2=5.577749960e-02 lk2=-6.377529522e-8
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=-2.663045674e-01 ldsub=1.067616350e-6
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.021762939e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-1.639286090e-9
+  nfactor={2.430472285e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-5.350714714e-7
+  eta0=-2.241626400e-01 leta0=4.546093453e-07 weta0=-1.387778781e-22 peta0=2.220446049e-28
+  etab=8.442995791e-01 letab=-1.709466317e-06 wetab=1.498801083e-21 petab=9.298117831e-28
+  u0=1.250070846e-02 lu0=-4.350787479e-9
+  ua=2.633023699e-11 lua=-9.458151364e-16
+  ub=5.976931819e-19 lub=4.788153150e-25
+  uc=-7.509174596e-11 luc=1.060590969e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=5.963848416e+04 lvsat=-1.254680371e-2
+  a0=1.369865781e+00 la0=-4.183103528e-7
+  ags=1.727992847e-01 lags=4.492250930e-7
+  a1=0.0
+  a2=5.953062352e-01 la2=4.142019269e-7
+  b0=0.0
+  b1=0.0
+  keta=-1.079934288e-02 lketa=-2.963762975e-9
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=4.550220723e-01 lpclm=3.593326501e-7
+  pdiblc1=7.492555200e-01 lpdiblc1=-7.269607298e-7
+  pdiblc2=0.00043
+  pdiblcb=-0.025
+  drout=1.096512000e-01 ldrout=9.112898038e-7
+  pscbe1=7.983183467e+08 lpscbe1=-1.229870506e+1
+  pscbe2=9.530520115e-09 lpscbe2=-3.620850560e-16
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=5.862313582e+00 lbeta0=1.848390856e-6
* Gidl Induced Drain Leakage Model Parameters
+  agidl=2.315918186e-11 lagidl=-8.599862589e-18
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.585366557e-01 lkt1=-2.101090483e-8
+  kt2=-5.625426130e-02 lkt2=7.876068592e-9
+  at=9.703221664e+04 lat=-3.610003518e-2
+  ute=9.359355551e-01 lute=-2.030761278e-06 wute=-3.552713679e-21 pute=-8.881784197e-28
+  ua1=6.136533540e-09 lua1=-6.721391901e-15
+  ub1=-4.270929418e-18 lub1=5.287314936e-24
+  uc1=-1.285649500e-10 luc1=2.000815094e-16 wuc1=4.135903063e-31 puc1=-4.135903063e-37
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=2.75e-6
+  sbref=2.74e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.104 pmos
* Model Flag Parameters
+  lmin=5.0e-07 lmax=1.0e-06 wmin=8.4e-07 wmax=8.6e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.092582479e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=2.169604366e-8
+  k1=5.229315034e-01 lk1=-6.902427879e-9
+  k2=-6.829846957e-03 lk2=3.045761312e-10
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=1.255329254e+00 ldsub=-4.898062988e-07 wdsub=-7.105427358e-21 pdsub=-3.552713679e-27
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={2.670066454e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-4.818574081e-7
+  nfactor={1.728101006e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.838195797e-7
+  eta0=-2.358444013e-02 leta0=2.493135462e-7
+  etab=-1.689932780e+00 letab=8.843711865e-7
+  u0=1.006938082e-02 lu0=-1.862275006e-9
+  ua=-5.806459616e-10 lua=-3.245628577e-16
+  ub=8.868137281e-19 lub=1.828946535e-25
+  uc=-9.986617302e-11 luc=3.596303128e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=-5.927833243e+04 lvsat=1.091669364e-1
+  a0=1.185060244e+00 la0=-2.291581900e-7
+  ags=-5.662276608e-02 lags=6.840431505e-7
+  a1=0.0
+  a2=1.050779681e+00 la2=-5.198425436e-8
+  b0=-9.183315919e-17 lb0=9.399307509e-23
+  b1=-3.817924830e-20 lb1=3.907722422e-26
+  keta=1.192995869e-02 lketa=-2.622765772e-8
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=1.588106337e+00 lpclm=-8.004017569e-7
+  pdiblc1=6.353741327e-02 lpdiblc1=-2.511453323e-8
+  pdiblc2=7.762209763e-04 lpdiblc2=-3.543640937e-10
+  pdiblcb=-1.404746093e-02 lpdiblcb=-1.121014279e-8
+  drout=1.039619329e+00 ldrout=-4.055117553e-8
+  pscbe1=8.256802058e+08 lpscbe1=-4.030411509e+1
+  pscbe2=3.429057487e-09 lpscbe2=5.882883972e-15
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=6.559046608e+00 lbeta0=1.135270669e-6
* Gidl Induced Drain Leakage Model Parameters
+  agidl=3.020804646e-11 lagidl=-1.581451648e-17
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.216831793e-01 lkt1=-5.873117501e-8
+  kt2=-6.301890653e-02 lkt2=1.479981827e-8
+  at=8.604123040e+04 lat=-2.485054094e-2
+  ute=-1.934483867e+00 lute=9.071704088e-7
+  ua1=-3.495144579e-09 lua1=3.136823287e-15 pua1=6.617444900e-36
+  ub1=4.257545597e-18 lub1=-3.441749811e-24 wub1=1.232595164e-38
+  uc1=3.311138654e-10 luc1=-2.704089518e-16 wuc1=-8.271806126e-31 puc1=4.135903063e-37
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.75e-6
+  sbref=1.74e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.105 pmos
* Model Flag Parameters
+  lmin=2.5e-07 lmax=5.0e-07 wmin=8.4e-07 wmax=8.6e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.045892418e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-2.747137143e-9
+  k1=4.352213524e-01 lk1=3.901559036e-8
+  k2=1.408936088e-02 lk2=-1.064704755e-08 pk2=-1.387778781e-29
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=-1.888704683e-01 ldsub=2.662611400e-7
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-8.564575735e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=1.062985797e-7
+  nfactor={1.710086311e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.932506331e-7
+  eta0=4.117672797e-01 leta0=2.139821381e-8
+  etab=-1.291129272e-03 letab=3.335097045e-10
+  u0=7.485205816e-03 lu0=-5.094077095e-10 wu0=-5.551115123e-23
+  ua=-1.063421140e-09 lua=-7.182039643e-17
+  ub=1.148080500e-18 lub=4.611627323e-26
+  uc=-6.419271038e-11 luc=1.728726011e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=1.425608788e+05 lvsat=3.500072552e-3
+  a0=8.919849864e-01 la0=-7.572743094e-8
+  ags=9.698322768e-01 lags=1.466734064e-7
+  a1=0.0
+  a2=1.121568012e+00 la2=-8.904336116e-8
+  b0=1.836663184e-16 lb0=-5.023641140e-23
+  b1=7.635849659e-20 lb1=-2.088557599e-26
+  keta=-4.524308758e-02 lketa=3.703575468e-9
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-5.731343976e-01 lpclm=3.310509927e-07 wpclm=8.881784197e-22 ppclm=-6.661338148e-28
+  pdiblc1=-4.101030779e-01 lpdiblc1=2.228457367e-07 wpdiblc1=-6.661338148e-22 ppdiblc1=-3.885780586e-28
+  pdiblc2=-9.175377595e-03 lpdiblc2=4.855496791e-09 wpdiblc2=-1.734723476e-24 ppdiblc2=-5.637851297e-30
+  pdiblcb=2.408596814e-01 lpdiblcb=-1.446591300e-07 wpdiblcb=4.440892099e-22 ppdiblcb=2.220446049e-28
+  drout=1.436421824e+00 ldrout=-2.482852179e-7
+  pscbe1=6.925891618e+08 lpscbe1=2.937170827e+1
+  pscbe2=2.103542680e-08 lpscbe2=-3.334402489e-15
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=8.528056950e+00 lbeta0=1.044543745e-7
* Gidl Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=7.372237654e+08 lbgidl=1.375686143e+2
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.00074326333
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.5407449e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-5.460023937e-01 lkt1=6.352420121e-9
+  kt2=-1.498550792e-02 lkt2=-1.034662657e-8
+  at=6.500485322e+03 lat=1.679062992e-2
+  ute=4.908242408e-01 lute=-3.625268917e-07 pute=8.881784197e-28
+  ua1=4.905387581e-09 lua1=-1.261023309e-15
+  ub1=-4.666106948e-18 lub1=1.229960769e-24
+  uc1=-2.811617509e-10 luc1=5.012957887e-17
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.1e-6
+  sbref=1.1e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.106 pmos
* Model Flag Parameters
+  lmin=1.8e-07 lmax=2.5e-07 wmin=8.4e-07 wmax=8.6e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.019148548e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-1.006212048e-8
+  k1=-9.713628067e-01 lk1=4.237444896e-7
+  k2=5.462543423e-01 lk2=-1.562048133e-07 wk2=4.440892099e-22 pk2=3.330669074e-28
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=2.165150868e+00 ldsub=-3.776107759e-7
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-9.008120908e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=1.184304273e-7
+  nfactor={2.343418770e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=2.002153880e-8
+  eta0=1.276514272e+00 leta0=-2.151273835e-7
+  etab=7.929135335e-02 letab=-2.170741094e-08 wetab=-6.245004514e-23 petab=9.107298249e-30
+  u0=1.377891457e-02 lu0=-2.230862929e-9
+  ua=1.617442340e-09 lua=-8.050901755e-16
+  ub=-7.945990585e-19 lub=5.774779860e-25
+  uc=-4.117135234e-12 luc=8.553888012e-19
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=3.707618922e+05 lvsat=-5.891746863e-2
+  a0=-8.914415674e-01 la0=4.120754001e-7
+  ags=2.250598986e+00 lags=-2.036419039e-7
+  a1=0.0
+  a2=1.234506918e+00 la2=-1.199344107e-7
+  b0=0.0
+  b1=0.0
+  keta=-1.261266502e-01 lketa=2.582684751e-8
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=6.811740897e-01 lpclm=-1.202746476e-8
+  pdiblc1=1.093397930e+00 lpdiblc1=-1.883918589e-7
+  pdiblc2=2.229218241e-02 lpdiblc2=-3.751510221e-09 ppdiblc2=2.775557562e-29
+  pdiblcb=-2.150238278e-02 lpdiblcb=-7.289785815e-8
+  drout=-8.416450324e-01 ldrout=3.748116287e-7
+  pscbe1=7.998956542e+08 lpscbe1=2.123647450e-2
+  pscbe2=1.310849154e-08 lpscbe2=-1.166227157e-15
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=1.053371402e+01 lbeta0=-4.441329485e-7
* Gidl Induced Drain Leakage Model Parameters
+  agidl=-6.666647741e-10 lagidl=1.823461490e-16
+  bgidl=1.938486425e+09 lbgidl=-1.910007484e+2
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.00074326333
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.5407449e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=3.924873623e-01 lkt1=-2.503432980e-7
+  kt2=7.350242203e-02 lkt2=-3.454984517e-8
+  at=1.453087251e+05 lat=-2.117619981e-2
+  ute=-3.115723385e+00 lute=6.239360150e-7
+  ua1=-1.009072480e-09 lua1=3.566998069e-16
+  ub1=7.124395827e-19 lub1=-2.411792780e-25 pub1=-7.703719778e-46
+  uc1=-3.186965368e-10 luc1=6.039609351e-17
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.1e-6
+  sbref=1.1e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.107 pmos
* Model Flag Parameters
+  lmin=1.5e-07 lmax=1.8e-07 wmin=8.4e-07 wmax=8.6e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-2.026e-8
+  vth0={-1.019405789e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-1.084588123e-08 wvth0=-4.039278319e-08 pvth0=8.907416548e-15
+  k1=2.384239477e+00 lk1=-2.808376021e-07 wk1=-1.045910090e-06 pk1=2.306440931e-13
+  k2=2.788564512e+00 lk2=-6.637268202e-07 wk2=-2.471885868e-06 pk2=5.451002717e-13
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=5.899118457e-01 ldsub=-6.178084732e-08 wdsub=-2.300892115e-07 pdsub=5.073927293e-14
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-1.668632019e+01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=3.609343152e-06 wvoff=1.344210252e-05 pvoff=-2.964252447e-12
+  nfactor={-3.614141450e+02+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=8.023751189e-05 wnfactor=2.988246952e-04 pnfactor=-6.589682180e-11
+  eta0=9.045906615e-01 leta0=-1.510803522e-07 weta0=-5.626610206e-07 peta0=1.240780083e-13
+  etab=-6.426754980e-01 letab=1.356875018e-07 wetab=5.053341779e-07 petab=-1.114362929e-13
+  u0=3.546844387e-02 lu0=-7.200181630e-09 wu0=-2.681528674e-08 pu0=5.913307032e-15
+  ua=-1.467343553e-08 lua=2.720125131e-15 wua=1.013043104e-14 pua=-2.233962654e-21
+  ub=1.405826812e-17 lub=-2.649639621e-24 wub=-9.867925890e-24 pub=2.176075017e-30
+  uc=2.793693865e-12 luc=-5.971367126e-19 wuc=-2.223881254e-18 puc=4.904102942e-25
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=-1.402307357e+07 lvsat=3.110289759e+00 wvsat=1.158350273e+01 pvsat=-2.554394021e-6
+  a0=9.565222028e+00 la0=-1.859407450e-06 wa0=-6.924901578e-06 pa0=1.527079296e-12
+  ags=1.249999977e+00 lags=6.870465086e-15 wags=7.028091886e-14 pags=-1.549834394e-20
+  a1=0.0
+  a2=-5.637236484e+00 la2=1.385404338e-06 wa2=5.159594558e-06 pa2=-1.137793792e-12
+  b0=0.0
+  b1=0.0
+  keta=5.127595502e-02 lketa=-1.113666167e-08 wketa=-4.147560895e-08 pketa=9.146201285e-15
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=6.162250608e-01 lpclm=1.290442483e-09 wpclm=4.805864056e-09 ppclm=-1.059789142e-15
+  pdiblc1=7.369041684e-01 lpdiblc1=-1.255142029e-07 wpdiblc1=-4.674465757e-07 ppdiblc1=1.030813189e-13
+  pdiblc2=4.376683139e-02 lpdiblc2=-8.800462992e-09 wpdiblc2=-3.277515210e-08 ppdiblc2=7.227576541e-15
+  pdiblcb=-2.022819590e+00 lpdiblcb=3.623434635e-07 wpdiblcb=1.349457693e-06 ppdiblcb=-2.975824105e-13
+  drout=1.000002593e+00 ldrout=-5.373826184e-13 wdrout=-1.188062981e-12 pdrout=2.619916444e-19
+  pscbe1=8.000000136e+08 lpscbe1=-2.994468689e-06 wpscbe1=-1.085488892e-05 ppscbe1=2.393722534e-12
+  pscbe2=-2.999218905e-08 lpscbe2=8.240920118e-15 wpscbe2=3.069125940e-14 ppscbe2=-6.768036523e-21
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=1.310307595e+01 lbeta0=-1.047827009e-06 wbeta0=-3.902373647e-06 pbeta0=8.605514367e-13
* Gidl Induced Drain Leakage Model Parameters
+  agidl=6.148185157e-08 lagidl=-1.350741332e-14 wagidl=-5.030500795e-14 pagidl=1.109326035e-20
+  bgidl=1.000000330e+09 lbgidl=-6.318053436e-05 wbgidl=-7.731658936e-06 pbgidl=1.704986572e-12
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-1.106e-8
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-8.015864343e+01 lkt1=1.749188092e-05 wkt1=6.514416875e-05 pkt1=-1.436559209e-11
+  kt2=-9.625899341e-02 lkt2=-2.053970327e-15 wkt2=-2.186541082e-14 pkt2=4.821759880e-21
+  at=7.812770834e+05 lat=-1.631887875e-01 wat=-6.077561245e-01 pat=1.340223806e-7
+  ute=-1.802674948e+00 lute=3.864998705e-07 wute=1.439422612e-06 pute=-3.174214743e-13
+  ua1=7.435796112e-10 lua1=5.781011115e-23 wua1=-4.454044932e-22 pua1=9.822059722e-29
+  ub1=-4.726031082e-19 lub1=6.614588398e-31 wub1=1.896854528e-30 pub1=-4.182943640e-37
+  uc1=-2.193904273e-11 luc1=9.015758513e-24 wuc1=2.397447348e-23 puc1=-5.286851059e-30
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.04e-6
+  sbref=1.04e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.108 pmos
* Model Flag Parameters
+  lmin=2.0e-05 lmax=0.0001 wmin=8.2e-07 wmax=8.4e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.126311+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+  k1=0.43165561
+  k2=0.026980026
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=3.2465718e-7
+  voff={-0.23051772+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.8768912+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+  eta0=0.08
+  etab=-0.07
+  u0=0.0095864
+  ua=-7.4757916e-10
+  ub=9.5046395e-19
+  uc=-1.0566299e-10
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=80156.0
+  a0=1.464
+  ags=0.11329
+  a1=0.0
+  a2=0.97
+  b0=-8.9873e-8
+  b1=3.3859e-9
+  keta=0.023361259
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=0.015
+  pdiblc1=0.39
+  pdiblc2=0.0012771588
+  pdiblcb=-0.225
+  drout=0.56
+  pscbe1=800000000.0
+  pscbe2=1.0060625e-8
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=0.0
+  alpha1=0.0
+  beta0=30.0
* Gidl Induced Drain Leakage Model Parameters
+  agidl=9.43573999999999e-11
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-0.43825
+  kt2=-0.058546
+  at=70990.0
+  ute=-0.08298
+  ua1=2.0902e-9
+  ub1=-1.2289e-18
+  uc1=-2.9789e-11
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.109 pmos
* Model Flag Parameters
+  lmin=8.0e-06 lmax=2.0e-05 wmin=8.2e-07 wmax=8.4e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.151793231e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=5.102439717e-07 wvth0=-7.105427358e-21
+  k1=4.210498003e-01 lk1=2.123656422e-7
+  k2=3.098838670e-02 lk2=-8.026149068e-8
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=-6.144535039e-06 lcit=1.295359998e-10 wcit=-6.776263578e-27 pcit=2.981555974e-31
+  voff={-2.428791561e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=2.475194627e-7
+  nfactor={1.918471956e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-8.325930941e-7
+  eta0=0.08
+  etab=-0.07
+  u0=9.965711908e-03 lu0=-7.595159576e-9
+  ua=-7.615294670e-10 lua=2.793342514e-16
+  ub=9.271909546e-19 lub=4.660072882e-25
+  uc=-1.283201274e-10 luc=4.536756436e-16
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=2.656289816e+04 lvsat=1.073122547e+0
+  a0=1.605375760e+00 la0=-2.830840351e-6
+  ags=2.825339191e-02 lags=1.702732223e-6
+  a1=0.0
+  a2=1.083666533e+00 la2=-2.276004104e-6
+  b0=-1.499644844e-07 lb0=1.203243040e-12
+  b1=5.649803031e-09 lb1=-4.533130761e-14
+  keta=4.023168533e-02 lketa=-3.378053190e-7
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-6.921953293e-02 lpclm=1.686371502e-06 ppclm=2.664535259e-27
+  pdiblc1=0.39
+  pdiblc2=1.917610060e-03 lpdiblc2=-1.282408862e-8
+  pdiblcb=-2.717239457e-01 lpdiblcb=9.355778616e-07 wpdiblcb=-1.776356839e-21
+  drout=0.56
+  pscbe1=8.000325956e+08 lpscbe1=-6.526776473e-1
+  pscbe2=1.315981805e-08 lpscbe2=-6.205675405e-14
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=-6.686266667e-11 lalpha0=1.338825943e-15
+  alpha1=-6.686266667e-11 lalpha1=1.338825943e-15
+  beta0=4.586076776e+01 lbeta0=-3.175884006e-4
* Gidl Induced Drain Leakage Model Parameters
+  agidl=-8.562847058e-09 lagidl=1.733477066e-13 wagidl=-1.737079286e-29 pagidl=3.176373552e-34
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=-4.251725813e-01 legidl=1.051580369e-05 pegidl=-1.421085472e-26
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.365640579e-01 lkt1=-3.375849616e-8
+  kt2=-6.268314622e-02 lkt2=8.284023011e-8
+  at=1.184558071e+05 lat=-9.504325371e-1
+  ute=-5.002598587e-02 lute=-6.598553610e-7
+  ua1=2.269041386e-09 lua1=-3.581034063e-15
+  ub1=-1.571912915e-18 lub1=6.868325966e-24
+  uc1=-4.384869988e-11 luc1=2.815246818e-16 wuc1=-2.067951531e-31 puc1=-1.654361225e-36
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.110 pmos
* Model Flag Parameters
+  lmin=4.0e-06 lmax=8.0e-06 wmin=8.2e-07 wmax=8.4e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.090414346e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=1.776925644e-8
+  k1=4.556728822e-01 lk1=-6.543334786e-8
+  k2=1.885398624e-02 lk2=1.709911408e-8
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.057269452e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-5.057204472e-8
+  nfactor={2.150233085e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-2.692133146e-06 wnfactor=-1.421085472e-20
+  eta0=0.08
+  etab=-0.07
+  u0=8.535573484e-03 lu0=3.879584672e-9
+  ua=-8.237874492e-10 lua=7.788624164e-16
+  ub=1.048518672e-18 lub=-5.074680762e-25
+  uc=-7.083802061e-11 luc=-7.533189791e-18
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=2.678104074e+05 lvsat=-8.625316685e-1
+  a0=1.347035279e+00 la0=-7.580403376e-7
+  ags=2.084960866e-01 lags=2.565513575e-7
+  a1=0.0
+  a2=0.8
+  b0=0.0
+  b1=0.0
+  keta=-8.364571240e-04 lketa=-8.294256640e-9
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=2.407132755e-01 lpclm=-8.003805848e-7
+  pdiblc1=0.39
+  pdiblc2=-1.397670217e-03 lpdiblc2=1.377612899e-08 ppdiblc2=1.387778781e-29
+  pdiblcb=-2.494013897e-01 lpdiblcb=7.564723865e-7
+  drout=0.56
+  pscbe1=1.227212561e+09 lpscbe1=-3.428139670e+3
+  pscbe2=-1.711599940e-08 lpscbe2=1.808618728e-13 wpscbe2=-5.293955920e-29 ppscbe2=2.117582368e-34
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=3.429576331e+00 lbeta0=2.285911254e-5
* Gidl Induced Drain Leakage Model Parameters
+  agidl=2.613220901e-08 lagidl=-1.050287696e-13
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=1.675517744e+00 legidl=-6.339127153e-6
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.061103840e-01 lkt1=-2.781041573e-7
+  kt2=-4.839276194e-02 lkt2=-3.181895402e-8
+  at=-9.120917488e+04 lat=7.318186388e-1
+  ute=-1.647219648e-01 lute=2.604101198e-7
+  ua1=5.703275549e-10 lua1=1.004863033e-14
+  ub1=8.239234094e-19 lub1=-1.235471470e-23 pub1=2.465190329e-44
+  uc1=-1.164852119e-11 luc1=2.316590399e-17
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.111 pmos
* Model Flag Parameters
+  lmin=2.0e-06 lmax=4.0e-06 wmin=8.2e-07 wmax=8.4e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.085843201e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-6.228379991e-10
+  k1=4.428072554e-01 lk1=-1.366824095e-8
+  k2=2.193345702e-02 lk2=4.708801823e-9
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=8.622137339e-01 ldsub=-1.215963003e-6
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.337857314e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=6.232304277e-8
+  nfactor={7.881674337e-01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=2.788165241e-6
+  eta0=1.604349200e-01 leta0=-3.236315093e-7
+  etab=-1.403185835e-01 letab=2.829282271e-7
+  u0=8.638994592e-03 lu0=3.463467775e-9
+  ua=-8.215637429e-10 lua=7.699152898e-16
+  ub=1.011504174e-18 lub=-3.585395030e-25
+  uc=-7.560382119e-11 luc=1.164210416e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=53438.0
+  a0=1.154071298e+00 la0=1.835409954e-8
+  ags=1.482758150e-01 lags=4.988488244e-7
+  a1=0.0
+  a2=0.8
+  b0=0.0
+  b1=0.0
+  keta=6.578345336e-03 lketa=-3.812786263e-08 pketa=-1.110223025e-28
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-5.559724103e-01 lpclm=2.405100206e-06 ppclm=-5.329070518e-27
+  pdiblc1=0.39
+  pdiblc2=3.641230659e-03 lpdiblc2=-6.497989463e-9
+  pdiblcb=-9.820554637e-02 lpdiblcb=1.481328872e-7
+  drout=0.56
+  pscbe1=-4.676991234e+07 lpscbe1=1.697754289e+3
+  pscbe2=4.653609693e-08 lpscbe2=-7.524360986e-14 ppscbe2=-4.235164736e-34
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=1.147359093e+01 lbeta0=-9.506141085e-6
* Gidl Induced Drain Leakage Model Parameters
+  agidl=3.821637237e-11 lagidl=-3.906838872e-17
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.816142056e-01 lkt1=2.568697892e-8
+  kt2=-6.028632264e-02 lkt2=1.603502535e-8
+  at=1.022950518e+05 lat=-4.674948746e-2
+  ute=-1.327375183e-01 lute=1.317200597e-7
+  ua1=3.323674104e-09 lua1=-1.029514575e-15
+  ub1=-2.842323112e-18 lub1=2.396501504e-24
+  uc1=1.818504214e-11 luc1=-9.687003470e-17 wuc1=-5.169878828e-32 puc1=-1.033975766e-37
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.112 pmos
* Model Flag Parameters
+  lmin=1.0e-06 lmax=2.0e-06 wmin=8.2e-07 wmax=8.4e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.101264296e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=3.058205737e-8
+  k1=3.540326720e-01 lk1=1.659689040e-7
+  k2=5.577749960e-02 lk2=-6.377529522e-8
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=-2.663045674e-01 ldsub=1.067616350e-06 pdsub=3.552713679e-27
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.021762939e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-1.639286090e-9
+  nfactor={2.430472285e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-5.350714714e-7
+  eta0=-2.241626400e-01 leta0=4.546093453e-07 weta0=2.636779683e-22 peta0=-6.383782392e-28
+  etab=8.442995791e-01 letab=-1.709466317e-06 wetab=1.228184221e-21 petab=1.214306433e-27
+  u0=1.250070846e-02 lu0=-4.350787479e-9
+  ua=2.633023699e-11 lua=-9.458151364e-16
+  ub=5.976931819e-19 lub=4.788153150e-25
+  uc=-7.509174596e-11 luc=1.060590969e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=5.963848416e+04 lvsat=-1.254680371e-2
+  a0=1.369865781e+00 la0=-4.183103528e-7
+  ags=1.727992847e-01 lags=4.492250930e-7
+  a1=0.0
+  a2=5.953062352e-01 la2=4.142019269e-7
+  b0=0.0
+  b1=0.0
+  keta=-1.079934288e-02 lketa=-2.963762975e-9
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=4.550220723e-01 lpclm=3.593326501e-7
+  pdiblc1=7.492555200e-01 lpdiblc1=-7.269607298e-7
+  pdiblc2=0.00043
+  pdiblcb=-0.025
+  drout=1.096512000e-01 ldrout=9.112898038e-7
+  pscbe1=7.983183467e+08 lpscbe1=-1.229870506e+1
+  pscbe2=9.530520115e-09 lpscbe2=-3.620850560e-16
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=5.862313582e+00 lbeta0=1.848390856e-6
* Gidl Induced Drain Leakage Model Parameters
+  agidl=2.315918186e-11 lagidl=-8.599862589e-18
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.585366557e-01 lkt1=-2.101090483e-8
+  kt2=-5.625426130e-02 lkt2=7.876068592e-9
+  at=9.703221664e+04 lat=-3.610003518e-2
+  ute=9.359355551e-01 lute=-2.030761278e-06 wute=8.881784197e-22 pute=6.217248938e-27
+  ua1=6.136533540e-09 lua1=-6.721391901e-15
+  ub1=-4.270929418e-18 lub1=5.287314936e-24 pub1=-2.465190329e-44
+  uc1=-1.285649500e-10 luc1=2.000815094e-16 wuc1=4.135903063e-31 puc1=4.135903063e-37
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=2.75e-6
+  sbref=2.74e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.113 pmos
* Model Flag Parameters
+  lmin=5.0e-07 lmax=1.0e-06 wmin=8.2e-07 wmax=8.4e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.092582479e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=2.169604366e-8
+  k1=5.229315034e-01 lk1=-6.902427879e-9
+  k2=-6.829846957e-03 lk2=3.045761312e-10
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=1.255329254e+00 ldsub=-4.898062988e-7
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={2.670066454e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-4.818574081e-07 pvoff=8.881784197e-28
+  nfactor={1.728101006e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.838195797e-7
+  eta0=-2.358444013e-02 leta0=2.493135462e-07 peta0=8.881784197e-28
+  etab=-1.689932780e+00 letab=8.843711865e-7
+  u0=1.006938082e-02 lu0=-1.862275006e-9
+  ua=-5.806459616e-10 lua=-3.245628577e-16
+  ub=8.868137281e-19 lub=1.828946535e-25
+  uc=-9.986617302e-11 luc=3.596303128e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=-5.927833243e+04 lvsat=1.091669364e-01 pvsat=-2.328306437e-22
+  a0=1.185060244e+00 la0=-2.291581900e-7
+  ags=-5.662276608e-02 lags=6.840431505e-7
+  a1=0.0
+  a2=1.050779681e+00 la2=-5.198425436e-8
+  b0=-9.183315919e-17 lb0=9.399307509e-23
+  b1=-3.817924830e-20 lb1=3.907722422e-26
+  keta=1.192995869e-02 lketa=-2.622765772e-08 pketa=-5.551115123e-29
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=1.588106337e+00 lpclm=-8.004017569e-7
+  pdiblc1=6.353741327e-02 lpdiblc1=-2.511453323e-8
+  pdiblc2=7.762209763e-04 lpdiblc2=-3.543640937e-10
+  pdiblcb=-1.404746093e-02 lpdiblcb=-1.121014279e-8
+  drout=1.039619329e+00 ldrout=-4.055117553e-8
+  pscbe1=8.256802058e+08 lpscbe1=-4.030411509e+1
+  pscbe2=3.429057487e-09 lpscbe2=5.882883972e-15
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=6.559046608e+00 lbeta0=1.135270669e-6
* Gidl Induced Drain Leakage Model Parameters
+  agidl=3.020804646e-11 lagidl=-1.581451648e-17
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.216831793e-01 lkt1=-5.873117501e-8
+  kt2=-6.301890653e-02 lkt2=1.479981827e-8
+  at=8.604123040e+04 lat=-2.485054094e-2
+  ute=-1.934483867e+00 lute=9.071704088e-7
+  ua1=-3.495144579e-09 lua1=3.136823287e-15 wua1=3.308722450e-30 pua1=-3.308722450e-36
+  ub1=4.257545597e-18 lub1=-3.441749811e-24 pub1=6.162975822e-45
+  uc1=3.311138654e-10 luc1=-2.704089518e-16 puc1=8.271806126e-37
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.75e-6
+  sbref=1.74e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.114 pmos
* Model Flag Parameters
+  lmin=2.5e-07 lmax=5.0e-07 wmin=8.2e-07 wmax=8.4e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.045892418e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-2.747137143e-9
+  k1=4.352213524e-01 lk1=3.901559036e-8
+  k2=1.408936088e-02 lk2=-1.064704755e-8
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=-1.888704683e-01 ldsub=2.662611400e-07 pdsub=8.881784197e-28
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-8.564575735e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=1.062985797e-7
+  nfactor={1.710086311e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.932506331e-7
+  eta0=4.117672797e-01 leta0=2.139821381e-8
+  etab=-1.291129272e-03 letab=3.335097045e-10
+  u0=7.485205816e-03 lu0=-5.094077095e-10
+  ua=-1.063421140e-09 lua=-7.182039643e-17
+  ub=1.148080500e-18 lub=4.611627323e-26
+  uc=-6.419271038e-11 luc=1.728726011e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=1.425608788e+05 lvsat=3.500072552e-3
+  a0=8.919849864e-01 la0=-7.572743094e-8
+  ags=9.698322768e-01 lags=1.466734064e-7
+  a1=0.0
+  a2=1.121568012e+00 la2=-8.904336116e-8
+  b0=1.836663184e-16 lb0=-5.023641140e-23
+  b1=7.635849659e-20 lb1=-2.088557599e-26
+  keta=-4.524308758e-02 lketa=3.703575468e-9
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-5.731343976e-01 lpclm=3.310509927e-07 wpclm=-8.881784197e-22 ppclm=6.661338148e-28
+  pdiblc1=-4.101030779e-01 lpdiblc1=2.228457367e-07 wpdiblc1=6.661338148e-22 ppdiblc1=-1.110223025e-28
+  pdiblc2=-9.175377595e-03 lpdiblc2=4.855496791e-09 wpdiblc2=-1.561251128e-23 ppdiblc2=-5.854691731e-30
+  pdiblcb=2.408596814e-01 lpdiblcb=-1.446591300e-07 wpdiblcb=4.440892099e-22 ppdiblcb=-3.330669074e-28
+  drout=1.436421824e+00 ldrout=-2.482852179e-7
+  pscbe1=6.925891618e+08 lpscbe1=2.937170827e+1
+  pscbe2=2.103542680e-08 lpscbe2=-3.334402489e-15
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=8.528056950e+00 lbeta0=1.044543745e-7
* Gidl Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=7.372237654e+08 lbgidl=1.375686143e+2
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.00074326333
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.5407449e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-5.460023937e-01 lkt1=6.352420121e-9
+  kt2=-1.498550792e-02 lkt2=-1.034662657e-8
+  at=6.500485322e+03 lat=1.679062992e-2
+  ute=4.908242408e-01 lute=-3.625268917e-07 wute=-1.776356839e-21 pute=4.440892099e-28
+  ua1=4.905387581e-09 lua1=-1.261023309e-15
+  ub1=-4.666106948e-18 lub1=1.229960769e-24
+  uc1=-2.811617509e-10 luc1=5.012957887e-17
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.1e-6
+  sbref=1.1e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.115 pmos
* Model Flag Parameters
+  lmin=1.8e-07 lmax=2.5e-07 wmin=8.2e-07 wmax=8.4e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-6.136775425e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-1.209665498e-07 wvth0=-3.330019835e-07 pvth0=9.108270251e-14
+  k1=-1.323742875e+00 lk1=5.201274859e-07 wk1=2.893998836e-07 pk1=-7.915665615e-14
+  k2=-5.144293646e-01 lk2=1.339133943e-07 wk2=8.711098293e-07 pk2=-2.382659605e-13
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=3.287138683e+00 ldsub=-6.844968832e-07 wdsub=-9.214571771e-07 pdsub=2.520369671e-13
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={6.645511476e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-1.945639995e-06 wvoff=-6.197584248e-06 pvoff=1.695163244e-12
+  nfactor={2.132878379e+02+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-5.767749598e-05 wnfactor=-1.732427450e-04 pnfactor=4.738535561e-11
+  eta0=3.719710767e+00 leta0=-8.833904888e-07 weta0=-2.006528872e-06 peta0=5.488257770e-13
+  etab=3.187780279e-01 letab=-8.721180617e-08 wetab=-1.966837002e-07 petab=5.379692568e-14
+  u0=-5.411772392e-03 lu0=3.018173770e-09 wu0=1.576077387e-08 pu0=-4.310886868e-15
+  ua=1.295367533e-09 lua=-7.169962742e-16 wua=2.645110211e-16 pua=-7.234905449e-23
+  ub=-7.292222104e-19 lub=5.595961105e-25 wub=-5.369217482e-26 pub=1.468588366e-32
+  uc=-1.253042192e-10 luc=3.400248001e-17 wuc=9.952755882e-17 puc=-2.722277789e-23
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=3.668737326e+06 lvsat=-9.609797092e-01 wvsat=-2.708534880e+00 pvsat=7.408384605e-7
+  a0=-3.205044165e+00 la0=1.044891983e-06 wa0=1.900097032e-06 pa0=-5.197145403e-13
+  ags=2.250599016e+00 lags=-2.036419122e-07 wags=-2.503131213e-14 pags=6.846562428e-21
+  a1=0.0
+  a2=2.169154490e+00 la2=-3.755792148e-07 wa2=-7.675998812e-07 pa2=2.099539195e-13
+  b0=0.0
+  b1=0.0
+  keta=-2.465179654e-01 lketa=5.875628005e-08 wketa=9.887401625e-08 pketa=-2.704402092e-14
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=6.693889164e-01 lpclm=-8.803984157e-09 wpclm=9.678832864e-09 ppclm=-2.647354365e-15
+  pdiblc1=2.785383071e+00 lpdiblc1=-6.511836349e-07 wpdiblc1=-1.389580021e-06 ppdiblc1=3.800779274e-13
+  pdiblc2=-1.387835366e-03 lpdiblc2=2.725448240e-09 wpdiblc2=1.944773556e-08 ppdiblc2=-5.319344629e-15
+  pdiblcb=-6.879811727e+00 lpdiblcb=1.802986914e-06 wpdiblcb=5.632537432e-06 ppdiblcb=-1.540611638e-12
+  drout=-8.416464080e-01 ldrout=3.748120050e-07 wdrout=1.129703094e-12 pdrout=-3.089963911e-19
+  pscbe1=7.998956583e+08 lpscbe1=2.123534760e-02 wpscbe1=-3.383621216e-06 ppscbe1=9.254913330e-13
+  pscbe2=-6.974408175e-09 lpscbe2=4.326847573e-15 wpscbe2=1.649352321e-14 ppscbe2=-4.511308469e-21
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=1.055619196e+01 lbeta0=-4.502811130e-07 wbeta0=-1.846049774e-08 pbeta0=5.049315343e-15
* Gidl Induced Drain Leakage Model Parameters
+  agidl=-2.737565562e-08 lagidl=7.487789324e-15 wagidl=2.193534633e-14 pagidl=-5.999755928e-21
+  bgidl=1.938486441e+09 lbgidl=-1.910007526e+02 wbgidl=-1.255871582e-05 pbgidl=3.435058594e-12
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.00074326333
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.5407449e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=3.503431887e+01 lkt1=-9.725577051e-06 wkt1=-2.845036624e-05 pkt1=7.781744175e-12
+  kt2=4.841924118e-01 lkt2=-1.468817712e-07 wkt2=-3.372881892e-07 pkt2=9.225506552e-14
+  at=-6.222650337e+04 lat=3.558883587e-02 wat=1.704428721e-01 pat=-4.661953438e-8
+  ute=-7.028629373e+00 lute=1.694194061e-06 wute=3.213560127e-06 pute=-8.789729658e-13
+  ua1=-4.563875964e-09 lua1=1.329009656e-15 wua1=2.919460567e-15 pua1=-7.985308542e-22
+  ub1=3.952316636e-18 lub1=-1.127350450e-24 wub1=-2.660820307e-24 pub1=7.277875704e-31
+  uc1=-3.851865440e-10 luc1=7.858244028e-17 wuc1=5.460638120e-17 puc1=-1.493593739e-23
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.1e-6
+  sbref=1.1e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.116 pmos
* Model Flag Parameters
+  lmin=1.5e-07 lmax=1.8e-07 wmin=8.2e-07 wmax=8.4e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-2.026e-8
+  vth0={-1.795143098e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=1.294659139e-07 wvth0=5.966985481e-07 pvth0=-1.063267320e-13
+  k1=1.231916698e+00 lk1=-3.797529189e-13 wk1=-9.953965721e-08 pk1=3.458469280e-19
+  k2=-3.799091694e-01 lk2=1.154347698e-07 wk2=1.302928486e-07 pk2=-9.480332564e-14
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=-7.615957108e-02 ldsub=1.709356880e-12 wdsub=3.169365931e-07 pdsub=-1.010960535e-18
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.914438770e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=1.169476025e-12 wvoff=2.131641919e-06 pvoff=-9.383077995e-19
+  nfactor={-1.726040546e+02+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=2.260159018e-05 wnfactor=1.437602548e-04 pnfactor=-1.856205310e-11
+  eta0=-6.208466612e-01 leta0=-2.611834482e-13 weta0=6.901379403e-07 peta0=1.597411927e-19
+  etab=-1.097401186e-01 letab=2.242988286e-13 wetab=6.764927297e-08 petab=-1.311298694e-19
+  u0=-7.226761977e-03 lu0=3.670522949e-09 wu0=8.249090357e-09 pu0=-3.014498258e-15
+  ua=-2.227607364e-09 lua=-4.584191544e-22 wua=-9.097914396e-17 pua=3.292879493e-28
+  ub=2.020361843e-18 lub=8.278891576e-31 wub=1.846947385e-26 pub=-4.930923246e-37
+  uc=4.176772084e-11 luc=-1.332166199e-24 wuc=-3.423215834e-17 puc=-2.739104635e-31
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=1.567620174e+06 lvsat=-5.779118691e-01 wvsat=-1.220697507e+00 pvsat=4.746227064e-7
+  a0=1.929051414e+00 la0=9.213504484e-13 wa0=-6.535284660e-07 pa0=-7.355759166e-19
+  ags=1.249999989e+00 lags=2.073733185e-15 wags=6.102618499e-14 pags=-1.155895291e-20
+  a1=0.0
+  a2=3.237378198e-01 la2=-1.520076864e-14 wa2=2.640132694e-07 pa2=1.201360789e-20
+  b0=0.0
+  b1=0.0
+  keta=4.218281402e-02 lketa=-1.111449523e-13 wketa=-3.400766685e-08 pketa=6.416587225e-20
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=6.261299533e-01 lpclm=8.669641005e-14 wpclm=-3.328746847e-09 ppclm=-5.606420572e-20
+  pdiblc1=-4.142237009e-01 lpdiblc1=3.634762766e-13 wpdiblc1=4.779425119e-07 ppdiblc1=-2.801234755e-19
+  pdiblc2=1.200367986e-02 lpdiblc2=7.651560968e-15 wpdiblc2=-6.688965112e-09 ppdiblc2=-3.585787722e-21
+  pdiblcb=1.979201262e+00 lpdiblcb=6.395183334e-13 wpdiblcb=-1.937289976e-06 ppdiblcb=-3.946861966e-19
+  drout=1.000004514e+00 ldrout=-8.567691552e-13 wdrout=-2.766096316e-12 pdrout=5.242948689e-19
+  pscbe1=7.999999852e+08 lpscbe1=2.968872070e-06 wpscbe1=1.251791382e-05 ppscbe1=-2.503814697e-12
+  pscbe2=1.428565304e-08 lpscbe2=-9.259324781e-23 wpscbe2=-5.672892524e-15 ppscbe2=5.001148277e-28
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=8.343718675e+00 lbeta0=1.570862707e-12 wbeta0=6.353218810e-09 pbeta0=-8.367560440e-19
* Gidl Induced Drain Leakage Model Parameters
+  agidl=9.415762829e-09 lagidl=-1.709634062e-22 wagidl=-7.544587114e-15 pagidl=1.369881918e-28
+  bgidl=1.000000352e+09 lbgidl=-6.917549896e-05 wbgidl=-2.573889160e-05 pbgidl=6.628479004e-12
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-1.106e-8
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-1.275250163e+01 lkt1=-3.622959802e-12 wkt1=9.785391861e-06 pkt1=2.909716002e-18
+  kt2=-2.375137447e-01 lkt2=-1.454123630e-13 wkt2=1.160085502e-07 pkt2=1.225579940e-19
+  at=1.126398909e+05 lat=2.957911044e-08 wat=-5.862312017e-02 pat=-2.560526552e-14
+  ute=1.295830162e+00 lute=6.090733606e-14 wute=-1.105292877e-06 pute=-2.684970912e-21
+  ua1=1.966235506e-09 lua1=1.483836552e-21 wua1=-1.004133498e-15 pua1=-1.072934993e-27
+  ub1=-1.586945149e-18 lub1=1.181096969e-31 wub1=9.151798138e-25 pub1=2.794307721e-38
+  uc1=9.299026423e-13 luc1=2.282398126e-23 wuc1=-1.878160053e-17 puc1=-1.662715749e-29
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.04e-6
+  sbref=1.04e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.117 pmos
* Model Flag Parameters
+  lmin=2.0e-05 lmax=0.0001 wmin=7.9e-07 wmax=8.2e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.126311+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+  k1=0.43165561
+  k2=0.026980026
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=3.2465718e-7
+  voff={-0.23051772+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.8768912+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+  eta0=0.08
+  etab=-0.07
+  u0=0.0095864
+  ua=-7.4757916e-10
+  ub=9.5046395e-19
+  uc=-1.0566299e-10
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=80156.0
+  a0=1.464
+  ags=0.11329
+  a1=0.0
+  a2=0.97
+  b0=-8.9873e-8
+  b1=3.3859e-9
+  keta=0.023361259
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=0.015
+  pdiblc1=0.39
+  pdiblc2=0.0012771588
+  pdiblcb=-0.225
+  drout=0.56
+  pscbe1=800000000.0
+  pscbe2=1.0060625e-8
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=0.0
+  alpha1=0.0
+  beta0=30.0
* Gidl Induced Drain Leakage Model Parameters
+  agidl=9.43573999999999e-11
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-0.43825
+  kt2=-0.058546
+  at=70990.0
+  ute=-0.08298
+  ua1=2.0902e-9
+  ub1=-1.2289e-18
+  uc1=-2.9789e-11
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.118 pmos
* Model Flag Parameters
+  lmin=8.0e-06 lmax=2.0e-05 wmin=7.9e-07 wmax=8.2e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.151793231e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=5.102439717e-7
+  k1=4.210498003e-01 lk1=2.123656422e-7
+  k2=3.098838670e-02 lk2=-8.026149068e-8
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=-6.144535039e-06 lcit=1.295359998e-10 wcit=-3.388131789e-27 pcit=-1.355252716e-32
+  voff={-2.428791561e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=2.475194627e-07 wvoff=8.881784197e-22
+  nfactor={1.918471956e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-8.325930941e-7
+  eta0=0.08
+  etab=-0.07
+  u0=9.965711908e-03 lu0=-7.595159576e-9
+  ua=-7.615294670e-10 lua=2.793342514e-16
+  ub=9.271909546e-19 lub=4.660072882e-25
+  uc=-1.283201274e-10 luc=4.536756436e-16 wuc=4.135903063e-31
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=2.656289816e+04 lvsat=1.073122547e+0
+  a0=1.605375760e+00 la0=-2.830840351e-06 wa0=7.105427358e-21
+  ags=2.825339191e-02 lags=1.702732223e-06 pags=3.552713679e-27
+  a1=0.0
+  a2=1.083666533e+00 la2=-2.276004104e-6
+  b0=-1.499644844e-07 lb0=1.203243040e-12
+  b1=5.649803031e-09 lb1=-4.533130761e-14
+  keta=4.023168533e-02 lketa=-3.378053190e-7
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-6.921953293e-02 lpclm=1.686371502e-06 wpclm=1.110223025e-22 ppclm=1.776356839e-27
+  pdiblc1=0.39
+  pdiblc2=1.917610060e-03 lpdiblc2=-1.282408862e-8
+  pdiblcb=-2.717239457e-01 lpdiblcb=9.355778616e-7
+  drout=0.56
+  pscbe1=8.000325956e+08 lpscbe1=-6.526776473e-1
+  pscbe2=1.315981805e-08 lpscbe2=-6.205675405e-14
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=-6.686266667e-11 lalpha0=1.338825943e-15
+  alpha1=-6.686266667e-11 lalpha1=1.338825943e-15
+  beta0=4.586076776e+01 lbeta0=-3.175884006e-4
* Gidl Induced Drain Leakage Model Parameters
+  agidl=-8.562847058e-09 lagidl=1.733477066e-13 wagidl=-1.033975766e-29 pagidl=1.985233470e-35
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=-4.251725813e-01 legidl=1.051580369e-05 pegidl=-3.552713679e-27
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.365640579e-01 lkt1=-3.375849616e-08 wkt1=-1.776356839e-21
+  kt2=-6.268314622e-02 lkt2=8.284023011e-8
+  at=1.184558071e+05 lat=-9.504325371e-1
+  ute=-5.002598587e-02 lute=-6.598553610e-7
+  ua1=2.269041386e-09 lua1=-3.581034063e-15
+  ub1=-1.571912915e-18 lub1=6.868325966e-24 wub1=6.162975822e-39
+  uc1=-4.384869988e-11 luc1=2.815246818e-16
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.119 pmos
* Model Flag Parameters
+  lmin=4.0e-06 lmax=8.0e-06 wmin=7.9e-07 wmax=8.2e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.090414346e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=1.776925644e-8
+  k1=4.556728822e-01 lk1=-6.543334786e-8
+  k2=1.885398624e-02 lk2=1.709911408e-8
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.057269452e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-5.057204472e-8
+  nfactor={2.150233085e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-2.692133146e-6
+  eta0=0.08
+  etab=-0.07
+  u0=8.535573484e-03 lu0=3.879584672e-9
+  ua=-8.237874492e-10 lua=7.788624164e-16
+  ub=1.048518672e-18 lub=-5.074680762e-25
+  uc=-7.083802061e-11 luc=-7.533189791e-18
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=2.678104074e+05 lvsat=-8.625316685e-1
+  a0=1.347035279e+00 la0=-7.580403376e-7
+  ags=2.084960866e-01 lags=2.565513575e-7
+  a1=0.0
+  a2=0.8
+  b0=0.0
+  b1=0.0
+  keta=-8.364571240e-04 lketa=-8.294256640e-9
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=2.407132755e-01 lpclm=-8.003805848e-7
+  pdiblc1=0.39
+  pdiblc2=-1.397670217e-03 lpdiblc2=1.377612899e-08 wpdiblc2=1.734723476e-24 ppdiblc2=6.938893904e-30
+  pdiblcb=-2.494013897e-01 lpdiblcb=7.564723865e-07 wpdiblcb=8.881784197e-22
+  drout=0.56
+  pscbe1=1.227212561e+09 lpscbe1=-3.428139670e+3
+  pscbe2=-1.711599940e-08 lpscbe2=1.808618728e-13 ppscbe2=-1.058791184e-34
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=3.429576331e+00 lbeta0=2.285911254e-5
* Gidl Induced Drain Leakage Model Parameters
+  agidl=2.613220901e-08 lagidl=-1.050287696e-13
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=1.675517744e+00 legidl=-6.339127153e-6
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.061103840e-01 lkt1=-2.781041573e-7
+  kt2=-4.839276194e-02 lkt2=-3.181895402e-8
+  at=-9.120917488e+04 lat=7.318186388e-1
+  ute=-1.647219648e-01 lute=2.604101198e-7
+  ua1=5.703275549e-10 lua1=1.004863033e-14
+  ub1=8.239234094e-19 lub1=-1.235471470e-23 pub1=-2.465190329e-44
+  uc1=-1.164852119e-11 luc1=2.316590399e-17
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.120 pmos
* Model Flag Parameters
+  lmin=2.0e-06 lmax=4.0e-06 wmin=7.9e-07 wmax=8.2e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.085843201e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-6.228379991e-10
+  k1=4.428072554e-01 lk1=-1.366824095e-8
+  k2=2.193345702e-02 lk2=4.708801823e-9
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=8.622137339e-01 ldsub=-1.215963003e-6
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.337857314e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=6.232304277e-8
+  nfactor={7.881674337e-01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=2.788165241e-6
+  eta0=1.604349200e-01 leta0=-3.236315093e-7
+  etab=-1.403185835e-01 letab=2.829282271e-7
+  u0=8.638994592e-03 lu0=3.463467775e-9
+  ua=-8.215637429e-10 lua=7.699152898e-16
+  ub=1.011504174e-18 lub=-3.585395030e-25
+  uc=-7.560382119e-11 luc=1.164210416e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=53438.0
+  a0=1.154071298e+00 la0=1.835409954e-8
+  ags=1.482758150e-01 lags=4.988488244e-7
+  a1=0.0
+  a2=0.8
+  b0=0.0
+  b1=0.0
+  keta=6.578345336e-03 lketa=-3.812786263e-08 wketa=1.387778781e-23 pketa=2.775557562e-29
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-5.559724103e-01 lpclm=2.405100206e-06 wpclm=-4.440892099e-22 ppclm=-8.881784197e-28
+  pdiblc1=0.39
+  pdiblc2=3.641230659e-03 lpdiblc2=-6.497989463e-9
+  pdiblcb=-9.820554637e-02 lpdiblcb=1.481328872e-7
+  drout=0.56
+  pscbe1=-4.676991234e+07 lpscbe1=1.697754289e+03 ppscbe1=-3.814697266e-18
+  pscbe2=4.653609693e-08 lpscbe2=-7.524360986e-14
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=1.147359093e+01 lbeta0=-9.506141085e-6
* Gidl Induced Drain Leakage Model Parameters
+  agidl=3.821637237e-11 lagidl=-3.906838872e-17
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.816142056e-01 lkt1=2.568697892e-8
+  kt2=-6.028632264e-02 lkt2=1.603502535e-8
+  at=1.022950518e+05 lat=-4.674948746e-2
+  ute=-1.327375183e-01 lute=1.317200597e-7
+  ua1=3.323674104e-09 lua1=-1.029514575e-15
+  ub1=-2.842323112e-18 lub1=2.396501504e-24
+  uc1=1.818504214e-11 luc1=-9.687003470e-17 puc1=-2.067951531e-37
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.121 pmos
* Model Flag Parameters
+  lmin=1.0e-06 lmax=2.0e-06 wmin=7.9e-07 wmax=8.2e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.101264296e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=3.058205737e-8
+  k1=3.540326720e-01 lk1=1.659689040e-7
+  k2=5.577749960e-02 lk2=-6.377529522e-8
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=-2.663045674e-01 ldsub=1.067616350e-06 pdsub=-1.776356839e-27
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.021762939e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-1.639286090e-9
+  nfactor={2.430472285e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-5.350714714e-7
+  eta0=-2.241626400e-01 leta0=4.546093453e-07 weta0=-2.775557562e-22 peta0=-2.567390744e-28
+  etab=8.442995791e-01 letab=-1.709466317e-06 wetab=-5.481726184e-22 petab=2.914335440e-28
+  u0=1.250070846e-02 lu0=-4.350787479e-9
+  ua=2.633023699e-11 lua=-9.458151364e-16
+  ub=5.976931819e-19 lub=4.788153150e-25
+  uc=-7.509174596e-11 luc=1.060590969e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=5.963848416e+04 lvsat=-1.254680371e-2
+  a0=1.369865781e+00 la0=-4.183103528e-7
+  ags=1.727992847e-01 lags=4.492250930e-7
+  a1=0.0
+  a2=5.953062352e-01 la2=4.142019269e-7
+  b0=0.0
+  b1=0.0
+  keta=-1.079934288e-02 lketa=-2.963762975e-9
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=4.550220723e-01 lpclm=3.593326501e-7
+  pdiblc1=7.492555200e-01 lpdiblc1=-7.269607298e-7
+  pdiblc2=0.00043
+  pdiblcb=-0.025
+  drout=1.096512000e-01 ldrout=9.112898038e-7
+  pscbe1=7.983183467e+08 lpscbe1=-1.229870506e+1
+  pscbe2=9.530520115e-09 lpscbe2=-3.620850560e-16
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=5.862313582e+00 lbeta0=1.848390856e-6
* Gidl Induced Drain Leakage Model Parameters
+  agidl=2.315918186e-11 lagidl=-8.599862589e-18
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.585366557e-01 lkt1=-2.101090483e-8
+  kt2=-5.625426130e-02 lkt2=7.876068592e-9
+  at=9.703221664e+04 lat=-3.610003518e-2
+  ute=9.359355551e-01 lute=-2.030761278e-06 wute=-4.440892099e-22 pute=-8.881784197e-28
+  ua1=6.136533540e-09 lua1=-6.721391901e-15
+  ub1=-4.270929418e-18 lub1=5.287314936e-24 pub1=-1.232595164e-44
+  uc1=-1.285649500e-10 luc1=2.000815094e-16 puc1=4.135903063e-37
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=2.75e-6
+  sbref=2.74e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.122 pmos
* Model Flag Parameters
+  lmin=5.0e-07 lmax=1.0e-06 wmin=7.9e-07 wmax=8.2e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.092582479e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=2.169604366e-8
+  k1=5.229315034e-01 lk1=-6.902427879e-9
+  k2=-6.829846957e-03 lk2=3.045761312e-10
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=1.255329254e+00 ldsub=-4.898062988e-7
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={2.670066454e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-4.818574081e-7
+  nfactor={1.728101006e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.838195797e-7
+  eta0=-2.358444013e-02 leta0=2.493135462e-7
+  etab=-1.689932780e+00 letab=8.843711865e-7
+  u0=1.006938082e-02 lu0=-1.862275006e-9
+  ua=-5.806459616e-10 lua=-3.245628577e-16
+  ub=8.868137281e-19 lub=1.828946535e-25
+  uc=-9.986617302e-11 luc=3.596303128e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=-5.927833243e+04 lvsat=1.091669364e-1
+  a0=1.185060244e+00 la0=-2.291581900e-7
+  ags=-5.662276608e-02 lags=6.840431505e-7
+  a1=0.0
+  a2=1.050779681e+00 la2=-5.198425436e-8
+  b0=-9.183315919e-17 lb0=9.399307509e-23
+  b1=-3.817924830e-20 lb1=3.907722422e-26
+  keta=1.192995869e-02 lketa=-2.622765772e-08 pketa=-5.551115123e-29
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=1.588106337e+00 lpclm=-8.004017569e-7
+  pdiblc1=6.353741327e-02 lpdiblc1=-2.511453323e-08 ppdiblc1=-1.110223025e-28
+  pdiblc2=7.762209763e-04 lpdiblc2=-3.543640937e-10
+  pdiblcb=-1.404746093e-02 lpdiblcb=-1.121014279e-8
+  drout=1.039619329e+00 ldrout=-4.055117553e-8
+  pscbe1=8.256802058e+08 lpscbe1=-4.030411509e+1
+  pscbe2=3.429057487e-09 lpscbe2=5.882883972e-15
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=6.559046608e+00 lbeta0=1.135270669e-6
* Gidl Induced Drain Leakage Model Parameters
+  agidl=3.020804646e-11 lagidl=-1.581451648e-17
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.216831793e-01 lkt1=-5.873117501e-8
+  kt2=-6.301890653e-02 lkt2=1.479981827e-8
+  at=8.604123040e+04 lat=-2.485054094e-2
+  ute=-1.934483867e+00 lute=9.071704088e-7
+  ua1=-3.495144579e-09 lua1=3.136823287e-15 wua1=6.617444900e-30 pua1=-4.963083675e-36
+  ub1=4.257545597e-18 lub1=-3.441749811e-24 wub1=-6.162975822e-39
+  uc1=3.311138654e-10 luc1=-2.704089518e-16 wuc1=4.135903063e-31 puc1=-4.135903063e-37
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.75e-6
+  sbref=1.74e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.123 pmos
* Model Flag Parameters
+  lmin=2.5e-07 lmax=5.0e-07 wmin=7.9e-07 wmax=8.2e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.045892418e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-2.747137143e-9
+  k1=4.352213524e-01 lk1=3.901559036e-8
+  k2=1.408936088e-02 lk2=-1.064704755e-08 pk2=1.387778781e-29
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=-1.888704683e-01 ldsub=2.662611400e-7
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-8.564575735e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=1.062985797e-07 wvoff=3.552713679e-21
+  nfactor={1.710086311e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.932506331e-7
+  eta0=4.117672797e-01 leta0=2.139821381e-8
+  etab=-1.291129272e-03 letab=3.335097045e-10
+  u0=7.485205816e-03 lu0=-5.094077095e-10
+  ua=-1.063421140e-09 lua=-7.182039643e-17
+  ub=1.148080500e-18 lub=4.611627323e-26
+  uc=-6.419271038e-11 luc=1.728726011e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=1.425608788e+05 lvsat=3.500072552e-3
+  a0=8.919849864e-01 la0=-7.572743094e-8
+  ags=9.698322768e-01 lags=1.466734064e-7
+  a1=0.0
+  a2=1.121568012e+00 la2=-8.904336116e-8
+  b0=1.836663184e-16 lb0=-5.023641140e-23
+  b1=7.635849659e-20 lb1=-2.088557599e-26
+  keta=-4.524308758e-02 lketa=3.703575468e-9
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-5.731343976e-01 lpclm=3.310509927e-07 wpclm=4.440892099e-22 ppclm=-2.220446049e-28
+  pdiblc1=-4.101030779e-01 lpdiblc1=2.228457367e-07 wpdiblc1=2.220446049e-22 ppdiblc1=-2.775557562e-28
+  pdiblc2=-9.175377595e-03 lpdiblc2=4.855496791e-09 wpdiblc2=-1.214306433e-23 ppdiblc2=1.084202172e-30
+  pdiblcb=2.408596814e-01 lpdiblcb=-1.446591300e-07 wpdiblcb=4.440892099e-22
+  drout=1.436421824e+00 ldrout=-2.482852179e-7
+  pscbe1=6.925891618e+08 lpscbe1=2.937170827e+1
+  pscbe2=2.103542680e-08 lpscbe2=-3.334402489e-15
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=8.528056950e+00 lbeta0=1.044543745e-7
* Gidl Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=7.372237654e+08 lbgidl=1.375686143e+2
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.00074326333
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.5407449e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-5.460023937e-01 lkt1=6.352420121e-9
+  kt2=-1.498550792e-02 lkt2=-1.034662657e-8
+  at=6.500485322e+03 lat=1.679062992e-2
+  ute=4.908242408e-01 lute=-3.625268917e-7
+  ua1=4.905387581e-09 lua1=-1.261023309e-15
+  ub1=-4.666106948e-18 lub1=1.229960769e-24
+  uc1=-2.811617509e-10 luc1=5.012957887e-17
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.1e-6
+  sbref=1.1e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.124 pmos
* Model Flag Parameters
+  lmin=1.8e-07 lmax=2.5e-07 wmin=7.9e-07 wmax=8.2e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.029269231e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-7.293911197e-9
+  k1=-9.625672899e-01 lk1=4.213387398e-7
+  k2=5.727293397e-01 lk2=-1.634462546e-07 wk2=-4.440892099e-22 pk2=-2.220446049e-28
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=2.137145701e+00 ldsub=-3.699508026e-7
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-1.089170690e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=1.699502713e-7
+  nfactor={-2.921819978e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.460169641e-6
+  eta0=1.215531322e+00 leta0=-1.984473271e-7
+  etab=7.331369097e-02 letab=-2.007240073e-08 wetab=1.647987302e-23 petab=-8.673617380e-30
+  u0=1.425792013e-02 lu0=-2.361880528e-9
+  ua=1.625481428e-09 lua=-8.072890268e-16
+  ub=-7.962308851e-19 lub=5.779243232e-25
+  uc=-1.092267674e-12 luc=2.802702628e-20
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=2.884433928e+05 lvsat=-3.640171267e-2
+  a0=-8.336933221e-01 la0=3.962801000e-7
+  ags=2.250598985e+00 lags=-2.036419037e-7
+  a1=0.0
+  a2=1.211177822e+00 la2=-1.135534364e-7
+  b0=0.0
+  b1=0.0
+  keta=-1.231216453e-01 lketa=2.500491856e-8
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=6.814682513e-01 lpclm=-1.210792385e-8
+  pdiblc1=1.051165451e+00 lpdiblc1=-1.768404313e-7
+  pdiblc2=2.288324307e-02 lpdiblc2=-3.913177133e-9
+  pdiblcb=1.496831658e-01 lpdiblcb=-1.197205294e-7
+  drout=-8.416449981e-01 ldrout=3.748116193e-7
+  pscbe1=7.998956541e+08 lpscbe1=2.123650263e-2
+  pscbe2=1.360976700e-08 lpscbe2=-1.303336022e-15
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=1.053315297e+01 lbeta0=-4.439794884e-7
* Gidl Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=1.938486425e+09 lbgidl=-1.910007483e+2
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.00074326333
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.5407449e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.721835984e-01 lkt1=-1.383849677e-8
+  kt2=6.325147130e-02 lkt2=-3.174600512e-8
+  at=1.504888693e+05 lat=-2.259307287e-2
+  ute=-3.018056026e+00 lute=5.972220390e-07 pute=1.776356839e-27
+  ua1=-9.203434720e-10 lua1=3.324306487e-16
+  ub1=6.315712371e-19 lub1=-2.190601681e-25
+  uc1=-3.170369254e-10 luc1=5.994215660e-17
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.1e-6
+  sbref=1.1e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.125 pmos
* Model Flag Parameters
+  lmin=1.5e-07 lmax=1.8e-07 wmin=7.9e-07 wmax=8.2e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-2.026e-8
+  vth0={-1.313143993e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=5.469689174e-08 wvth0=2.104861606e-07 pvth0=-4.641640813e-14
+  k1=3.187794420e-01 lk1=1.739705304e-07 wk1=6.321316583e-07 pk1=-1.393976733e-13
+  k2=-2.343119070e-01 lk2=8.698360709e-10 wk2=1.362983893e-08 pk2=-3.005652080e-15
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=2.831294506e+00 ldsub=-5.539264412e-07 wdsub=-2.012724951e-06 pdsub=4.438461061e-13
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-1.146439752e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=1.967751696e-07 wvoff=7.149938099e-07 pvoff=-1.576704350e-13
+  nfactor={-2.266678388e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=5.936296868e-06 wnfactor=2.361971794e-05 pnfactor=-5.208620201e-12
+  eta0=5.710310891e+00 leta0=-1.206212398e-06 weta0=-4.382841334e-06 peta0=9.665041709e-13
+  etab=5.108517495e-01 letab=-1.182349385e-07 wetab=-4.296136144e-07 petab=9.473839425e-14
+  u0=-6.166418921e-05 lu0=5.985866220e-10 wu0=2.507898122e-09 pu0=-5.530416939e-16
+  ua=-3.062213224e-09 lua=1.590086471e-16 wua=5.777671626e-16 pua=-1.274092147e-22
+  ub=2.189775517e-18 lub=-3.227586245e-26 wub=-1.172769596e-25 pub=2.586191513e-32
+  uc=-2.722694536e-10 luc=5.983036117e-17 wuc=2.173970365e-16 puc=-4.794039450e-23
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=-2.153950831e+05 lvsat=7.166411754e-02 wvsat=2.079826933e-01 pvsat=-4.586434353e-8
+  a0=-4.066283983e+00 la0=1.142232220e-06 wa0=4.150365918e-06 pa0=-9.152386923e-13
+  ags=1.250000065e+00 lags=-1.235200386e-14
+  a1=0.0
+  a2=2.745729274e+00 la2=-4.614378268e-07 wa2=-1.676660667e-06 pa2=3.697372102e-13
+  b0=0.0
+  b1=0.0
+  keta=-2.697922500e-01 lketa=5.943737803e-08 wketa=2.159692167e-07 pketa=-4.762553166e-14
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=5.955905271e-01 lpclm=5.818458548e-09 wpclm=2.114164028e-08 ppclm=-4.662154515e-15
+  pdiblc1=3.970288360e+00 lpdiblc1=-8.353368741e-07 wpdiblc1=-3.035244236e-06 ppdiblc1=6.693320589e-13
+  pdiblc2=-4.935934427e-02 lpdiblc2=1.169089103e-08 wpdiblc2=4.247950796e-08 ppdiblc2=-9.367581094e-15
+  pdiblcb=-1.579302345e+01 lpdiblcb=3.385964893e-06 wpdiblcb=1.230309606e-05 ppdiblcb=-2.713078744e-12
+  drout=1.000001062e+00 ldrout=-2.024409511e-13
+  pscbe1=8.000000008e+08 lpscbe1=-1.559181213e-7
+  pscbe2=-3.775600725e-08 lpscbe2=9.914977023e-15 wpscbe2=3.602663270e-14 ppscbe2=-7.944593043e-21
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=8.401966736e+00 lbeta0=-1.109585119e-08 wbeta0=-4.031932164e-08 pbeta0=8.891216809e-15
* Gidl Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=1.000000320e+09 lbgidl=-6.090304565e-5
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-1.106e-8
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-1.559664757e+00 lkt1=2.248169204e-07 wkt1=8.168850748e-07 pkt1=-1.801394967e-13
+  kt2=8.267244544e-01 lkt2=-2.027588072e-07 wkt2=-7.367357200e-07 pkt2=1.624649610e-13
+  at=-4.251548531e+05 lat=1.024606843e-01 wat=3.722967500e-01 pat=-8.209887930e-8
+  ute=-8.843847175e+00 lute=1.931811385e-06 wute=7.019346662e-06 pute=-1.547906326e-12
+  ua1=-7.245475874e-09 lua1=1.755016736e-15 wua1=6.376952903e-15 pua1=-1.406245654e-21
+  ub1=6.808684109e-18 lub1=-1.599535167e-24 wub1=-5.812002834e-24 pub1=1.281662865e-30
+  uc1=-1.713684412e-10 luc1=3.282630327e-17 wuc1=1.192762380e-16 puc1=-2.630279601e-23
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.04e-6
+  sbref=1.04e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.126 pmos
* Model Flag Parameters
+  lmin=2.0e-05 lmax=0.0001 wmin=7.5e-07 wmax=7.9e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.126311+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+  k1=0.43165561
+  k2=0.026980026
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=3.2465718e-7
+  voff={-0.23051772+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.8768912+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+  eta0=0.08
+  etab=-0.07
+  u0=0.0095864
+  ua=-7.4757916e-10
+  ub=9.5046395e-19
+  uc=-1.0566299e-10
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=80156.0
+  a0=1.464
+  ags=0.11329
+  a1=0.0
+  a2=0.97
+  b0=-8.9873e-8
+  b1=3.3859e-9
+  keta=0.023361259
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=0.015
+  pdiblc1=0.39
+  pdiblc2=0.0012771588
+  pdiblcb=-0.225
+  drout=0.56
+  pscbe1=800000000.0
+  pscbe2=1.0060625e-8
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=0.0
+  alpha1=0.0
+  beta0=30.0
* Gidl Induced Drain Leakage Model Parameters
+  agidl=9.43573999999999e-11
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-0.43825
+  kt2=-0.058546
+  at=70990.0
+  ute=-0.08298
+  ua1=2.0902e-9
+  ub1=-1.2289e-18
+  uc1=-2.9789e-11
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.127 pmos
* Model Flag Parameters
+  lmin=8.0e-06 lmax=2.0e-05 wmin=7.5e-07 wmax=7.9e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.151793231e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=5.102439717e-7
+  k1=4.210498003e-01 lk1=2.123656422e-7
+  k2=3.098838670e-02 lk2=-8.026149068e-8
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=-6.144535039e-06 lcit=1.295359998e-10 wcit=1.694065895e-27 pcit=6.776263578e-32
+  voff={-2.428791561e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=2.475194627e-7
+  nfactor={1.918471956e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-8.325930941e-7
+  eta0=0.08
+  etab=-0.07
+  u0=9.965711908e-03 lu0=-7.595159576e-09 wu0=2.775557562e-23
+  ua=-7.615294670e-10 lua=2.793342514e-16
+  ub=9.271909546e-19 lub=4.660072882e-25
+  uc=-1.283201274e-10 luc=4.536756436e-16
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=2.656289816e+04 lvsat=1.073122547e+0
+  a0=1.605375760e+00 la0=-2.830840351e-6
+  ags=2.825339191e-02 lags=1.702732223e-6
+  a1=0.0
+  a2=1.083666533e+00 la2=-2.276004104e-6
+  b0=-1.499644844e-07 lb0=1.203243040e-12
+  b1=5.649803031e-09 lb1=-4.533130761e-14
+  keta=4.023168533e-02 lketa=-3.378053190e-7
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-6.921953293e-02 lpclm=1.686371502e-6
+  pdiblc1=0.39
+  pdiblc2=1.917610060e-03 lpdiblc2=-1.282408862e-08 ppdiblc2=2.775557562e-29
+  pdiblcb=-2.717239457e-01 lpdiblcb=9.355778616e-7
+  drout=0.56
+  pscbe1=8.000325955e+08 lpscbe1=-6.526776473e-1
+  pscbe2=1.315981805e-08 lpscbe2=-6.205675405e-14
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=-6.686266667e-11 lalpha0=1.338825943e-15
+  alpha1=-6.686266667e-11 lalpha1=1.338825943e-15
+  beta0=4.586076776e+01 lbeta0=-3.175884006e-4
* Gidl Induced Drain Leakage Model Parameters
+  agidl=-8.562847058e-09 lagidl=1.733477066e-13 wagidl=9.926167351e-30 pagidl=6.617444900e-35
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=-4.251725813e-01 legidl=1.051580369e-05 wegidl=4.440892099e-22 pegidl=1.065814104e-26
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.365640579e-01 lkt1=-3.375849616e-8
+  kt2=-6.268314622e-02 lkt2=8.284023011e-8
+  at=1.184558071e+05 lat=-9.504325371e-1
+  ute=-5.002598587e-02 lute=-6.598553610e-7
+  ua1=2.269041386e-09 lua1=-3.581034063e-15
+  ub1=-1.571912915e-18 lub1=6.868325966e-24
+  uc1=-4.384869988e-11 luc1=2.815246818e-16
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.128 pmos
* Model Flag Parameters
+  lmin=4.0e-06 lmax=8.0e-06 wmin=7.5e-07 wmax=7.9e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.090414346e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=1.776925644e-8
+  k1=4.556728822e-01 lk1=-6.543334786e-8
+  k2=1.885398624e-02 lk2=1.709911408e-8
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.057269452e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-5.057204472e-8
+  nfactor={2.150233085e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-2.692133146e-6
+  eta0=0.08
+  etab=-0.07
+  u0=8.535573484e-03 lu0=3.879584672e-9
+  ua=-8.237874492e-10 lua=7.788624164e-16
+  ub=1.048518672e-18 lub=-5.074680762e-25
+  uc=-7.083802061e-11 luc=-7.533189791e-18
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=2.678104074e+05 lvsat=-8.625316685e-1
+  a0=1.347035279e+00 la0=-7.580403376e-7
+  ags=2.084960866e-01 lags=2.565513575e-7
+  a1=0.0
+  a2=0.8
+  b0=0.0
+  b1=0.0
+  keta=-8.364571240e-04 lketa=-8.294256640e-9
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=2.407132755e-01 lpclm=-8.003805848e-7
+  pdiblc1=0.39
+  pdiblc2=-1.397670217e-03 lpdiblc2=1.377612899e-08 wpdiblc2=-1.734723476e-24 ppdiblc2=6.938893904e-30
+  pdiblcb=-2.494013897e-01 lpdiblcb=7.564723865e-7
+  drout=0.56
+  pscbe1=1.227212561e+09 lpscbe1=-3.428139670e+3
+  pscbe2=-1.711599940e-08 lpscbe2=1.808618728e-13 wpscbe2=-2.646977960e-29 ppscbe2=1.058791184e-34
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=3.429576331e+00 lbeta0=2.285911254e-5
* Gidl Induced Drain Leakage Model Parameters
+  agidl=2.613220901e-08 lagidl=-1.050287696e-13
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=1.675517744e+00 legidl=-6.339127153e-06 pegidl=-1.421085472e-26
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.061103840e-01 lkt1=-2.781041573e-7
+  kt2=-4.839276194e-02 lkt2=-3.181895402e-8
+  at=-9.120917488e+04 lat=7.318186388e-1
+  ute=-1.647219648e-01 lute=2.604101198e-7
+  ua1=5.703275549e-10 lua1=1.004863033e-14
+  ub1=8.239234094e-19 lub1=-1.235471470e-23 pub1=-1.232595164e-44
+  uc1=-1.164852119e-11 luc1=2.316590399e-17
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.129 pmos
* Model Flag Parameters
+  lmin=2.0e-06 lmax=4.0e-06 wmin=7.5e-07 wmax=7.9e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.085843201e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-6.228379991e-10
+  k1=4.428072554e-01 lk1=-1.366824095e-8
+  k2=2.193345702e-02 lk2=4.708801823e-9
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=8.622137339e-01 ldsub=-1.215963003e-6
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.337857314e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=6.232304277e-8
+  nfactor={7.881674337e-01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=2.788165241e-6
+  eta0=1.604349200e-01 leta0=-3.236315093e-7
+  etab=-1.403185835e-01 letab=2.829282271e-7
+  u0=8.638994592e-03 lu0=3.463467775e-9
+  ua=-8.215637429e-10 lua=7.699152898e-16
+  ub=1.011504174e-18 lub=-3.585395030e-25
+  uc=-7.560382119e-11 luc=1.164210416e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=53438.0
+  a0=1.154071298e+00 la0=1.835409954e-8
+  ags=1.482758150e-01 lags=4.988488244e-7
+  a1=0.0
+  a2=0.8
+  b0=0.0
+  b1=0.0
+  keta=6.578345336e-03 lketa=-3.812786263e-08 pketa=-2.775557562e-29
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-5.559724103e-01 lpclm=2.405100206e-06 ppclm=-3.552713679e-27
+  pdiblc1=0.39
+  pdiblc2=3.641230659e-03 lpdiblc2=-6.497989463e-9
+  pdiblcb=-9.820554637e-02 lpdiblcb=1.481328872e-07 ppdiblcb=-4.440892099e-28
+  drout=0.56
+  pscbe1=-4.676991234e+07 lpscbe1=1.697754289e+3
+  pscbe2=4.653609693e-08 lpscbe2=-7.524360986e-14 ppscbe2=-2.117582368e-34
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=1.147359093e+01 lbeta0=-9.506141085e-6
* Gidl Induced Drain Leakage Model Parameters
+  agidl=3.821637237e-11 lagidl=-3.906838872e-17
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.816142056e-01 lkt1=2.568697892e-8
+  kt2=-6.028632264e-02 lkt2=1.603502535e-8
+  at=1.022950518e+05 lat=-4.674948746e-2
+  ute=-1.327375183e-01 lute=1.317200597e-7
+  ua1=3.323674104e-09 lua1=-1.029514575e-15
+  ub1=-2.842323112e-18 lub1=2.396501504e-24
+  uc1=1.818504214e-11 luc1=-9.687003470e-17 wuc1=2.584939414e-32 puc1=1.033975766e-37
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.130 pmos
* Model Flag Parameters
+  lmin=1.0e-06 lmax=2.0e-06 wmin=7.5e-07 wmax=7.9e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.101264296e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=3.058205737e-8
+  k1=3.540326720e-01 lk1=1.659689040e-7
+  k2=5.577749960e-02 lk2=-6.377529522e-8
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=-2.663045674e-01 ldsub=1.067616350e-06 pdsub=8.881784197e-28
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.021762939e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-1.639286090e-9
+  nfactor={2.430472285e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-5.350714714e-7
+  eta0=-2.241626400e-01 leta0=4.546093453e-07 weta0=-5.204170428e-23 peta0=4.683753385e-29
+  etab=8.442995791e-01 letab=-1.709466317e-06 wetab=-6.800116026e-22 petab=-1.066854938e-27
+  u0=1.250070846e-02 lu0=-4.350787479e-9
+  ua=2.633023699e-11 lua=-9.458151364e-16
+  ub=5.976931819e-19 lub=4.788153150e-25
+  uc=-7.509174596e-11 luc=1.060590969e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=5.963848416e+04 lvsat=-1.254680371e-2
+  a0=1.369865781e+00 la0=-4.183103528e-7
+  ags=1.727992847e-01 lags=4.492250930e-7
+  a1=0.0
+  a2=5.953062352e-01 la2=4.142019269e-7
+  b0=0.0
+  b1=0.0
+  keta=-1.079934288e-02 lketa=-2.963762975e-9
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=4.550220723e-01 lpclm=3.593326501e-7
+  pdiblc1=7.492555200e-01 lpdiblc1=-7.269607298e-7
+  pdiblc2=0.00043
+  pdiblcb=-0.025
+  drout=1.096512000e-01 ldrout=9.112898038e-7
+  pscbe1=7.983183467e+08 lpscbe1=-1.229870506e+1
+  pscbe2=9.530520115e-09 lpscbe2=-3.620850560e-16
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=5.862313582e+00 lbeta0=1.848390856e-6
* Gidl Induced Drain Leakage Model Parameters
+  agidl=2.315918186e-11 lagidl=-8.599862589e-18
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.585366557e-01 lkt1=-2.101090483e-8
+  kt2=-5.625426130e-02 lkt2=7.876068592e-9
+  at=9.703221664e+04 lat=-3.610003518e-2
+  ute=9.359355551e-01 lute=-2.030761278e-06 wute=-8.881784197e-22 pute=1.332267630e-27
+  ua1=6.136533540e-09 lua1=-6.721391901e-15 pua1=1.323488980e-35
+  ub1=-4.270929418e-18 lub1=5.287314936e-24 wub1=-6.162975822e-39 pub1=-6.162975822e-45
+  uc1=-1.285649500e-10 luc1=2.000815094e-16 wuc1=-1.033975766e-31 puc1=-1.033975766e-37
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=2.75e-6
+  sbref=2.74e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.131 pmos
* Model Flag Parameters
+  lmin=5.0e-07 lmax=1.0e-06 wmin=7.5e-07 wmax=7.9e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.092582479e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=2.169604366e-8
+  k1=5.229315034e-01 lk1=-6.902427879e-9
+  k2=-6.829846957e-03 lk2=3.045761312e-10
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=1.255329254e+00 ldsub=-4.898062988e-7
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={2.670066454e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-4.818574081e-7
+  nfactor={1.728101006e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.838195797e-7
+  eta0=-2.358444013e-02 leta0=2.493135462e-7
+  etab=-1.689932780e+00 letab=8.843711865e-7
+  u0=1.006938082e-02 lu0=-1.862275006e-9
+  ua=-5.806459616e-10 lua=-3.245628577e-16
+  ub=8.868137281e-19 lub=1.828946535e-25
+  uc=-9.986617302e-11 luc=3.596303128e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=-5.927833243e+04 lvsat=1.091669364e-1
+  a0=1.185060244e+00 la0=-2.291581900e-7
+  ags=-5.662276608e-02 lags=6.840431505e-7
+  a1=0.0
+  a2=1.050779681e+00 la2=-5.198425436e-8
+  b0=-9.183315919e-17 lb0=9.399307509e-23
+  b1=-3.817924830e-20 lb1=3.907722422e-26
+  keta=1.192995869e-02 lketa=-2.622765772e-8
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=1.588106337e+00 lpclm=-8.004017569e-7
+  pdiblc1=6.353741327e-02 lpdiblc1=-2.511453323e-8
+  pdiblc2=7.762209763e-04 lpdiblc2=-3.543640937e-10
+  pdiblcb=-1.404746093e-02 lpdiblcb=-1.121014279e-8
+  drout=1.039619329e+00 ldrout=-4.055117553e-8
+  pscbe1=8.256802058e+08 lpscbe1=-4.030411509e+1
+  pscbe2=3.429057487e-09 lpscbe2=5.882883972e-15
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=6.559046608e+00 lbeta0=1.135270669e-6
* Gidl Induced Drain Leakage Model Parameters
+  agidl=3.020804646e-11 lagidl=-1.581451648e-17
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.216831793e-01 lkt1=-5.873117501e-8
+  kt2=-6.301890653e-02 lkt2=1.479981827e-8
+  at=8.604123040e+04 lat=-2.485054094e-2
+  ute=-1.934483867e+00 lute=9.071704088e-7
+  ua1=-3.495144579e-09 lua1=3.136823287e-15 pua1=8.271806126e-37
+  ub1=4.257545597e-18 lub1=-3.441749811e-24 wub1=-3.081487911e-39
+  uc1=3.311138654e-10 luc1=-2.704089518e-16 wuc1=4.135903063e-31 puc1=-2.067951531e-37
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.75e-6
+  sbref=1.74e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.132 pmos
* Model Flag Parameters
+  lmin=2.5e-07 lmax=5.0e-07 wmin=7.5e-07 wmax=7.9e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.045892418e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-2.747137143e-9
+  k1=4.352213524e-01 lk1=3.901559036e-8
+  k2=1.408936088e-02 lk2=-1.064704755e-08 pk2=6.938893904e-30
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=-1.888704683e-01 ldsub=2.662611400e-7
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-8.564575735e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=1.062985797e-7
+  nfactor={1.710086311e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.932506331e-7
+  eta0=4.117672797e-01 leta0=2.139821381e-8
+  etab=-1.291129272e-03 letab=3.335097045e-10
+  u0=7.485205816e-03 lu0=-5.094077095e-10
+  ua=-1.063421140e-09 lua=-7.182039643e-17
+  ub=1.148080500e-18 lub=4.611627323e-26
+  uc=-6.419271038e-11 luc=1.728726011e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=1.425608788e+05 lvsat=3.500072552e-3
+  a0=8.919849864e-01 la0=-7.572743094e-8
+  ags=9.698322768e-01 lags=1.466734064e-7
+  a1=0.0
+  a2=1.121568012e+00 la2=-8.904336116e-8
+  b0=1.836663184e-16 lb0=-5.023641140e-23
+  b1=7.635849659e-20 lb1=-2.088557599e-26
+  keta=-4.524308758e-02 lketa=3.703575468e-9
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-5.731343976e-01 lpclm=3.310509927e-07 wpclm=2.220446049e-22 ppclm=5.551115123e-29
+  pdiblc1=-4.101030779e-01 lpdiblc1=2.228457367e-07 wpdiblc1=4.440892099e-22
+  pdiblc2=-9.175377595e-03 lpdiblc2=4.855496791e-09 wpdiblc2=9.107298249e-24 ppdiblc2=-2.059984128e-30
+  pdiblcb=2.408596814e-01 lpdiblcb=-1.446591300e-07 ppdiblcb=1.665334537e-28
+  drout=1.436421824e+00 ldrout=-2.482852179e-7
+  pscbe1=6.925891618e+08 lpscbe1=2.937170827e+1
+  pscbe2=2.103542680e-08 lpscbe2=-3.334402489e-15
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=8.528056950e+00 lbeta0=1.044543745e-7
* Gidl Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=7.372237654e+08 lbgidl=1.375686143e+2
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.00074326333
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.5407449e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-5.460023937e-01 lkt1=6.352420121e-9
+  kt2=-1.498550792e-02 lkt2=-1.034662657e-8
+  at=6.500485322e+03 lat=1.679062992e-2
+  ute=4.908242408e-01 lute=-3.625268917e-07 pute=-4.440892099e-28
+  ua1=4.905387581e-09 lua1=-1.261023309e-15
+  ub1=-4.666106948e-18 lub1=1.229960769e-24
+  uc1=-2.811617509e-10 luc1=5.012957887e-17
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.1e-6
+  sbref=1.1e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.133 pmos
* Model Flag Parameters
+  lmin=1.8e-07 lmax=2.5e-07 wmin=7.5e-07 wmax=7.9e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.029269231e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-7.293911197e-9
+  k1=-9.625672899e-01 lk1=4.213387398e-7
+  k2=5.727293397e-01 lk2=-1.634462546e-07 wk2=-4.440892099e-22 pk2=1.110223025e-28
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=2.137145701e+00 ldsub=-3.699508026e-7
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-1.089170690e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=1.699502713e-7
+  nfactor={-2.921819978e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.460169641e-6
+  eta0=1.215531322e+00 leta0=-1.984473271e-7
+  etab=7.331369097e-02 letab=-2.007240073e-08 wetab=-6.158268340e-23 petab=-2.428612866e-29
+  u0=1.425792013e-02 lu0=-2.361880528e-9
+  ua=1.625481428e-09 lua=-8.072890268e-16
+  ub=-7.962308851e-19 lub=5.779243232e-25
+  uc=-1.092267674e-12 luc=2.802702628e-20
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=2.884433928e+05 lvsat=-3.640171267e-2
+  a0=-8.336933221e-01 la0=3.962801000e-7
+  ags=2.250598985e+00 lags=-2.036419037e-7
+  a1=0.0
+  a2=1.211177822e+00 la2=-1.135534364e-7
+  b0=0.0
+  b1=0.0
+  keta=-1.231216453e-01 lketa=2.500491856e-8
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=6.814682513e-01 lpclm=-1.210792385e-8
+  pdiblc1=1.051165451e+00 lpdiblc1=-1.768404313e-7
+  pdiblc2=2.288324307e-02 lpdiblc2=-3.913177133e-09 wpdiblc2=5.551115123e-23
+  pdiblcb=1.496831658e-01 lpdiblcb=-1.197205294e-7
+  drout=-8.416449981e-01 ldrout=3.748116193e-7
+  pscbe1=7.998956541e+08 lpscbe1=2.123650263e-2
+  pscbe2=1.360976700e-08 lpscbe2=-1.303336022e-15
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=1.053315297e+01 lbeta0=-4.439794884e-7
* Gidl Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=1.938486425e+09 lbgidl=-1.910007483e+2
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.00074326333
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.5407449e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.721835984e-01 lkt1=-1.383849677e-8
+  kt2=6.325147130e-02 lkt2=-3.174600512e-8
+  at=1.504888693e+05 lat=-2.259307287e-2
+  ute=-3.018056026e+00 lute=5.972220390e-7
+  ua1=-9.203434720e-10 lua1=3.324306487e-16 pua1=-4.135903063e-37
+  ub1=6.315712371e-19 lub1=-2.190601681e-25
+  uc1=-3.170369254e-10 luc1=5.994215660e-17
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.1e-6
+  sbref=1.1e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.134 pmos
* Model Flag Parameters
+  lmin=1.5e-07 lmax=1.8e-07 wmin=7.5e-07 wmax=7.9e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-2.026e-8
+  vth0={-1.026501304e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-8.513553884e-09 wvth0=-1.059331889e-08 pvth0=2.336038682e-15
+  k1=3.187794420e-01 lk1=1.739705304e-07 wk1=6.321316583e-07 pk1=-1.393976733e-13
+  k2=-5.917828312e-02 lk2=-3.775063066e-08 wk2=-1.214458214e-07 pk2=2.678123254e-14
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=2.831294506e+00 ldsub=-5.539264412e-07 wdsub=-2.012724951e-06 pdsub=4.438461061e-13
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-1.146439752e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=1.967751696e-07 wvoff=7.149938099e-07 pvoff=-1.576704350e-13
+  nfactor={2.909554634e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=2.962026982e-07 wnfactor=3.893404182e-06 pnfactor=-8.585734902e-13
+  eta0=5.710310891e+00 leta0=-1.206212398e-06 weta0=-4.382841334e-06 peta0=9.665041709e-13
+  etab=5.108517495e-01 letab=-1.182349385e-07 wetab=-4.296136144e-07 petab=9.473839425e-14
+  u0=4.110143461e-03 lu0=-3.213804012e-10 wu0=-7.097003082e-10 pu0=1.565031120e-16
+  ua=-3.062213224e-09 lua=1.590086471e-16 wua=5.777671626e-16 pua=-1.274092147e-22
+  ub=2.189775517e-18 lub=-3.227586245e-26 wub=-1.172769596e-25 pub=2.586191513e-32
+  uc=-2.722694536e-10 luc=5.983036117e-17 wuc=2.173970365e-16 puc=-4.794039450e-23
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=-1.120963484e+06 lvsat=2.713600613e-01 wvsat=9.064222450e-01 pvsat=-1.998842335e-7
+  a0=-4.066283983e+00 la0=1.142232220e-06 wa0=4.150365918e-06 pa0=-9.152386923e-13
+  ags=1.250000065e+00 lags=-1.235200386e-14
+  a1=0.0
+  a2=2.745729274e+00 la2=-4.614378268e-07 wa2=-1.676660667e-06 pa2=3.697372102e-13
+  b0=0.0
+  b1=0.0
+  keta=-2.697922500e-01 lketa=5.943737803e-08 wketa=2.159692167e-07 pketa=-4.762553166e-14
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=5.955905271e-01 lpclm=5.818458548e-09 wpclm=2.114164028e-08 ppclm=-4.662154515e-15
+  pdiblc1=3.970288360e+00 lpdiblc1=-8.353368741e-07 wpdiblc1=-3.035244236e-06 ppdiblc1=6.693320589e-13
+  pdiblc2=-4.935934427e-02 lpdiblc2=1.169089103e-08 wpdiblc2=4.247950796e-08 ppdiblc2=-9.367581094e-15
+  pdiblcb=-1.579302345e+01 lpdiblcb=3.385964893e-06 wpdiblcb=1.230309606e-05 ppdiblcb=-2.713078744e-12
+  drout=1.000001062e+00 ldrout=-2.024409795e-13 wdrout=-8.526512829e-20 pdrout=2.131628207e-26
+  pscbe1=8.000000008e+08 lpscbe1=-1.559181213e-7
+  pscbe2=-3.775600725e-08 lpscbe2=9.914977023e-15 wpscbe2=3.602663270e-14 ppscbe2=-7.944593043e-21
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=8.401966736e+00 lbeta0=-1.109585119e-08 wbeta0=-4.031932164e-08 pbeta0=8.891216808e-15
* Gidl Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=1.000000320e+09 lbgidl=-6.090304565e-5
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-1.106e-8
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-1.559664757e+00 lkt1=2.248169204e-07 wkt1=8.168850748e-07 pkt1=-1.801394967e-13
+  kt2=8.267244544e-01 lkt2=-2.027588072e-07 wkt2=-7.367357200e-07 pkt2=1.624649610e-13
+  at=-4.251548531e+05 lat=1.024606843e-01 wat=3.722967500e-01 pat=-8.209887930e-8
+  ute=-8.843847175e+00 lute=1.931811385e-06 wute=7.019346662e-06 pute=-1.547906326e-12
+  ua1=-7.245475874e-09 lua1=1.755016736e-15 wua1=6.376952903e-15 pua1=-1.406245654e-21
+  ub1=6.808684109e-18 lub1=-1.599535167e-24 wub1=-5.812002834e-24 pub1=1.281662865e-30
+  uc1=-1.713684412e-10 luc1=3.282630327e-17 wuc1=1.192762380e-16 puc1=-2.630279601e-23
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.04e-6
+  sbref=1.04e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.135 pmos
* Model Flag Parameters
+  lmin=2.0e-05 lmax=0.0001 wmin=7.0e-07 wmax=7.5e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.126311+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+  k1=0.43165561
+  k2=0.026980026
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=3.2465718e-7
+  voff={-0.23051772+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.8768912+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+  eta0=0.08
+  etab=-0.07
+  u0=0.0095864
+  ua=-7.4757916e-10
+  ub=9.5046395e-19
+  uc=-1.0566299e-10
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=80156.0
+  a0=1.464
+  ags=0.11329
+  a1=0.0
+  a2=0.97
+  b0=-8.9873e-8
+  b1=3.3859e-9
+  keta=0.023361259
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=0.015
+  pdiblc1=0.39
+  pdiblc2=0.0012771588
+  pdiblcb=-0.225
+  drout=0.56
+  pscbe1=800000000.0
+  pscbe2=1.0060625e-8
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=0.0
+  alpha1=0.0
+  beta0=30.0
* Gidl Induced Drain Leakage Model Parameters
+  agidl=9.43573999999999e-11
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-0.43825
+  kt2=-0.058546
+  at=70990.0
+  ute=-0.08298
+  ua1=2.0902e-9
+  ub1=-1.2289e-18
+  uc1=-2.9789e-11
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.136 pmos
* Model Flag Parameters
+  lmin=8.0e-06 lmax=2.0e-05 wmin=7.0e-07 wmax=7.5e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-9.888904645e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-2.751642841e-06 wvth0=-1.191262322e-07 pvth0=2.385326493e-12
+  k1=4.756564958e-01 lk1=-8.810526164e-07 wk1=-3.993234740e-08 pk1=7.995861568e-13
+  k2=6.836158540e-02 lk2=-8.286044823e-07 wk2=-2.732997376e-08 pk2=5.472422762e-13
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=-6.144535039e-06 lcit=1.295359998e-10 wcit=-3.388131789e-27 pcit=-2.710505431e-32
+  voff={-1.644528585e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-1.322851075e-06 wvoff=-5.735095548e-08 pvoff=1.148368004e-12
+  nfactor={-1.060811764e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=5.882315405e-05 wnfactor=2.178666764e-06 pnfactor=-4.362457752e-11
+  eta0=0.08
+  etab=-0.07
+  u0=8.128341260e-04 lu0=1.756776717e-07 wu0=6.693243241e-09 pu0=-1.340222899e-13
+  ua=1.283819901e-09 lua=-4.067575973e-14 wua=-1.495706723e-15 pua=2.994931349e-20
+  ub=-4.692614964e-18 lub=1.129943035e-22 wub=4.109606714e-24 pub=-8.228879223e-29
+  uc=-4.507886468e-10 luc=6.910630491e-15 wuc=2.358121991e-16 puc=-4.721790285e-21
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=-8.776011276e+05 lvsat=1.917766900e+01 wvsat=6.611898354e-01 pvsat=-1.323934789e-5
+  a0=1.317149436e+00 la0=2.940465199e-06 wa0=2.107718399e-07 pa0=-4.220394152e-12
+  ags=-1.122964394e+00 lags=2.475416459e-05 wags=8.418533331e-07 pags=-1.685686705e-11
+  a1=0.0
+  a2=1.083666533e+00 la2=-2.276004104e-6
+  b0=1.358995297e-07 lb0=-4.520760764e-12 wb0=-2.090443493e-13 pb0=4.185803709e-18
+  b1=8.336895610e-09 lb1=-9.913635962e-14 wb1=-1.964995565e-15 pb1=3.934612799e-20
+  keta=1.222295640e-01 lketa=-1.979691482e-06 wketa=-5.996275270e-08 pketa=1.200665378e-12
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-6.921953293e-02 lpclm=1.686371502e-06 wpclm=2.775557562e-23
+  pdiblc1=0.39
+  pdiblc2=2.026251140e-03 lpdiblc2=-1.499946546e-08 wpdiblc2=-7.944617972e-11 ppdiblc2=1.590792169e-15
+  pdiblcb=-9.083582647e-01 lpdiblcb=1.368323788e-05 wpdiblcb=4.655528517e-07 ppdiblcb=-9.322006837e-12
+  drout=0.56
+  pscbe1=8.004767243e+08 lpscbe1=-9.545697770e+00 wpscbe1=-3.247788906e-01 ppscbe1=6.503216611e-6
+  pscbe2=7.173623340e-08 lpscbe2=-1.234962778e-12 wpscbe2=-4.283529241e-14 ppscbe2=8.577133342e-19
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=-6.686266667e-11 lalpha0=1.338825943e-15
+  alpha1=-6.686266667e-11 lalpha1=1.338825943e-15
+  beta0=1.599172902e+01 lbeta0=2.804948942e-04 wbeta0=2.184239170e-05 pbeta0=-4.373615671e-10
* Gidl Induced Drain Leakage Model Parameters
+  agidl=-1.270808056e-07 lagidl=2.546494420e-12 wagidl=8.666886459e-14 pagidl=-1.735415743e-18
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=-7.580880078e+00 legidl=1.537982559e-04 wegidl=5.232768532e-06 pegidl=-1.047784454e-10
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-3.299115814e-01 lkt1=-2.169316491e-06 wkt1=-7.799196975e-08 pkt1=1.561673766e-12
+  kt2=-2.807034184e-02 lkt2=-6.102299507e-07 wkt2=-2.531137469e-08 pkt2=5.068228173e-13
+  at=6.811258234e+05 lat=-1.221706686e+01 wat=-4.114648282e-01 pat=8.238974216e-6
+  ute=-8.394121972e+00 lute=1.664183175e-04 wute=6.101803760e-06 pute=-1.221795896e-10
+  ua1=-1.825770657e-08 lua1=4.074367141e-13 wua1=1.501063603e-14 pua1=-3.005657707e-19
+  ub1=1.310277777e-17 lub1=-2.869706365e-22 wub1=-1.073119041e-23 pub1=2.148762058e-28
+  uc1=6.456217551e-10 luc1=-1.352410076e-14 wuc1=-5.041904386e-16 puc1=1.009566733e-20
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.137 pmos
* Model Flag Parameters
+  lmin=4.0e-06 lmax=8.0e-06 wmin=7.0e-07 wmax=7.5e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.826055678e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=3.965368993e-06 wvth0=5.379539081e-07 pvth0=-2.886769154e-12
+  k1=3.911231088e-01 lk1=-2.027972957e-07 wk1=4.720344188e-08 pk1=1.004504088e-13
+  k2=-1.481909608e-01 lk2=9.089092033e-07 wk2=1.221552925e-07 pk2=-6.521557476e-13
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-4.156687847e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=6.927849331e-07 wvoff=1.535245889e-07 pvoff=-5.435961439e-13
+  nfactor={2.084474039e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.169364817e-04 wnfactor=-1.367076974e-05 pnfactor=8.354369328e-11
+  eta0=0.08
+  etab=-0.07
+  u0=5.160227398e-02 lu0=-2.318324147e-07 wu0=-3.149347221e-08 pu0=1.723695852e-13
+  ua=-4.920767924e-09 lua=9.106874780e-15 wua=2.996007106e-15 pua=-6.090042257e-21
+  ub=1.641019926e-17 lub=-5.632454851e-23 wub=-1.123356689e-23 pub=4.081746804e-29
+  uc=4.219816178e-10 luc=-9.205918246e-17 wuc=-3.603852026e-16 puc=6.181149171e-23
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=3.052433313e+06 lvsat=-1.235504093e+01 wvsat=-2.036316761e+00 pvsat=8.404150236e-6
+  a0=3.770080004e+00 la0=-1.674067227e-05 wa0=-1.771904762e-06 pa0=1.168765122e-11
+  ags=2.439365090e+00 lags=-3.828257273e-06 wags=-1.631372038e-06 pags=2.987106177e-12
+  a1=0.0
+  a2=0.8
+  b0=-1.817310007e-06 lb0=1.115085502e-11 wb0=1.328947923e-12 pb0=-8.154308050e-18
+  b1=1.691847152e-08 lb1=-1.679908056e-13 wb1=-1.237200451e-14 pb1=1.228469724e-19
+  keta=-1.149748278e-01 lketa=-7.647730010e-08 wketa=8.346619462e-08 pketa=4.986035056e-14
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=9.119689207e+00 lpclm=-7.204102155e-05 wpclm=-6.492946487e-06 ppclm=5.209628600e-11
+  pdiblc1=0.39
+  pdiblc2=-2.360080879e-02 lpdiblc2=1.906197624e-07 wpdiblc2=1.623653355e-08 ppdiblc2=-1.293207975e-13
+  pdiblcb=-5.818810603e-01 lpdiblcb=1.106374150e-05 wpdiblcb=2.431330737e-07 ppdiblcb=-7.537417300e-12
+  drout=0.56
+  pscbe1=7.048171672e+09 lpscbe1=-5.013805106e+04 wpscbe1=-4.256704411e+03 ppscbe1=3.415765032e-2
+  pscbe2=-4.497359603e-07 lpscbe2=2.949079797e-12 wpscbe2=3.163628640e-13 ppscbe2=-2.024320258e-18
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=-1.270555759e-09 lalpha0=1.099668154e-14 walpha0=1.002249051e-15 palpha0=-8.041565304e-21
+  alpha1=-1.270555759e-09 lalpha1=1.099668154e-14 walpha1=1.002249051e-15 palpha1=-8.041565304e-21
+  beta0=3.793327977e+02 lbeta0=-2.634779437e-03 wbeta0=-2.748875005e-04 pbeta0=1.943456658e-9
* Gidl Induced Drain Leakage Model Parameters
+  agidl=3.815295249e-07 lagidl=-1.534350739e-12 wagidl=-2.598921060e-13 pagidl=1.045223135e-18
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=2.314264023e+01 legidl=-9.271252383e-05 wegidl=-1.569830560e-05 pegidl=6.316244653e-11
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-3.014696393e-01 lkt1=-2.397520983e-06 wkt1=-7.652084669e-08 pkt1=1.549870181e-12
+  kt2=-1.830001519e-01 lkt2=6.328524787e-07 wkt2=9.843461525e-08 pkt2=-4.860556079e-13
+  at=-1.637860103e+06 lat=6.389363097e+00 wat=1.131022517e+00 pat=-4.137203851e-6
+  ute=2.373027882e+01 lute=-9.133245478e-05 wute=-1.747374502e-05 pute=6.697929750e-11
+  ua1=4.875201832e-08 lua1=-1.302171537e-13 wua1=-3.523392137e-14 pua1=1.025724404e-19
+  ub1=-2.788007638e-17 lub1=4.185611345e-23 wub1=2.099043133e-23 pub1=-3.964286072e-29
+  uc1=-7.730163667e-09 luc1=5.367918108e-14 wuc1=5.644334007e-15 puc1=-3.923714153e-20
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.138 pmos
* Model Flag Parameters
+  lmin=2.0e-06 lmax=4.0e-06 wmin=7.0e-07 wmax=7.5e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-8.103091478e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-1.215074866e-07 wvth0=-2.014903380e-07 pvth0=8.839955872e-14
+  k1=1.225807115e+00 lk1=-3.561165090e-06 wk1=-5.725858736e-07 pk1=2.594185116e-12
+  k2=-2.330807718e-01 lk2=1.250465056e-06 wk2=1.864847652e-07 pk2=-9.109866673e-13
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=8.443064175e-01 ldsub=-1.143912557e-06 wdsub=1.309511903e-08 pdsub=-5.268847333e-14
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-3.893048602e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=5.867091554e-07 wvoff=1.137267844e-07 pvoff=-3.834688814e-13
+  nfactor={-1.941557006e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=4.505168257e-05 wnfactor=1.477442753e-05 pnfactor=-3.090612684e-11
+  eta0=1.604349200e-01 leta0=-3.236315093e-7
+  etab=-1.403357992e-01 letab=2.829974947e-07 wetab=1.258935134e-11 petab=-5.065350689e-17
+  u0=-3.869121542e-02 lu0=1.314652458e-07 wu0=3.461125734e-08 pu0=-9.360411620e-14
+  ua=-1.023266084e-08 lua=3.047938215e-14 wua=6.882071794e-15 pua=-2.172570125e-20
+  ub=6.362971760e-18 lub=-1.589932770e-23 wub=-3.913378405e-24 pub=1.136454327e-29
+  uc=7.174654981e-10 luc=-1.280944484e-15 wuc=-5.799493872e-16 puc=9.452323797e-22
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=-3.614778172e+05 lvsat=1.380898776e+00 wvsat=3.034163195e-01 pvsat=-1.009812610e-6
+  a0=-2.207241251e+00 la0=7.309199343e-06 wa0=2.458033750e-06 pa0=-5.331590983e-12
+  ags=2.772491850e+00 lags=-5.168599455e-06 wags=-1.919015708e-06 pags=4.144446238e-12
+  a1=0.0
+  a2=0.8
+  b0=1.367112853e-06 lb0=-1.661734049e-12 wb0=-9.997313503e-13 pb0=1.215179581e-18
+  b1=-1.977438415e-08 lb1=-2.035636690e-14 wb1=1.446045345e-14 pb1=1.488604113e-20
+  keta=-2.145978629e-01 lketa=3.243579738e-07 wketa=1.617399681e-07 pketa=-2.650757426e-13
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-1.638822495e+01 lpclm=3.059058122e-05 wpclm=1.157768298e-05 ppclm=-2.061125308e-11
+  pdiblc1=0.39
+  pdiblc2=4.755176576e-02 lpdiblc2=-9.566404433e-08 wpdiblc2=-3.211054483e-08 ppdiblc2=6.520463928e-14
+  pdiblcb=4.386559709e+00 lpdiblcb=-8.926879302e-06 wpdiblcb=-3.279583258e-06 ppdiblcb=6.636302314e-12
+  drout=0.56
+  pscbe1=-1.158438255e+10 lpscbe1=2.483040349e+04 wpscbe1=8.437133066e+03 ppscbe1=-1.691625864e-2
+  pscbe2=5.618995403e-07 lpscbe2=-1.121255872e-12 wpscbe2=-3.768708560e-13 ppscbe2=7.649194792e-19
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=2.841111517e-09 lalpha0=-5.546693978e-15 walpha0=-2.004498102e-15 palpha0=4.056141999e-21
+  alpha1=2.841111517e-09 lalpha1=-5.546693978e-15 walpha1=-2.004498102e-15 palpha1=4.056141999e-21
+  beta0=-5.777699435e+02 lbeta0=1.216142584e-03 wbeta0=4.308972979e-04 pbeta0=-8.962825945e-10
* Gidl Induced Drain Leakage Model Parameters
+  agidl=3.361923060e-10 lagidl=-6.117412458e-16 wagidl=-2.179014569e-16 pagidl=4.187796255e-22
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-1.109550467e+00 lkt1=8.538083898e-07 wkt1=4.591922059e-07 pkt1=-6.055820004e-13
+  kt2=-2.043323612e-02 lkt2=-2.123875818e-08 wkt2=-2.914344628e-08 pkt2=2.725727423e-14
+  at=-7.201323731e+05 lat=2.696867222e+00 wat=6.014181479e-01 pat=-2.006330078e-6
+  ute=-6.939730642e-01 lute=6.939011178e-06 wute=4.104158401e-07 pute=-4.977981391e-12
+  ua1=9.274082300e-09 lua1=2.862311143e-14 wua1=-4.351366902e-15 pua1=-2.168413512e-20
+  ub1=-1.561623263e-17 lub1=-7.487707165e-24 wub1=9.341202360e-24 pub1=7.228045041e-30
+  uc1=1.221739784e-08 luc1=-2.658023158e-14 wuc1=-8.920942740e-15 puc1=1.936654077e-20
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.139 pmos
* Model Flag Parameters
+  lmin=1.0e-06 lmax=2.0e-06 wmin=7.0e-07 wmax=7.5e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-8.717528304e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=2.825034048e-09 wvth0=-1.678353087e-07 pvth0=2.029793396e-14
+  k1=-1.722928233e+00 lk1=2.405659863e-06 wk1=1.518823355e-06 pk1=-1.637823287e-12
+  k2=8.533724819e-01 lk2=-9.479948323e-07 wk2=-5.832588779e-07 pk2=6.466049893e-13
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=-7.437436148e+00 ldsub=1.561435916e-05 wdsub=5.244047733e-06 pdsub=-1.063762571e-11
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-1.604132786e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=1.235424622e-07 wvoff=-3.054012376e-08 pvoff=-9.154190742e-14
+  nfactor={1.372368471e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=2.986873184e-06 wnfactor=7.737616924e-07 pnfactor=-2.575499512e-12
+  eta0=3.541233154e+00 leta0=-7.164744352e-06 weta0=-2.753528513e-06 peta0=5.571820017e-12
+  etab=1.234464833e+01 letab=-2.498061760e-05 wetab=-8.409883035e-06 petab=1.701754134e-11
+  u0=2.669302544e-02 lu0=-8.410732975e-10 wu0=-1.037844402e-08 pu0=-2.566555709e-15
+  ua=4.906545040e-09 lua=-1.551037253e-16 wua=-3.568764440e-15 pua=-5.782251150e-22
+  ub=-9.740529492e-19 lub=-1.052711464e-24 wub=1.149373937e-24 pub=1.119962651e-30
+  uc=5.319927074e-10 luc=-9.056365829e-16 wuc=-4.439438624e-16 puc=6.700224801e-22
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=6.627622624e+05 lvsat=-6.916715100e-01 wvsat=-4.410475315e-01 pvsat=4.966248822e-7
+  a0=5.987898701e+00 la0=-9.273830252e-06 wa0=-3.377038169e-06 pa0=6.475793748e-12
+  ags=-8.459669049e-01 lags=2.153424205e-06 wags=7.449951890e-07 pags=-1.246233093e-12
+  a1=0.0
+  a2=-2.193736375e+00 la2=6.057885430e-06 wa2=2.039548768e-06 pa2=-4.127067723e-12
+  b0=-2.810613383e-07 lb0=1.673379391e-12 wb0=2.055322870e-13 pb0=-1.223695494e-18
+  b1=3.753279024e-07 lb1=-8.198537458e-13 wb1=-2.744667858e-13 pb1=5.995360884e-19
+  keta=8.066116310e-02 lketa=-2.731045704e-07 wketa=-6.688250713e-08 pketa=1.975464085e-13
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-5.879381478e+00 lpclm=9.325726280e-06 wpclm=4.632171953e-06 ppclm=-6.556872602e-12
+  pdiblc1=5.565324206e+00 lpdiblc1=-1.047237204e-05 wpdiblc1=-3.521856180e-06 ppdiblc1=7.126546418e-12
+  pdiblc2=1.177911272e-04 lpdiblc2=3.195520255e-10 wpdiblc2=2.283096068e-10 ppdiblc2=-2.336794488e-16
+  pdiblcb=-2.814182070e+00 lpdiblcb=5.643965702e-06 wpdiblcb=2.039650751e-06 ppdiblcb=-4.127274087e-12
+  drout=-3.566972320e+00 ldrout=8.351011029e-06 wdrout=2.688611835e-06 pdrout=-5.440459820e-12
+  pscbe1=7.754050805e+08 lpscbe1=-1.798739729e+02 wpscbe1=1.675582996e+01 ppscbe1=1.225431013e-4
+  pscbe2=6.273955912e-09 lpscbe2=3.063610230e-15 wpscbe2=2.381434218e-15 ppscbe2=-2.505115043e-21
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=2.247271270e+01 lbeta0=1.539564340e-06 wbeta0=-1.214671978e-05 pbeta0=2.258361835e-13
* Gidl Induced Drain Leakage Model Parameters
+  agidl=-5.838036797e-12 lagidl=8.036399338e-17 wagidl=2.120485408e-17 pagidl=-6.505677688e-23
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-9.010568288e-01 lkt1=4.319173427e-07 wkt1=3.236026120e-07 pkt1=-3.312137455e-13
+  kt2=-1.288452720e-02 lkt2=-3.651372165e-08 wkt2=-3.171507219e-08 pkt2=3.246101069e-14
+  at=1.036991479e+06 lat=-8.587080362e-01 wat=-6.873658899e-01 pat=6.015501981e-7
+  ute=6.607555321e+00 lute=-7.835777541e-06 wute=-4.147496730e-06 pute=4.245045853e-12
+  ua1=4.782992954e-08 lua1=-4.939541657e-14 wua1=-3.048921308e-14 pua1=3.120631937e-20
+  ub1=-4.056123588e-17 lub1=4.298900582e-23 wub1=2.653808499e-23 pub1=-2.757019090e-29
+  uc1=-1.926575420e-09 luc1=2.040381186e-15 wuc1=1.314834713e-15 puc1=-1.345759625e-21
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=2.75e-6
+  sbref=2.74e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.140 pmos
* Model Flag Parameters
+  lmin=5.0e-07 lmax=1.0e-06 wmin=7.0e-07 wmax=7.5e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-6.782773743e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-1.952009647e-07 wvth0=-3.029697225e-07 pvth0=1.586107091e-13
+  k1=7.506913696e-01 lk1=-1.261392730e-07 wk1=-1.665544129e-07 pk1=8.719456623e-14
+  k2=-1.425600885e-01 lk2=7.136207217e-08 wk2=9.925572517e-08 pk2=-5.196235724e-14
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=1.566922168e+01 ldsub=-8.035767261e-06 wdsub=-1.054047594e-05 pdsub=5.518149965e-12
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={6.028607049e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-6.576837253e-07 wvoff=-2.456006698e-07 pvoff=1.285768626e-13
+  nfactor={6.606009485e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-2.369863067e-06 wnfactor=-3.567077889e-06 pnfactor=1.867436617e-12
+  eta0=-7.554376028e+00 leta0=4.191833558e-06 weta0=5.507057026e-06 peta0=-2.883054494e-12
+  etab=-2.469056143e+01 letab=1.292566030e-05 wetab=1.681971571e-05 petab=-8.805457570e-12
+  u0=4.614104972e-02 lu0=-2.074651511e-08 wu0=-2.637820146e-08 pu0=1.380951603e-14
+  ua=1.099077177e-08 lua=-6.382431469e-15 wua=-8.461853788e-15 pua=4.429949695e-21
+  ub=-5.393667030e-18 lub=3.470851940e-24 wub=4.592739725e-24 pub=-2.404391101e-30
+  uc=-6.896249989e-10 luc=3.447135718e-16 wuc=4.312741161e-16 puc=-2.257806253e-22
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=-1.829092460e+05 lvsat=1.738901923e-01 wvsat=9.040782546e-02 pvsat=-4.733030479e-8
+  a0=-7.072681445e+00 la0=4.093934739e-06 wa0=6.038655281e-06 pa0=-3.161356813e-12
+  ags=1.266320318e+00 lags=-8.544012715e-09 wags=-9.674312347e-07 pags=5.064696000e-13
+  a1=0.0
+  a2=6.628864902e+00 la2=-2.972223429e-06 wa2=-4.079097536e-06 pa2=2.135489142e-12
+  b0=2.771414980e-06 lb0=-1.450891170e-12 wb0=-2.026658175e-12 pb0=1.060996088e-18
+  b1=-8.713962622e-07 lb1=4.561933712e-13 wb1=6.372276875e-13 pb1=-3.336014389e-19
+  keta=-3.411283420e-01 lketa=1.586054239e-07 wketa=2.581816497e-07 pketa=-1.351632572e-13
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=6.554116152e+00 lpclm=-3.400207215e-06 wpclm=-3.631503929e-06 ppclm=1.901164937e-12
+  pdiblc1=-9.568599959e+00 lpdiblc1=5.017502024e-06 wpdiblc1=7.043712361e-06 ppdiblc1=-3.687524295e-12
+  pdiblc2=7.762209763e-04 lpdiblc2=-3.543640937e-10
+  pdiblcb=5.564316679e+00 lpdiblcb=-2.931595337e-06 wpdiblcb=-4.079301501e-06 ppdiblcb=2.135595922e-12
+  drout=8.392866369e+00 ldrout=-3.890123066e-06 wdrout=-5.377223670e-06 pdrout=2.815084136e-12
+  pscbe1=4.436252978e+08 lpscbe1=1.597092704e+02 wpscbe1=2.793860567e+02 ppscbe1=-1.462641884e-4
+  pscbe2=3.614130874e-09 lpscbe2=5.785994353e-15 wpscbe2=-1.353389859e-16 ppscbe2=7.085266590e-23
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=3.994354498e+01 lbeta0=-1.634218192e-05 wbeta0=-2.441314890e-05 pbeta0=1.278077171e-11
* Gidl Induced Drain Leakage Model Parameters
+  agidl=1.487772919e-10 lagidl=-7.788788786e-17 wagidl=-8.670636926e-17 pagidl=4.539251844e-23
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.216831793e-01 lkt1=-5.873117501e-8
+  kt2=-6.301890653e-02 lkt2=1.479981827e-8
+  at=3.649594374e+05 lat=-1.708698007e-01 wat=-2.039650751e-01 pat=1.067797961e-7
+  ute=-1.934483867e+00 lute=9.071704088e-7
+  ua1=-3.495144579e-09 lua1=3.136823287e-15 pua1=-1.654361225e-36
+  ub1=5.373218425e-18 lub1=-4.025826850e-24 wub1=-8.158603002e-25 pub1=4.271191844e-31
+  uc1=3.311138654e-10 luc1=-2.704089518e-16 wuc1=-2.067951531e-31 puc1=1.033975766e-37
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.75e-6
+  sbref=1.74e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.141 pmos
* Model Flag Parameters
+  lmin=2.5e-07 lmax=5.0e-07 wmin=7.0e-07 wmax=7.5e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.045892418e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-2.747137143e-9
+  k1=4.352213524e-01 lk1=3.901559036e-8
+  k2=1.408936088e-02 lk2=-1.064704755e-8
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=-1.888704683e-01 ldsub=2.662611400e-7
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-8.564575735e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=1.062985797e-7
+  nfactor={1.710086311e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.932506331e-7
+  eta0=4.117672797e-01 leta0=2.139821381e-8
+  etab=-1.291129272e-03 letab=3.335097045e-10
+  u0=7.485205816e-03 lu0=-5.094077095e-10
+  ua=-1.063421140e-09 lua=-7.182039643e-17
+  ub=1.148080500e-18 lub=4.611627323e-26
+  uc=-6.419271038e-11 luc=1.728726011e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=1.425608788e+05 lvsat=3.500072552e-3
+  a0=8.919849864e-01 la0=-7.572743094e-8
+  ags=9.698322768e-01 lags=1.466734064e-7
+  a1=0.0
+  a2=1.121568012e+00 la2=-8.904336116e-8
+  b0=1.836663184e-16 lb0=-5.023641140e-23
+  b1=7.635849659e-20 lb1=-2.088557599e-26
+  keta=-4.524308758e-02 lketa=3.703575468e-9
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-5.731343976e-01 lpclm=3.310509927e-07 wpclm=2.220446049e-22 ppclm=-1.665334537e-28
+  pdiblc1=-4.101030779e-01 lpdiblc1=2.228457367e-07 ppdiblc1=-8.326672685e-29
+  pdiblc2=-9.175377595e-03 lpdiblc2=4.855496791e-09 wpdiblc2=1.734723476e-24 ppdiblc2=3.144186300e-30
+  pdiblcb=2.408596814e-01 lpdiblcb=-1.446591300e-07 wpdiblcb=1.110223025e-22 ppdiblcb=2.775557562e-29
+  drout=1.436421824e+00 ldrout=-2.482852179e-7
+  pscbe1=6.925891618e+08 lpscbe1=2.937170827e+1
+  pscbe2=2.103542680e-08 lpscbe2=-3.334402489e-15
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=8.528056950e+00 lbeta0=1.044543745e-7
* Gidl Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=7.372237654e+08 lbgidl=1.375686143e+2
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.00074326333
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.5407449e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-5.460023937e-01 lkt1=6.352420121e-9
+  kt2=-1.498550792e-02 lkt2=-1.034662657e-8
+  at=6.500485322e+03 lat=1.679062992e-2
+  ute=4.908242408e-01 lute=-3.625268917e-07 pute=-2.220446049e-28
+  ua1=4.905387581e-09 lua1=-1.261023309e-15
+  ub1=-4.666106948e-18 lub1=1.229960769e-24
+  uc1=-2.811617509e-10 luc1=5.012957887e-17
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.1e-6
+  sbref=1.1e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.142 pmos
* Model Flag Parameters
+  lmin=1.8e-07 lmax=2.5e-07 wmin=7.0e-07 wmax=7.5e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.260936797e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=5.607180137e-08 wvth0=1.694120041e-07 pvth0=-4.633757136e-14
+  k1=-2.388367963e+00 lk1=8.113237399e-07 wk1=1.042648110e-06 pk1=-2.851851110e-13
+  k2=1.334853916e+00 lk2=-3.719025686e-07 wk2=-5.573203631e-07 pk2=1.524382657e-13
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=6.676943852e+00 ldsub=-1.611676393e-06 wdsub=-3.319827273e-06 pdsub=9.080391558e-13
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-5.970464504e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=1.505081755e-06 wvoff=3.569553490e-06 pvoff=-9.763442706e-13
+  nfactor={-8.338248924e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=2.346777190e-05 wnfactor=5.883863453e-05 pnfactor=-1.609354332e-11
+  eta0=1.110121481e+01 leta0=-2.902379475e-06 weta0=-7.229123536e-06 peta0=1.977309870e-12
+  etab=1.042326804e+00 letab=-2.851168675e-07 wetab=-7.086121574e-07 petab=1.938195973e-13
+  u0=1.434860387e-02 lu0=-2.386684346e-09 wu0=-6.631448256e-11 pu0=1.813833727e-17
+  ua=3.222999760e-10 lua=-4.508428360e-16 wua=9.529801071e-16 pua=-2.606591189e-22
+  ub=-5.317012365e-19 lub=5.055701737e-25 wub=-1.934431252e-25 pub=5.291056360e-32
+  uc=-4.914405300e-10 luc=1.341480837e-16 wuc=3.585779545e-16 puc=-9.807824210e-23
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=-7.107366610e+05 lvsat=2.368940156e-01 wvsat=7.306723963e-01 pvsat=-1.998535138e-7
+  a0=-1.019501200e+01 la0=2.956787986e-06 wa0=6.845670235e-06 pa0=-1.872427723e-12
+  ags=2.250598975e+00 lags=-2.036419008e-07 wags=7.580119643e-15 pags=-2.073313965e-21
+  a1=0.0
+  a2=4.992957653e+00 la2=-1.147945856e-06 wa2=-2.765509701e-06 pa2=7.564222134e-13
+  b0=0.0
+  b1=0.0
+  keta=-6.102501342e-01 lketa=1.582443028e-07 wketa=3.562234243e-07 pketa=-9.743423102e-14
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=6.337829886e-01 lpclm=9.349492092e-10 wpclm=3.487089744e-08 ppclm=-9.537887867e-15
+  pdiblc1=7.897290898e+00 lpdiblc1=-2.049392664e-06 wpdiblc1=-5.006379848e-06 ppdiblc1=1.369345016e-12
+  pdiblc2=-7.293104918e-02 lpdiblc2=2.229394808e-08 wpdiblc2=7.006630912e-08 ppdiblc2=-1.916453687e-14
+  pdiblcb=-2.760046981e+01 lpdiblcb=7.470501312e-06 wpdiblcb=2.029290987e-05 ppdiblcb=-5.550516707e-12
+  drout=-8.416496816e-01 ldrout=3.748129004e-07 wdrout=3.424960241e-12 pdrout=-9.367951250e-19
+  pscbe1=7.998956527e+08 lpscbe1=2.123688588e-02 wpscbe1=1.024650574e-06 ppscbe1=-2.802619934e-13
+  pscbe2=-6.764984646e-08 lpscbe2=2.092279345e-14 wpscbe2=5.942288006e-14 ppscbe2=-1.625334615e-20
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=1.062410412e+01 lbeta0=-4.688564472e-07 wbeta0=-6.651003022e-08 pbeta0=1.819182347e-14
* Gidl Induced Drain Leakage Model Parameters
+  agidl=-1.305110520e-13 lagidl=3.569738293e-20 wagidl=9.543907799e-20 pagidl=-2.610449661e-26
+  bgidl=1.938486420e+09 lbgidl=-1.910007469e+02 wbgidl=3.803092957e-06 pbgidl=-1.040224075e-12
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.00074326333
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.5407449e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-1.022859020e+01 lkt1=2.654733838e-06 wkt1=7.134586971e-06 pkt1=-1.951452228e-12
+  kt2=1.724989142e+00 lkt2=-4.862644929e-07 wkt2=-1.215182230e-06 pkt2=3.323766436e-13
+  at=-6.892421477e+05 lat=2.070901549e-01 wat=6.140717803e-01 pat=-1.679609133e-7
+  ute=-1.885049126e+01 lute=4.927709725e-06 wute=1.157781658e-05 pute=-3.166764391e-12
+  ua1=-1.530382061e-08 lua1=4.266599314e-15 wua1=1.051823409e-14 pua1=-2.876947388e-21
+  ub1=1.374079099e-17 lub1=-3.804693956e-24 wub1=-9.586405349e-24 pub1=2.622073591e-30
+  uc1=-5.860694786e-10 luc1=1.335279405e-16 wuc1=1.967359732e-16 puc1=-5.381122340e-23
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.1e-6
+  sbref=1.1e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.143 pmos
* Model Flag Parameters
+  lmin=1.5e-07 lmax=1.8e-07 wmin=7.0e-07 wmax=7.5e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-2.026e-8
+  vth0={-4.170736186e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-1.253332362e-07 wvth0=-4.562507215e-07 pvth0=8.776300138e-14
+  k1=3.923540565e+00 lk1=-5.128085587e-07 wk1=-2.003929217e-06 pk1=3.628246447e-13
+  k2=-1.984709832e+00 lk2=3.290626543e-07 wk2=1.286641485e-06 pk2=-2.414590520e-13
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=-8.646388305e+00 ldsub=1.632801688e-06 wdsub=6.380583114e-06 pdsub=-1.155246946e-12
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={1.119462482e+01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-2.154444452e-06 wvoff=-8.309681160e-06 pvoff=1.561710640e-12
+  nfactor={2.053570187e+02+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-3.824480436e-05 wnfactor=-1.441507578e-04 pnfactor=2.732538583e-11
+  eta0=-1.928303368e+01 leta0=3.555519609e-06 weta0=1.389409174e-05 peta0=-2.515617117e-12
+  etab=-1.939042449e+00 letab=3.485189043e-07 wetab=1.361925416e-06 petab=-2.465856219e-13
+  u0=8.135153008e-04 lu0=3.987139427e-10 wu0=1.701031560e-09 pu0=-3.700817190e-16
+  ua=2.325375246e-10 lua=-4.687072656e-16 wua=-1.831591807e-15 pua=3.316218562e-22
+  ub=1.520982037e-18 lub=9.514267123e-26 wub=3.717929856e-25 pub=-6.731569083e-32
+  uc=9.674468586e-10 luc=-1.763603906e-16 wuc=-6.891727905e-16 puc=1.247792890e-22
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=2.715878168e+06 lvsat=-4.989553591e-01 wvsat=-1.899352624e+00 pvsat=3.634258647e-7
+  a0=1.960134241e+01 la0=-3.366923961e-06 wa0=-1.315710657e-05 pa0=2.382180966e-12
+  ags=1.250000091e+00 lags=-1.734492727e-14 wags=-1.916431813e-14 pags=3.651187797e-21
+  a1=0.0
+  a2=-6.815504052e+00 la2=1.360168346e-06 wa2=5.315201549e-06 pa2=-9.623523792e-13
+  b0=0.0
+  b1=0.0
+  keta=9.617837140e-01 lketa=-1.752024746e-07 wketa=-6.846478017e-07 pketa=1.239600227e-13
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=7.161501427e-01 lpclm=-1.715055943e-08 wpclm=-6.702023098e-08 ppclm=1.213444520e-14
+  pdiblc1=-1.333833501e+01 lpdiblc1=2.462302050e-06 wpdiblc1=9.622067394e-06 ppdiblc1=-1.742138953e-12
+  pdiblc2=1.928818345e-01 lpdiblc2=-3.446089834e-08 wpdiblc2=-1.346646833e-07 ppdiblc2=2.438193022e-14
+  pdiblcb=5.436592266e+01 lpdiblcb=-9.980717520e-06 wpdiblcb=-3.900217678e-05 ppdiblcb=7.061601838e-12
+  drout=1.000012903e+00 ldrout=-2.458418830e-12 wdrout=-8.659109056e-12 pdrout=1.649733457e-18
+  pscbe1=8.000000043e+08 lpscbe1=-8.308391571e-07 wpscbe1=-2.590553284e-06 ppscbe1=4.935512543e-13
+  pscbe2=1.676875032e-07 lpscbe2=-2.922612059e-14 wpscbe2=-1.142084541e-13 ppscbe2=2.067819569e-20
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=8.172020727e+00 lbeta0=3.271346236e-08 wbeta0=1.278337559e-07 pbeta0=-2.314530753e-14
* Gidl Induced Drain Leakage Model Parameters
+  agidl=3.299627887e-13 lagidl=-6.286451050e-20 wagidl=-2.412925484e-19 pagidl=4.597105632e-26
+  bgidl=1.000000333e+09 lbgidl=-6.340809631e-05 wbgidl=-9.615112305e-06 pbgidl=1.831874847e-12
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-1.106e-8
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=2.310683730e+01 lkt1=-4.474645051e-06 wkt1=-1.722103721e-05 pkt1=3.256445458e-12
+  kt2=-3.374541169e+00 lkt2=5.976663193e-07 wkt2=2.335532195e-06 pkt2=-4.228635221e-13
+  at=1.697883648e+06 lat=-3.020206109e-01 wat=-1.180221861e+00 pat=2.136869664e-7
+  ute=3.118429147e+01 lute=-5.694349590e-06 wute=-2.225211034e-05 pute=4.028891662e-12
+  ua1=2.911935419e-08 lua1=-5.173210687e-15 wua1=-2.021562911e-14 pua1=3.660173070e-21
+  ub1=-2.633452210e-17 lub1=4.714908480e-24 wub1=1.842469586e-23 pub1=-3.335912970e-30
+  uc1=5.088094453e-10 luc1=-9.676118767e-17 wuc1=-3.781188054e-16 puc1=6.846090766e-23
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.04e-6
+  sbref=1.04e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.144 pmos
* Model Flag Parameters
+  lmin=2.0e-05 lmax=0.0001 wmin=6.4e-07 wmax=7.0e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.126311+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+  k1=0.43165561
+  k2=0.026980026
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=3.2465718e-7
+  voff={-0.23051772+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.8768912+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+  eta0=0.08
+  etab=-0.07
+  u0=0.0095864
+  ua=-7.4757916e-10
+  ub=9.5046395e-19
+  uc=-1.0566299e-10
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=80156.0
+  a0=1.464
+  ags=0.11329
+  a1=0.0
+  a2=0.97
+  b0=-8.9873e-8
+  b1=3.3859e-9
+  keta=0.023361259
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=0.015
+  pdiblc1=0.39
+  pdiblc2=0.0012771588
+  pdiblcb=-0.225
+  drout=0.56
+  pscbe1=800000000.0
+  pscbe2=1.0060625e-8
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=0.0
+  alpha1=0.0
+  beta0=30.0
* Gidl Induced Drain Leakage Model Parameters
+  agidl=9.43573999999999e-11
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-0.43825
+  kt2=-0.058546
+  at=70990.0
+  ute=-0.08298
+  ua1=2.0902e-9
+  ub1=-1.2289e-18
+  uc1=-2.9789e-11
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.145 pmos
* Model Flag Parameters
+  lmin=8.0e-06 lmax=2.0e-05 wmin=6.4e-07 wmax=7.0e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.163749012e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=7.496407775e-7
+  k1=4.170420989e-01 lk1=2.926139320e-7
+  k2=2.824548822e-02 lk2=-2.533900806e-8
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=-6.144535039e-06 lcit=1.295359998e-10 wcit=-3.388131789e-27 pcit=5.421010862e-32
+  voff={-2.486350287e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=3.627722941e-7
+  nfactor={2.137127920e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-5.210855164e-6
+  eta0=0.08
+  etab=-0.07
+  u0=1.063746106e-02 lu0=-2.104594218e-8
+  ua=-9.116420042e-10 lua=3.285115641e-15
+  ub=1.339640455e-18 lub=-7.792683529e-24
+  uc=-1.046534774e-10 luc=-2.021399574e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=9.292141765e+04 lvsat=-2.556085955e-1
+  a0=1.626529302e+00 la0=-3.254408731e-6
+  ags=1.127437120e-01 lags=1.093860960e-8
+  a1=0.0
+  a2=1.083666533e+00 la2=-2.276004104e-6
+  b0=-1.709446520e-07 lb0=1.623339844e-12
+  b1=5.452591595e-09 lb1=-4.138244049e-14
+  keta=3.421368674e-02 lketa=-2.173038039e-7
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-6.921953293e-02 lpclm=1.686371502e-06 wpclm=-2.775557562e-23 ppclm=4.440892099e-28
+  pdiblc1=0.39
+  pdiblc2=1.909636661e-03 lpdiblc2=-1.266443309e-8
+  pdiblcb=-0.225
+  drout=0.56
+  pscbe1=800000000.0
+  pscbe2=8.860770435e-09 lpscbe2=2.402531188e-14
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=-6.686266667e-11 lalpha0=1.338825943e-15
+  alpha1=-6.686266667e-11 lalpha1=1.338825943e-15
+  beta0=4.805292000e+01 lbeta0=-3.614830047e-04 pbeta0=4.547473509e-25
* Gidl Induced Drain Leakage Model Parameters
+  agidl=1.354378090e-10 lagidl=-8.225743918e-16
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.443915098e-01 lkt1=1.229746438e-7
+  kt2=-6.522345350e-02 lkt2=1.337061237e-7
+  at=7.716025872e+04 lat=-1.235502988e-1
+  ute=5.623649524e-01 lute=-1.292207756e-05 pute=-4.440892099e-27
+  ua1=3.775543044e-09 lua1=-3.374650014e-14
+  ub1=-2.648919653e-18 lub1=2.843379192e-23
+  uc1=-9.445040192e-11 luc1=1.294748875e-15 wuc1=5.169878828e-32
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.146 pmos
* Model Flag Parameters
+  lmin=4.0e-06 lmax=8.0e-06 wmin=6.4e-07 wmax=7.0e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.036424065e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-2.719534781e-7
+  k1=4.604103273e-01 lk1=-5.535191579e-8
+  k2=3.111376993e-02 lk2=-4.835272375e-8
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-1.903188674e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-1.051285932e-7
+  nfactor={7.782034620e-01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=5.692502402e-6
+  eta0=0.08
+  etab=-0.07
+  u0=5.374816804e-03 lu0=2.117898927e-8
+  ua=-5.231013447e-10 lua=1.676518894e-16
+  ub=-7.890771535e-20 lub=3.589066086e-24
+  uc=-1.070071013e-10 luc=-1.329647545e-18
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=6.344101412e+04 lvsat=-1.907198821e-2
+  a0=1.169202877e+00 la0=4.149589883e-7
+  ags=4.476786908e-02 lags=5.563441444e-7
+  a1=0.0
+  a2=0.8
+  b0=1.333762438e-07 lb0=-8.183849488e-13 wb0=5.293955920e-29 pb0=-2.117582368e-34
+  b1=-1.241682582e-09 lb1=1.232920225e-14 pb1=6.617444900e-36
+  keta=7.540400483e-03 lketa=-3.290158170e-9
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-4.109336388e-01 lpclm=4.428121465e-06 ppclm=-1.776356839e-27
+  pdiblc1=0.39
+  pdiblc2=2.318653116e-04 lpdiblc2=7.971988815e-10
+  pdiblcb=-0.225
+  drout=0.56
+  pscbe1=800000000.0
+  pscbe2=1.463489899e-08 lpscbe2=-2.230352405e-14
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=2.005880000e-10 lalpha0=-8.070698298e-16
+  alpha1=2.005880000e-10 lalpha1=-8.070698298e-16
+  beta0=-2.415876000e+01 lbeta0=2.179088540e-04 wbeta0=1.421085472e-20 pbeta0=5.684341886e-26
* Gidl Induced Drain Leakage Model Parameters
+  agidl=4.884466474e-11 lagidl=-1.277925667e-16
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.137901907e-01 lkt1=-1.225556520e-7
+  kt2=-3.851363950e-02 lkt2=-8.060060310e-8
+  at=2.230282385e+04 lat=3.165994270e-1
+  ute=-1.918426857e+00 lute=6.982605139e-06 wute=-1.776356839e-21
+  ua1=-2.965829131e-09 lua1=2.034303433e-14
+  ub1=2.930570959e-18 lub1=-1.633336259e-23 wub1=1.540743956e-39 pub1=1.232595164e-44
+  uc1=5.548297096e-10 luc1=-3.914763086e-15 wuc1=2.067951531e-31 puc1=8.271806126e-37
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.147 pmos
* Model Flag Parameters
+  lmin=2.0e-06 lmax=4.0e-06 wmin=6.4e-07 wmax=7.0e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.106065230e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=8.249143277e-9
+  k1=3.853412315e-01 lk1=2.466900923e-7
+  k2=4.064949326e-02 lk2=-8.671989728e-8
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=8.635279899e-01 ldsub=-1.221250938e-6
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.223718520e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=2.383723148e-8
+  nfactor={2.270962668e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-3.136441188e-7
+  eta0=1.604349200e-01 leta0=-3.236315093e-7
+  etab=-1.403173200e-01 letab=2.829231434e-7
+  u0=1.211265930e-02 lu0=-5.930854756e-9
+  ua=-1.308633256e-10 lua=-1.410525625e-15
+  ub=6.187485939e-19 lub=7.820319721e-25
+  uc=-1.338088641e-10 luc=1.065077811e-16
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=8.388955365e+04 lvsat=-1.013470960e-1
+  a0=1.400765170e+00 la0=-5.167365282e-7
+  ags=-4.432097709e-02 lags=9.147948988e-7
+  a1=0.0
+  a2=0.8
+  b0=-1.003353178e-07 lb0=1.219581936e-13
+  b1=1.451284080e-09 lb1=1.493997030e-15
+  keta=2.281093733e-02 lketa=-6.473146857e-8
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=6.059902523e-01 lpclm=3.365078504e-7
+  pdiblc1=0.39
+  pdiblc2=4.185431636e-04 lpdiblc2=4.609681023e-11
+  pdiblcb=-4.273520000e-01 lpdiblcb=8.141673190e-7
+  drout=0.56
+  pscbe1=800000000.0
+  pscbe2=8.712478508e-09 lpscbe2=1.525453199e-15
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=-1.011760000e-10 lalpha0=4.070836595e-16
+  alpha1=-1.011760000e-10 lalpha1=4.070836595e-16
+  beta0=5.471942625e+01 lbeta0=-9.945910591e-5
* Gidl Induced Drain Leakage Model Parameters
+  agidl=1.634728531e-11 lagidl=2.961289373e-18
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.355286288e-01 lkt1=-3.509061145e-8
+  kt2=-6.321122536e-02 lkt2=1.877062754e-8
+  at=1.626547485e+05 lat=-2.481093488e-1
+  ute=-9.154724880e-02 lute=-3.678815031e-7
+  ua1=2.886961000e-09 lua1=-3.205783819e-15 wua1=3.308722450e-30
+  ub1=-1.904818744e-18 lub1=3.121924585e-24
+  uc1=-8.771411122e-10 luc1=1.846800155e-15
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.148 pmos
* Model Flag Parameters
+  lmin=1.0e-06 lmax=2.0e-06 wmin=6.4e-07 wmax=7.0e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.118108631e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=3.261920430e-8
+  k1=5.064652470e-01 lk1=1.593224533e-9
+  k2=-2.759691298e-03 lk2=1.119455858e-9
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=2.600000202e-01 ldsub=-2.071113148e-14
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.052413704e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-1.082664065e-8
+  nfactor={2.508128773e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-7.935544749e-7
+  eta0=-5.005130400e-01 leta0=1.013809907e-06 weta0=1.977584763e-22 peta0=2.576064362e-28
+  etab=2.645421120e-04 letab=-1.547066255e-09 petab=-8.673617380e-31
+  u0=1.145910416e-02 lu0=-4.608372862e-9
+  ua=-3.318390994e-10 lua=-1.003847127e-15
+  ub=7.130469709e-19 lub=5.912173203e-25
+  uc=-1.196469642e-10 luc=7.785089353e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=1.537394825e+04 lvsat=3.729560184e-2
+  a0=1.030938530e+00 la0=2.316150734e-7
+  ags=2.475687006e-01 lags=3.241502982e-7
+  a1=0.0
+  a2=0.8
+  b0=2.062768896e-08 lb0=-1.228128700e-13
+  b1=-2.754611245e-08 lb1=6.017080885e-14 wb1=-6.617444900e-30 pb1=-1.323488980e-35
+  keta=-1.751182380e-02 lketa=1.686244502e-8
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=9.199174115e-01 lpclm=-2.987300348e-7
+  pdiblc1=3.957940034e-01 lpdiblc1=-1.172428182e-8
+  pdiblc2=4.529136727e-04 lpdiblc2=-2.345260230e-11
+  pdiblcb=1.797040000e-01 lpdiblcb=-4.142226381e-07 wpdiblcb=1.110223025e-22
+  drout=3.794864141e-01 ldrout=3.652728512e-7
+  pscbe1=800000000.0
+  pscbe2=9.769526283e-09 lpscbe2=-6.135041137e-16
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=4.643241089e+00 lbeta0=1.871056290e-6
* Gidl Induced Drain Leakage Model Parameters
+  agidl=2.528734937e-11 lagidl=-1.512910906e-17
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.260591597e-01 lkt1=-5.425227153e-8
+  kt2=-5.943725826e-02 lkt2=1.113392964e-8
+  at=2.804660864e+04 lat=2.427291432e-2
+  ute=5.196833265e-01 lute=-1.604718797e-06 pute=4.440892099e-28
+  ua1=3.076566596e-09 lua1=-3.589454534e-15
+  ub1=-1.607506698e-18 lub1=2.520307714e-24 pub1=1.540743956e-45
+  uc1=3.394859767e-12 luc1=6.501800488e-17
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=2.75e-6
+  sbref=2.74e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.149 pmos
* Model Flag Parameters
+  lmin=5.0e-07 lmax=1.0e-06 wmin=6.4e-07 wmax=7.0e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.318215689e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=2.374327807e-07 wvth0=1.330023330e-07 pvth0=-1.361305479e-13
+  k1=-3.047362452e-01 lk1=8.318741759e-07 wk1=5.524788691e-07 pk1=-5.654731721e-13
+  k2=4.002227781e-01 lk2=-4.113411612e-07 wk2=-2.705270439e-07 pk2=2.768898400e-13
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=7.572714005e+00 ldsub=-7.484709039e-06 wdsub=-5.024551965e-06 pdsub=5.142729427e-12
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={5.119371148e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-5.460674046e-06 wvoff=-3.322572773e-06 pvoff=3.400719684e-12
+  nfactor={1.001902646e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-8.481108477e-06 wnfactor=-5.892270791e-06 pnfactor=6.030857000e-12
+  eta0=-4.289659422e+00 leta0=4.892077011e-06 weta0=3.282897014e-06 peta0=-3.360110752e-12
+  etab=-5.618112549e-03 letab=4.473948444e-09 wetab=2.555010427e-09 petab=-2.615104272e-15
+  u0=2.988221817e-02 lu0=-2.346479851e-08 wu0=-1.530151477e-08 pu0=1.566140640e-14
+  ua=2.974418634e-09 lua=-4.387868043e-15 wua=-3.000536854e-15 pua=3.071109481e-21
+  ub=-1.750169136e-18 lub=3.112368270e-24 wub=2.110526628e-24 pub=-2.160166214e-30
+  uc=-2.426354036e-10 luc=2.037320210e-16 wuc=1.267526206e-16 puc=-1.297338422e-22
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=-6.247725462e+05 lvsat=6.924983419e-01 wvsat=3.914369197e-01 pvsat=-4.006435160e-7
+  a0=5.769610677e+00 la0=-4.618510642e-06 wa0=-2.710438758e-06 pa0=2.774188277e-12
+  ags=-1.537163700e-01 lags=7.348735937e-07 wags=-4.362963324e-16 pags=4.465601222e-22
+  a1=0.0
+  a2=-4.338442546e+00 la2=5.259298714e-06 wa2=3.392621944e-06 pa2=-3.472416412e-12
+  b0=-2.034000366e-07 lb0=1.064839877e-13 wb0=6.478143980e-22 pb0=-6.630510384e-28
+  b1=6.395362368e-08 lb1=-3.348100107e-14 wb1=2.693035377e-25 pb1=-2.756562848e-31
+  keta=-2.029414668e-02 lketa=1.971020813e-08 wketa=3.960629574e-08 pketa=-4.053783582e-14
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=5.270649158e+00 lpclm=-4.751790991e-06 wpclm=-2.757113803e-06 ppclm=2.821961120e-12
+  pdiblc1=1.359239429e+00 lpdiblc1=-9.978299443e-07 wpdiblc1=-4.011186353e-07 ppdiblc1=4.105529456e-13
+  pdiblc2=8.411932156e-03 lpdiblc2=-8.169667200e-09 wpdiblc2=-5.201996227e-09 ppdiblc2=5.324347178e-15
+  pdiblcb=-2.478369146e+00 lpdiblcb=2.306368389e-06 wpdiblcb=1.399955156e-06 ppdiblcb=-1.432882102e-12
+  drout=-4.380787899e+00 ldrout=5.237508817e-06 wdrout=3.325109321e-06 pdrout=-3.403315892e-12
+  pscbe1=-5.764093430e+09 lpscbe1=6.718480908e+03 wpscbe1=4.508531010e+03 ppscbe1=-4.614571659e-3
+  pscbe2=6.919512782e-07 lpscbe2=-6.988401709e-13 wpscbe2=-4.690801641e-13 ppscbe2=4.801129295e-19
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=1.014046269e+00 lbeta0=5.585609772e-06 wbeta0=2.108428552e-06 pbeta0=-2.158018792e-12
* Gidl Induced Drain Leakage Model Parameters
+  agidl=2.178139562e-10 lagidl=-2.121839417e-16 wagidl=-1.337391156e-16 pagidl=1.368846596e-22
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=1.202709299e-01 lkt1=-6.134320449e-07 wkt1=-3.692181599e-07 pkt1=3.779021710e-13
+  kt2=-3.318357464e-01 lkt2=2.899392302e-07 wkt2=1.831373861e-07 pkt2=-1.874447775e-13
+  at=5.147056721e+05 lat=-4.738323703e-01 wat=-3.059829918e-01 pat=3.131797118e-7
+  ute=-2.335023866e+00 lute=1.317131108e-06 wute=2.728766862e-07 pute=-2.792947458e-13
+  ua1=-1.250504413e-08 lua1=1.235863567e-14 wua1=6.138192284e-15 pua1=-6.282562567e-21
+  ub1=1.989883382e-17 lub1=-1.949186193e-23 wub1=-1.071175535e-23 pub1=1.096369584e-29
+  uc1=1.611051657e-09 luc1=-1.580450880e-15 wuc1=-8.719857791e-16 puc1=8.924948846e-22
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.75e-6
+  sbref=1.74e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.150 pmos
* Model Flag Parameters
+  lmin=2.5e-07 lmax=5.0e-07 wmin=6.4e-07 wmax=7.0e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-6.554394620e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-1.095438296e-07 wvth0=-2.660046661e-07 pvth0=7.275759627e-14
+  k1=2.057125288e+00 lk1=-4.046075742e-07 wk1=-1.104957738e-06 pk1=3.022280406e-13
+  k2=-7.800928274e-01 lk2=2.065776646e-07 wk2=5.410540878e-07 pk2=-1.479891141e-13
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=-1.493937237e+01 ldsub=4.300818420e-06 wdsub=1.004910393e-05 pdsub=-2.748630907e-12
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-1.061048467e+01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=2.774220070e-06 wvoff=6.645145545e-06 pvoff=-1.817580210e-12
+  nfactor={-1.558776474e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=4.924558853e-06 wnfactor=1.178454158e-05 pnfactor=-3.223307813e-12
+  eta0=1.004931884e+01 leta0=-2.614664890e-06 weta0=-6.565794029e-06 peta0=1.795875983e-12
+  etab=6.209576546e-03 letab=-1.718083351e-09 wetab=-5.110020854e-09 petab=1.397692904e-15
+  u0=-3.743522178e-02 lu0=1.177722765e-08 wu0=3.060302955e-08 pu0=-8.370540641e-15
+  ua=-9.872052212e-09 lua=2.337516375e-15 wua=6.001073708e-15 pua=-1.641413681e-21
+  ub=7.343921890e-18 lub=-1.648570264e-24 wub=-4.221053256e-24 pub=1.154542486e-30
+  uc=3.079130582e-10 luc=-8.449110970e-17 wuc=-2.535052412e-16 puc=6.933875356e-23
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=1.291696377e+06 lvsat=-3.108114690e-01 wvsat=-7.828738394e-01 pvsat=2.141316526e-7
+  a0=-7.065009452e+00 la0=2.100669688e-06 wa0=5.420877515e-06 pa0=-1.482718418e-12
+  ags=9.698322756e-01 lags=1.466734067e-07 wags=8.725926648e-16 pags=-2.386721931e-22
+  a1=0.0
+  a2=1.108123741e+01 la2=-2.813212134e-06 wa2=-6.785243888e-06 pa2=1.855899908e-12
+  b0=2.085445334e-15 lb0=-5.704110078e-22 wb0=-1.295628794e-21 pb0=3.543803876e-28
+  b1=8.670150949e-19 lb1=-2.371459687e-25 wb1=-5.386522020e-25 pb1=1.473321503e-31
+  keta=7.102852124e-02 lketa=-2.809903498e-08 wketa=-7.921259149e-08 pketa=2.166622802e-14
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-8.667152067e+00 lpclm=2.544926706e-06 wpclm=5.514227606e-06 ppclm=-1.508251535e-12
+  pdiblc1=-1.587661044e+00 lpdiblc1=5.449313916e-07 wpdiblc1=8.022372707e-07 ppdiblc1=-2.194279383e-13
+  pdiblc2=-2.444679995e-02 lpdiblc2=9.032536234e-09 wpdiblc2=1.040399245e-08 ppdiblc2=-2.845700016e-15
+  pdiblcb=4.350687052e+00 lpdiblcb=-1.268779112e-06 wpdiblcb=-2.799910313e-06 ppdiblcb=7.658314687e-13
+  drout=1.119789542e+01 ldrout=-2.918243477e-06 wdrout=-6.650218642e-06 pdrout=1.818967803e-12
+  pscbe1=1.392821608e+10 lpscbe1=-3.590836966e+03 wpscbe1=-9.017062020e+03 ppscbe1=2.466346804e-3
+  pscbe2=-1.356036181e-06 lpscbe2=3.733222236e-13 wpscbe2=9.381603281e-13 ppscbe2=-2.566056129e-19
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=1.471773905e+01 lbeta0=-1.588547474e-06 wbeta0=-4.216857105e-06 pbeta0=1.153394755e-12
* Gidl Induced Drain Leakage Model Parameters
+  agidl=-3.926159173e-10 lagidl=1.073883057e-16 wagidl=2.674782312e-16 pagidl=-7.316064580e-23
+  bgidl=7.372237654e+08 lbgidl=1.375686143e+2
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.00074326333
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.5407449e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-1.629910612e+00 lkt1=3.028229960e-07 wkt1=7.384363198e-07 pkt1=-2.019771022e-13
+  kt2=5.226481719e-01 lkt2=-1.574001907e-07 wkt2=-3.662747723e-07 pkt2=1.001834757e-13
+  at=-8.917691980e+05 lat=2.624853537e-01 wat=6.119659837e-01 pat=-1.673849359e-7
+  ute=1.291904239e+00 lute=-5.816382927e-07 wute=-5.457533723e-07 pute=1.492744624e-13
+  ua1=2.292518668e-08 lua1=-6.189798757e-15 wua1=-1.227638457e-14 pua1=3.357836707e-21
+  ub1=-3.611244660e-17 lub1=9.831163589e-24 wub1=2.142351070e-23 pub1=-5.859758648e-30
+  uc1=-2.841037334e-09 luc1=7.503067483e-16 wuc1=1.743971558e-15 puc1=-4.770111006e-22
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.1e-6
+  sbref=1.1e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.151 pmos
* Model Flag Parameters
+  lmin=1.8e-07 lmax=2.5e-07 wmin=6.4e-07 wmax=7.0e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.012266656e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-1.194445551e-8
+  k1=-8.579247482e-01 lk1=3.927169118e-7
+  k2=5.167953973e-01 lk2=-1.481472026e-07 wk2=1.110223025e-22 pk2=5.551115123e-29
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=1.803960266e+00 ldsub=-2.788179225e-7
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-7.309221625e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=7.196213411e-8
+  nfactor={2.983359543e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.550150614e-7
+  eta0=4.900000008e-01 leta0=-7.095923849e-17
+  etab=2.195759126e-03 letab=-6.202240101e-10 wetab=-8.673617380e-25 petab=1.084202172e-31
+  u0=1.425126466e-02 lu0=-2.360060124e-9
+  ua=1.721124685e-09 lua=-8.334493704e-16
+  ub=-8.156452782e-19 lub=5.832345480e-25
+  uc=3.489543344e-11 luc=-9.815328983e-18 wuc=1.292469707e-32 puc=5.654554969e-39
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=3.617753405e+05 lvsat=-5.645946701e-2
+  a0=-1.466462483e-01 la0=2.083589844e-7
+  ags=2.250598986e+00 lags=-2.036419039e-7
+  a1=0.0
+  a2=9.336249622e-01 la2=-3.763717830e-8
+  b0=0.0
+  b1=0.0
+  keta=-8.737025015e-02 lketa=1.522619697e-08 wketa=1.110223025e-22
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=6.849679741e-01 lpclm=-1.306516802e-8
+  pdiblc1=5.487137542e-01 lpdiblc1=-3.940984321e-8
+  pdiblc2=2.991525761e-02 lpdiblc2=-5.836573751e-9
+  pdiblcb=2.186325871e+00 lpdiblcb=-6.767830420e-7
+  drout=-8.416446543e-01 ldrout=3.748115253e-7
+  pscbe1=7.998956542e+08 lpscbe1=2.123647450e-2
+  pscbe2=1.957358274e-08 lpscbe2=-2.934558902e-15
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=1.052647787e+01 lbeta0=-4.421537155e-7
* Gidl Induced Drain Leakage Model Parameters
+  agidl=9.578483481e-15 lagidl=-2.619906802e-21
+  bgidl=1.938486425e+09 lbgidl=-1.910007484e+2
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.00074326333
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.5407449e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=2.438598179e-01 lkt1=-2.096906920e-7
+  kt2=-5.870698811e-02 lkt2=1.612072696e-9
+  at=2.121185134e+05 lat=-3.945001311e-2
+  ute=-1.856079955e+00 lute=2.793983441e-7
+  ua1=1.352904843e-10 lua1=4.369364895e-17
+  ub1=-3.305422621e-19 lub1=4.409711620e-26
+  uc1=-2.972920545e-10 luc1=5.454153952e-17
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.1e-6
+  sbref=1.1e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.152 pmos
* Model Flag Parameters
+  lmin=1.5e-07 lmax=1.8e-07 wmin=6.4e-07 wmax=7.0e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-2.026e-8
+  vth0={-1.253367155e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=4.022530760e-08 wvth0=1.134926485e-07 pvth0=-2.502739885e-14
+  k1=5.421836102e-02 lk1=2.243747076e-07 wk1=6.321316589e-07 pk1=-1.393976734e-13
+  k2=1.094714173e+00 lk2=-2.879645683e-07 wk2=-8.112838655e-07 pk2=1.789043180e-13
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=3.673666038e+00 ldsub=-7.144150654e-07 wdsub=-2.012724948e-06 pdsub=4.438461056e-13
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-7.477819189e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=1.565798854e-06 wvoff=4.411332113e-06 pvoff=-9.727869576e-13
+  nfactor={-9.378406977e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=2.117119006e-05 wnfactor=5.964568986e-05 pnfactor=-1.315306753e-11
+  eta0=7.544625565e+00 leta0=-1.555686030e-06 weta0=-4.382841332e-06 peta0=9.665041706e-13
+  etab=6.906546923e-01 letab=-1.524909952e-07 wetab=-4.296136149e-07 petab=9.473839435e-14
+  u0=1.010419726e-02 lu0=-1.642684346e-09 wu0=-4.628449918e-09 pu0=1.020665776e-15
+  ua=-3.304021960e-09 lua=2.050780466e-16 wua=5.777671459e-16 pua=-1.274092110e-22
+  ub=2.238859668e-18 lub=-4.162737417e-26 wub=-1.172769433e-25 pub=2.586191154e-32
+  uc=-3.632548687e-10 luc=7.716490245e-17 wuc=2.173970366e-16 puc=-4.794039452e-23
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=-1.691861975e+06 lvsat=3.916925817e-01 wvsat=1.103517319e+00 pvsat=-2.433476393e-7
+  a0=-5.803301371e+00 la0=1.473168772e-06 wa0=4.150365909e-06 pa0=-9.152386902e-13
+  ags=1.250000062e+00 lags=-1.182880638e-14 wags=4.842775070e-16 pags=-1.067927968e-22
+  a1=0.0
+  a2=3.447448506e+00 la2=-5.951293749e-07 wa2=-1.676660665e-06 pa2=3.697372099e-13
+  b0=0.0
+  b1=0.0
+  keta=-3.601802273e-01 lketa=7.665809545e-08 wketa=2.159692165e-07 pketa=-4.762553162e-14
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=5.867423976e-01 lpclm=7.504204276e-09 wpclm=2.114164239e-08 ppclm=-4.662154979e-15
+  pdiblc1=5.240605014e+00 lpdiblc1=-1.077357603e-06 wpdiblc1=-3.035244235e-06 ppdiblc1=6.693320587e-13
+  pdiblc2=-6.713793942e-02 lpdiblc2=1.507806899e-08 wpdiblc2=4.247950810e-08 ppdiblc2=-9.367581126e-15
+  pdiblcb=-2.094213764e+01 lpdiblcb=4.366974129e-06 wpdiblcb=1.230309608e-05 ppdiblcb=-2.713078747e-12
+  drout=1.000000221e+00 ldrout=-4.311984192e-14 wdrout=-1.930837357e-14 pdrout=4.257882935e-21
+  pscbe1=8.000000018e+08 lpscbe1=-3.814220428e-07 wpscbe1=-8.497085571e-07 ppscbe1=1.873769760e-13
+  pscbe2=-5.283394308e-08 lpscbe2=1.278762535e-14 wpscbe2=3.602663267e-14 ppscbe2=-7.944593037e-21
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=8.418842974e+00 lbeta0=-1.431111250e-08 wbeta0=-4.031932991e-08 pbeta0=8.891218632e-15
* Gidl Induced Drain Leakage Model Parameters
+  agidl=-2.421667034e-14 lagidl=4.613760032e-21
+  bgidl=1.000000301e+09 lbgidl=-5.672953796e-05 wbgidl=1.232560730e-05 pbgidl=-2.718044281e-12
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-1.106e-8
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-1.650650532e+01 lkt1=3.466584391e-06 wkt1=9.766423937e-06 pkt1=-2.153691807e-12
+  kt2=1.135064268e+00 lkt2=-2.615037085e-07 wkt2=-7.367357205e-07 pkt2=1.624649611e-13
+  at=-5.809691612e+05 lat=1.321464263e-01 wat=3.722967503e-01 pat=-8.209887937e-8
+  ute=-1.178159732e+01 lute=2.491511542e-06 wute=7.019346647e-06 pute=-1.547906323e-12
+  ua1=-9.914368045e-09 lua1=2.263494073e-15 wua1=6.376952908e-15 pua1=-1.406245655e-21
+  ub1=9.241134442e-18 lub1=-2.062965604e-24 wub1=-5.812002826e-24 pub1=1.281662863e-30
+  uc1=-2.212881416e-10 luc1=4.233700458e-17 wuc1=1.192762379e-16 puc1=-2.630279597e-23
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.04e-6
+  sbref=1.04e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.153 pmos
* Model Flag Parameters
+  lmin=2.0e-05 lmax=0.0001 wmin=6.3e-07 wmax=6.4e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.126311+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+  k1=0.43165561
+  k2=0.026980026
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=3.2465718e-7
+  voff={-0.23051772+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.8768912+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+  eta0=0.08
+  etab=-0.07
+  u0=0.0095864
+  ua=-7.4757916e-10
+  ub=9.5046395e-19
+  uc=-1.0566299e-10
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=80156.0
+  a0=1.464
+  ags=0.11329
+  a1=0.0
+  a2=0.97
+  b0=-8.9873e-8
+  b1=3.3859e-9
+  keta=0.023361259
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=0.015
+  pdiblc1=0.39
+  pdiblc2=0.0012771588
+  pdiblcb=-0.225
+  drout=0.56
+  pscbe1=800000000.0
+  pscbe2=1.0060625e-8
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=0.0
+  alpha1=0.0
+  beta0=30.0
* Gidl Induced Drain Leakage Model Parameters
+  agidl=9.43573999999999e-11
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-0.43825
+  kt2=-0.058546
+  at=70990.0
+  ute=-0.08298
+  ua1=2.0902e-9
+  ub1=-1.2289e-18
+  uc1=-2.9789e-11
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.154 pmos
* Model Flag Parameters
+  lmin=8.0e-06 lmax=2.0e-05 wmin=6.3e-07 wmax=6.4e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.163749012e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=7.496407775e-7
+  k1=4.170420989e-01 lk1=2.926139320e-7
+  k2=2.824548822e-02 lk2=-2.533900806e-08 wk2=-2.220446049e-22
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=-6.144535039e-06 lcit=1.295359998e-10 wcit=-1.016439537e-26 pcit=5.421010862e-32
+  voff={-2.486350287e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=3.627722941e-07 wvoff=-1.776356839e-21
+  nfactor={2.137127920e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-5.210855164e-6
+  eta0=0.08
+  etab=-0.07
+  u0=1.063746106e-02 lu0=-2.104594218e-8
+  ua=-9.116420042e-10 lua=3.285115641e-15
+  ub=1.339640455e-18 lub=-7.792683529e-24
+  uc=-1.046534774e-10 luc=-2.021399574e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=9.292141765e+04 lvsat=-2.556085955e-1
+  a0=1.626529302e+00 la0=-3.254408731e-6
+  ags=1.127437120e-01 lags=1.093860960e-8
+  a1=0.0
+  a2=1.083666533e+00 la2=-2.276004104e-6
+  b0=-1.709446520e-07 lb0=1.623339844e-12 pb0=6.776263578e-33
+  b1=5.452591595e-09 lb1=-4.138244049e-14
+  keta=3.421368674e-02 lketa=-2.173038039e-7
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-6.921953293e-02 lpclm=1.686371502e-06 wpclm=-1.110223025e-22
+  pdiblc1=0.39
+  pdiblc2=1.909636661e-03 lpdiblc2=-1.266443309e-8
+  pdiblcb=-0.225
+  drout=0.56
+  pscbe1=800000000.0
+  pscbe2=8.860770435e-09 lpscbe2=2.402531188e-14
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=-6.686266667e-11 lalpha0=1.338825943e-15
+  alpha1=-6.686266667e-11 lalpha1=1.338825943e-15
+  beta0=4.805292000e+01 lbeta0=-3.614830047e-4
* Gidl Induced Drain Leakage Model Parameters
+  agidl=1.354378090e-10 lagidl=-8.225743918e-16 pagidl=-6.617444900e-36
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.443915098e-01 lkt1=1.229746438e-7
+  kt2=-6.522345350e-02 lkt2=1.337061237e-7
+  at=7.716025872e+04 lat=-1.235502988e-1
+  ute=5.623649524e-01 lute=-1.292207756e-05 wute=-8.881784197e-22 pute=2.131628207e-26
+  ua1=3.775543044e-09 lua1=-3.374650014e-14
+  ub1=-2.648919653e-18 lub1=2.843379192e-23 pub1=-9.860761315e-44
+  uc1=-9.445040192e-11 luc1=1.294748875e-15 puc1=3.308722450e-36
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.155 pmos
* Model Flag Parameters
+  lmin=4.0e-06 lmax=8.0e-06 wmin=6.3e-07 wmax=6.4e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.036424065e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-2.719534781e-7
+  k1=4.604103273e-01 lk1=-5.535191579e-8
+  k2=3.111376993e-02 lk2=-4.835272375e-8
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-1.903188674e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-1.051285932e-7
+  nfactor={7.782034620e-01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=5.692502402e-6
+  eta0=0.08
+  etab=-0.07
+  u0=5.374816804e-03 lu0=2.117898927e-8
+  ua=-5.231013447e-10 lua=1.676518894e-16
+  ub=-7.890771535e-20 lub=3.589066086e-24
+  uc=-1.070071013e-10 luc=-1.329647545e-18
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=6.344101412e+04 lvsat=-1.907198821e-2
+  a0=1.169202877e+00 la0=4.149589883e-7
+  ags=4.476786908e-02 lags=5.563441444e-7
+  a1=0.0
+  a2=0.8
+  b0=1.333762438e-07 lb0=-8.183849488e-13
+  b1=-1.241682582e-09 lb1=1.232920225e-14
+  keta=7.540400483e-03 lketa=-3.290158170e-9
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-4.109336388e-01 lpclm=4.428121465e-06 ppclm=1.421085472e-26
+  pdiblc1=0.39
+  pdiblc2=2.318653116e-04 lpdiblc2=7.971988815e-10
+  pdiblcb=-0.225
+  drout=0.56
+  pscbe1=800000000.0
+  pscbe2=1.463489899e-08 lpscbe2=-2.230352405e-14
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=2.005880000e-10 lalpha0=-8.070698298e-16
+  alpha1=2.005880000e-10 lalpha1=-8.070698298e-16
+  beta0=-2.415876000e+01 lbeta0=2.179088540e-04 wbeta0=-2.842170943e-20
* Gidl Induced Drain Leakage Model Parameters
+  agidl=4.884466474e-11 lagidl=-1.277925667e-16
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.137901907e-01 lkt1=-1.225556520e-7
+  kt2=-3.851363950e-02 lkt2=-8.060060310e-8
+  at=2.230282385e+04 lat=3.165994270e-1
+  ute=-1.918426857e+00 lute=6.982605139e-06 pute=5.684341886e-26
+  ua1=-2.965829131e-09 lua1=2.034303433e-14 pua1=5.293955920e-35
+  ub1=2.930570959e-18 lub1=-1.633336259e-23 wub1=1.232595164e-38 pub1=4.930380658e-44
+  uc1=5.548297096e-10 luc1=-3.914763086e-15 wuc1=-8.271806126e-31 puc1=-3.308722450e-36
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.156 pmos
* Model Flag Parameters
+  lmin=2.0e-06 lmax=4.0e-06 wmin=6.3e-07 wmax=6.4e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.106065230e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=8.249143276e-9
+  k1=3.853412315e-01 lk1=2.466900923e-7
+  k2=4.064949326e-02 lk2=-8.671989728e-8
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=8.635279899e-01 ldsub=-1.221250938e-6
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.223718520e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=2.383723148e-8
+  nfactor={2.270962668e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-3.136441188e-7
+  eta0=1.604349200e-01 leta0=-3.236315093e-7
+  etab=-1.403173200e-01 letab=2.829231434e-7
+  u0=1.211265930e-02 lu0=-5.930854756e-9
+  ua=-1.308633256e-10 lua=-1.410525625e-15
+  ub=6.187485939e-19 lub=7.820319721e-25
+  uc=-1.338088641e-10 luc=1.065077811e-16
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=8.388955365e+04 lvsat=-1.013470960e-1
+  a0=1.400765170e+00 la0=-5.167365282e-7
+  ags=-4.432097709e-02 lags=9.147948988e-7
+  a1=0.0
+  a2=0.8
+  b0=-1.003353178e-07 lb0=1.219581936e-13
+  b1=1.451284080e-09 lb1=1.493997030e-15
+  keta=2.281093733e-02 lketa=-6.473146857e-08 wketa=1.110223025e-22
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=6.059902523e-01 lpclm=3.365078504e-7
+  pdiblc1=0.39
+  pdiblc2=4.185431636e-04 lpdiblc2=4.609681023e-11
+  pdiblcb=-4.273520000e-01 lpdiblcb=8.141673190e-7
+  drout=0.56
+  pscbe1=800000000.0
+  pscbe2=8.712478508e-09 lpscbe2=1.525453199e-15
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=-1.011760000e-10 lalpha0=4.070836595e-16
+  alpha1=-1.011760000e-10 lalpha1=4.070836595e-16
+  beta0=5.471942625e+01 lbeta0=-9.945910591e-5
* Gidl Induced Drain Leakage Model Parameters
+  agidl=1.634728531e-11 lagidl=2.961289373e-18
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.355286288e-01 lkt1=-3.509061145e-8
+  kt2=-6.321122536e-02 lkt2=1.877062754e-8
+  at=1.626547485e+05 lat=-2.481093488e-1
+  ute=-9.154724880e-02 lute=-3.678815031e-7
+  ua1=2.886961000e-09 lua1=-3.205783819e-15
+  ub1=-1.904818744e-18 lub1=3.121924585e-24
+  uc1=-8.771411122e-10 luc1=1.846800155e-15
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.157 pmos
* Model Flag Parameters
+  lmin=1.0e-06 lmax=2.0e-06 wmin=6.3e-07 wmax=6.4e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.118108631e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=3.261920430e-8
+  k1=5.064652470e-01 lk1=1.593224533e-9
+  k2=-2.759691298e-03 lk2=1.119455858e-9
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=2.600000202e-01 ldsub=-2.071113414e-14
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.052413704e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-1.082664065e-8
+  nfactor={2.508128773e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-7.935544749e-7
+  eta0=-5.005130400e-01 leta0=1.013809907e-06 weta0=4.440892099e-22 peta0=3.483324740e-27
+  etab=2.645421120e-04 letab=-1.547066255e-9
+  u0=1.145910416e-02 lu0=-4.608372862e-9
+  ua=-3.318390994e-10 lua=-1.003847127e-15
+  ub=7.130469709e-19 lub=5.912173203e-25
+  uc=-1.196469642e-10 luc=7.785089353e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=1.537394825e+04 lvsat=3.729560184e-2
+  a0=1.030938530e+00 la0=2.316150734e-7
+  ags=2.475687006e-01 lags=3.241502982e-7
+  a1=0.0
+  a2=0.8
+  b0=2.062768896e-08 lb0=-1.228128700e-13 pb0=-4.235164736e-34
+  b1=-2.754611245e-08 lb1=6.017080885e-14 wb1=5.293955920e-29 pb1=-1.058791184e-34
+  keta=-1.751182380e-02 lketa=1.686244502e-8
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=9.199174115e-01 lpclm=-2.987300348e-07 wpclm=-7.105427358e-21
+  pdiblc1=3.957940034e-01 lpdiblc1=-1.172428182e-8
+  pdiblc2=4.529136727e-04 lpdiblc2=-2.345260230e-11
+  pdiblcb=1.797040000e-01 lpdiblcb=-4.142226381e-7
+  drout=3.794864141e-01 ldrout=3.652728512e-7
+  pscbe1=800000000.0
+  pscbe2=9.769526283e-09 lpscbe2=-6.135041137e-16
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=4.643241089e+00 lbeta0=1.871056290e-6
* Gidl Induced Drain Leakage Model Parameters
+  agidl=2.528734937e-11 lagidl=-1.512910906e-17
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.260591597e-01 lkt1=-5.425227153e-8
+  kt2=-5.943725826e-02 lkt2=1.113392964e-8
+  at=2.804660864e+04 lat=2.427291432e-2
+  ute=5.196833265e-01 lute=-1.604718797e-6
+  ua1=3.076566596e-09 lua1=-3.589454534e-15
+  ub1=-1.607506698e-18 lub1=2.520307714e-24 pub1=6.162975822e-45
+  uc1=3.394859767e-12 luc1=6.501800488e-17
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=2.75e-6
+  sbref=2.74e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.158 pmos
* Model Flag Parameters
+  lmin=5.0e-07 lmax=1.0e-06 wmin=6.3e-07 wmax=6.4e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.104135008e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=1.831692178e-8
+  k1=5.845342661e-01 lk1=-7.831197791e-8
+  k2=-3.521780815e-02 lk2=3.434098762e-08 wk2=-1.110223025e-22 pk2=-4.163336342e-29
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=-5.148096000e-01 ldsub=7.930331218e-7
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.286451354e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=1.312758095e-8
+  nfactor={5.348218125e-01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.226164665e-6
+  eta0=9.944947238e-01 leta0=-5.163604397e-7
+  etab=-1.505565344e-03 letab=2.646741292e-10
+  u0=5.252885488e-03 lu0=1.743816071e-9
+  ua=-1.855248330e-09 lua=5.553926879e-16
+  ub=1.646936524e-18 lub=-3.646373153e-25 wub=-1.232595164e-38
+  uc=-3.861426543e-11 luc=-5.087694348e-18
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=5.284690706e+03 lvsat=4.762215872e-2
+  a0=1.406885884e+00 la0=-1.531745618e-7
+  ags=-1.537163707e-01 lags=7.348735944e-7
+  a1=0.0
+  a2=1.122324950e+00 la2=-3.299060332e-7
+  b0=-2.034000355e-07 lb0=1.064839866e-13
+  b1=6.395362368e-08 lb1=-3.348100107e-14
+  keta=4.345618449e-02 lketa=-4.553953082e-08 wketa=4.163336342e-23 pketa=7.632783294e-29
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=8.327961674e-01 lpclm=-2.095596990e-7
+  pdiblc1=7.135984939e-01 lpdiblc1=-3.370035339e-07 ppdiblc1=-1.776356839e-27
+  pdiblc2=3.879409928e-05 lpdiblc2=4.004070635e-10
+  pdiblcb=-0.225
+  drout=9.713112154e-01 ldrout=-2.404716693e-7
+  pscbe1=1.492842356e+09 lpscbe1=-7.091380085e+2
+  pscbe2=-6.308059837e-08 lpscbe2=7.395005547e-14 wpscbe2=-2.117582368e-28 ppscbe2=2.117582368e-34
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=4.407774865e+00 lbeta0=2.112060679e-6
* Gidl Induced Drain Leakage Model Parameters
+  agidl=2.547348960e-12 lagidl=8.145736160e-18
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.740229702e-01 lkt1=-5.160352257e-9
+  kt2=-3.705763611e-02 lkt2=-1.177206122e-8
+  at=2.219515839e+04 lat=3.026199068e-2
+  ute=-1.895801293e+00 lute=8.675780209e-07 pute=-7.105427358e-27
+  ua1=-2.625004008e-09 lua1=2.246217010e-15 pua1=6.617444900e-36
+  ub1=2.657182254e-18 lub1=-1.844686722e-24 wub1=1.232595164e-38
+  uc1=2.075025205e-10 luc1=-1.438902680e-16
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.75e-6
+  sbref=1.74e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.159 pmos
* Model Flag Parameters
+  lmin=2.5e-07 lmax=5.0e-07 wmin=6.3e-07 wmax=6.4e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.083600825e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=7.566866302e-9
+  k1=2.785842657e-01 lk1=8.185896632e-8
+  k2=9.078834505e-02 lk2=-3.162575371e-8
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=1.235674842e+00 ldsub=-1.233804932e-7
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={8.554790169e-02+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-1.513587578e-7
+  nfactor={3.380644558e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-2.636804585e-7
+  eta0=-5.189894481e-01 leta0=2.759787940e-07 weta0=1.554312234e-21 peta0=5.828670879e-28
+  etab=-2.015517863e-03 letab=5.316444720e-10
+  u0=1.182344359e-02 lu0=-1.696002504e-9
+  ua=-2.127182843e-10 lua=-3.045046414e-16
+  ub=5.497105694e-19 lub=2.097824166e-25
+  uc=-1.001292182e-10 luc=2.711661375e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=3.158190353e+04 lvsat=3.385504186e-2
+  a0=1.660440134e+00 la0=-2.859152828e-7
+  ags=9.698322770e-01 lags=1.466734064e-7
+  a1=0.0
+  a2=1.597024138e-01 la2=1.740461171e-7
+  b0=0.0
+  b1=0.0
+  keta=-5.647214109e-02 lketa=6.774946183e-9
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=2.085539131e-01 lpclm=1.172436059e-7
+  pdiblc1=-2.963791728e-01 lpdiblc1=1.917399742e-07 ppdiblc1=2.220446049e-28
+  pdiblc2=-7.700523841e-03 lpdiblc2=4.452094792e-09 wpdiblc2=1.387778781e-23 ppdiblc2=-1.040834086e-29
+  pdiblcb=-1.560512404e-01 lpdiblcb=-3.609605461e-8
+  drout=4.936971948e-01 ldrout=9.568822735e-9
+  pscbe1=-5.856554958e+08 lpscbe1=3.789971870e+02 ppscbe1=4.768371582e-19
+  pscbe2=1.540275727e-07 lpscbe2=-3.971041422e-14
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=7.930281860e+00 lbeta0=2.679578173e-7
* Gidl Induced Drain Leakage Model Parameters
+  agidl=3.791729715e-11 lagidl=-1.037113912e-17
+  bgidl=7.372237654e+08 lbgidl=1.375686143e+2
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.00074326333
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.5407449e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.413228120e-01 lkt1=-2.227953908e-8
+  kt2=-6.690804875e-02 lkt2=3.855226801e-9
+  at=9.325182934e+04 lat=-6.937597694e-3
+  ute=4.134590933e-01 lute=-3.413659765e-07 pute=8.881784197e-28
+  ua1=3.165106439e-09 lua1=-7.850216110e-16
+  ub1=-1.629143462e-18 lub1=3.992905164e-25
+  uc1=-3.393906100e-11 luc1=-1.749077126e-17
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.1e-6
+  sbref=1.1e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.160 pmos
* Model Flag Parameters
+  lmin=1.8e-07 lmax=2.5e-07 wmin=6.3e-07 wmax=6.4e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.012266656e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-1.194445551e-8
+  k1=-8.579247482e-01 lk1=3.927169118e-7
+  k2=5.167953973e-01 lk2=-1.481472026e-07 wk2=1.332267630e-21 pk2=-1.110223025e-28
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=1.803960266e+00 ldsub=-2.788179225e-7
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-7.309221625e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=7.196213411e-8
+  nfactor={2.983359543e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.550150614e-7
+  eta0=4.900000008e-01 leta0=-7.096190302e-17
+  etab=2.195759126e-03 letab=-6.202240101e-10 wetab=-1.734723476e-24 petab=-1.301042607e-30
+  u0=1.425126466e-02 lu0=-2.360060124e-9
+  ua=1.721124685e-09 lua=-8.334493704e-16
+  ub=-8.156452782e-19 lub=5.832345480e-25
+  uc=3.489543344e-11 luc=-9.815328983e-18 wuc=7.754818243e-32
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=3.617753405e+05 lvsat=-5.645946701e-2
+  a0=-1.466462483e-01 la0=2.083589844e-7
+  ags=2.250598986e+00 lags=-2.036419039e-7
+  a1=0.0
+  a2=9.336249622e-01 la2=-3.763717830e-8
+  b0=0.0
+  b1=0.0
+  keta=-8.737025015e-02 lketa=1.522619697e-08 pketa=-1.110223025e-28
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=6.849679741e-01 lpclm=-1.306516802e-8
+  pdiblc1=5.487137542e-01 lpdiblc1=-3.940984321e-8
+  pdiblc2=2.991525761e-02 lpdiblc2=-5.836573751e-9
+  pdiblcb=2.186325871e+00 lpdiblcb=-6.767830420e-7
+  drout=-8.416446543e-01 ldrout=3.748115253e-7
+  pscbe1=7.998956542e+08 lpscbe1=2.123647450e-2
+  pscbe2=1.957358274e-08 lpscbe2=-2.934558902e-15
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=1.052647787e+01 lbeta0=-4.421537155e-7
* Gidl Induced Drain Leakage Model Parameters
+  agidl=9.578483481e-15 lagidl=-2.619906802e-21
+  bgidl=1.938486425e+09 lbgidl=-1.910007484e+2
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.00074326333
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.5407449e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=2.438598179e-01 lkt1=-2.096906920e-7
+  kt2=-5.870698811e-02 lkt2=1.612072696e-9
+  at=2.121185134e+05 lat=-3.945001311e-2
+  ute=-1.856079955e+00 lute=2.793983441e-07 wute=1.421085472e-20
+  ua1=1.352904843e-10 lua1=4.369364895e-17
+  ub1=-3.305422621e-19 lub1=4.409711620e-26
+  uc1=-2.972920545e-10 luc1=5.454153952e-17 puc1=-4.135903063e-37
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.1e-6
+  sbref=1.1e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.161 pmos
* Model Flag Parameters
+  lmin=1.5e-07 lmax=1.8e-07 wmin=6.3e-07 wmax=6.4e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-2.026e-8
+  vth0={1.302789072e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-5.234582635e-07 wvth0=-1.474575643e-06 pvth0=3.251734208e-13
+  k1=2.666255590e-01 lk1=1.775346723e-07 wk1=5.001690142e-07 pk1=-1.102972710e-13
+  k2=-6.537104039e+00 lk2=1.395003984e-06 wk2=3.930151099e-06 pk2=-8.666769204e-13
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=-5.155565786e+00 ldsub=1.232607137e-06 wdsub=3.472629566e-06 pdsub=-7.657842719e-13
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={3.155670232e+01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-7.042093830e-06 wvoff=-1.983972314e-05 pvoff=4.375055746e-12
+  nfactor={3.999130933e+02+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-8.769890834e-05 wnfactor=-2.470745340e-04 pnfactor=5.448487624e-11
+  eta0=-1.093665024e+01 leta0=2.519804911e-06 weta0=7.099057850e-06 peta0=-1.565484237e-12
+  etab=-6.496892491e-01 letab=1.430816508e-07 wetab=4.031045463e-07 petab=-8.889261456e-14
+  u0=-5.499844497e-02 lu0=1.271375032e-08 wu0=3.581799883e-08 pu0=-7.898585101e-15
+  ua=4.539382406e-09 lua=-1.524549484e-15 wua=-4.295120371e-15 pua=9.471599442e-22
+  ub=-2.519919023e-19 lub=5.076552140e-25 wub=1.430219393e-24 pub=-3.153919806e-31
+  uc=4.871909564e-10 luc=-1.103754109e-16 wuc=-3.109611420e-16 puc=6.857315104e-23
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=1.450144756e+07 lvsat=-3.179256036e+00 wvsat=-8.956932479e+00 pvsat=1.975182750e-6
+  a0=5.978140540e+00 la0=-1.124874798e-06 wa0=-3.169114070e-06 pa0=6.988530347e-13
+  ags=1.250000067e+00 lags=-1.292610818e-14 wags=-2.607123406e-15 pags=5.749143384e-22
+  a1=0.0
+  a2=8.547183238e+00 la2=-1.719722878e-06 wa2=-4.844983061e-06 pa2=1.068415665e-12
+  b0=0.0
+  b1=0.0
+  keta=1.996439956e+00 lketa=-4.430237873e-07 wketa=-1.248132918e-06 pketa=2.752382710e-13
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=6.633270215e-01 lpclm=-9.384236998e-09 wpclm=-2.643824011e-08 ppclm=5.830160708e-15
+  pdiblc1=-6.508220492e+00 lpdiblc1=1.513493398e-06 wpdiblc1=4.263972085e-06 ppdiblc1=-9.402911241e-13
+  pdiblc2=3.424791438e-02 lpdiblc2=-7.279539492e-09 wpdiblc2=-2.050868406e-08 ppdiblc2=4.522575010e-15
+  pdiblcb=3.875064344e+01 lpdiblcb=-8.796477954e-06 wpdiblcb=-2.478235740e-05 ppdiblcb=5.465005455e-12
+  drout=1.000000053e+00 ldrout=-5.914387202e-15 wdrout=8.551069186e-14 pdrout=-1.885682366e-20
+  pscbe1=7.861069041e+07 lpscbe1=1.590807706e+02 wpscbe1=4.481789794e+02 ppscbe1=-9.883242854e-5
+  pscbe2=1.562207896e-07 lpscbe2=-3.331312430e-14 wpscbe2=-9.385321921e-14 ppscbe2=2.069651190e-20
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=-5.199897891e+00 lbeta0=2.988893623e-06 wbeta0=8.420623045e-06 pbeta0=-1.856915794e-12
* Gidl Induced Drain Leakage Model Parameters
+  agidl=-2.421667034e-14 lagidl=4.613760032e-21
+  bgidl=1.000000428e+09 lbgidl=-8.465629578e-05 wbgidl=-6.635260010e-05 pbgidl=1.463207245e-11
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-1.106e-8
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=7.730602693e+01 lkt1=-1.722095522e-05 wkt1=-4.851667560e-05 pkt1=1.069889730e-11
+  kt2=-1.639495691e+00 lkt2=3.503422538e-07 wkt2=9.870206947e-07 pkt2=-2.176578036e-13
+  at=1.423147657e+06 lat=-3.098014146e-01 wat=-8.728049138e-01 pat=1.924709396e-7
+  ute=1.151482381e+01 lute=-2.645815245e-06 wute=-7.454067500e-06 pute=1.643770965e-12
+  ua1=1.510530450e-08 lua1=-3.253844117e-15 wua1=-9.167069095e-15 pua1=2.021522077e-21
+  ub1=-2.011491469e-17 lub1=4.410630350e-24 wub1=1.242608853e-23 pub1=-2.740201043e-30
+  uc1=-4.826448999e-10 luc1=9.997139693e-17 wuc1=2.816498738e-16 puc1=-6.210943017e-23
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.04e-6
+  sbref=1.04e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.162 pmos
* Model Flag Parameters
+  lmin=2.0e-05 lmax=0.0001 wmin=5.5e-07 wmax=6.3e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.126311+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+  k1=0.43165561
+  k2=0.026980026
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=3.2465718e-7
+  voff={-0.23051772+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.8768912+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+  eta0=0.08
+  etab=-0.07
+  u0=0.0095864
+  ua=-7.4757916e-10
+  ub=9.5046395e-19
+  uc=-1.0566299e-10
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=80156.0
+  a0=1.464
+  ags=0.11329
+  a1=0.0
+  a2=0.97
+  b0=-8.9873e-8
+  b1=3.3859e-9
+  keta=0.023361259
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=0.015
+  pdiblc1=0.39
+  pdiblc2=0.0012771588
+  pdiblcb=-0.225
+  drout=0.56
+  pscbe1=800000000.0
+  pscbe2=1.0060625e-8
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=0.0
+  alpha1=0.0
+  beta0=30.0
* Gidl Induced Drain Leakage Model Parameters
+  agidl=9.43573999999999e-11
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-0.43825
+  kt2=-0.058546
+  at=70990.0
+  ute=-0.08298
+  ua1=2.0902e-9
+  ub1=-1.2289e-18
+  uc1=-2.9789e-11
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.163 pmos
* Model Flag Parameters
+  lmin=8.0e-06 lmax=2.0e-05 wmin=5.5e-07 wmax=6.3e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.163749012e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=7.496407775e-07 wvth0=8.881784197e-22
+  k1=4.170420989e-01 lk1=2.926139320e-7
+  k2=2.824548822e-02 lk2=-2.533900806e-8
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=-6.144535039e-06 lcit=1.295359998e-10 wcit=8.470329473e-28 pcit=4.743384505e-32
+  voff={-2.486350287e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=3.627722941e-7
+  nfactor={2.137127920e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-5.210855164e-6
+  eta0=0.08
+  etab=-0.07
+  u0=1.063746106e-02 lu0=-2.104594218e-8
+  ua=-9.116420042e-10 lua=3.285115641e-15
+  ub=1.339640455e-18 lub=-7.792683529e-24
+  uc=-1.046534774e-10 luc=-2.021399574e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=9.292141765e+04 lvsat=-2.556085955e-1
+  a0=1.626529302e+00 la0=-3.254408731e-6
+  ags=1.127437120e-01 lags=1.093860960e-8
+  a1=0.0
+  a2=1.083666533e+00 la2=-2.276004104e-6
+  b0=-1.709446520e-07 lb0=1.623339844e-12
+  b1=5.452591595e-09 lb1=-4.138244049e-14
+  keta=3.421368674e-02 lketa=-2.173038039e-07 wketa=-2.775557562e-23
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-6.921953293e-02 lpclm=1.686371502e-06 wpclm=-1.387778781e-23 ppclm=-3.330669074e-28
+  pdiblc1=0.39
+  pdiblc2=1.909636661e-03 lpdiblc2=-1.266443309e-8
+  pdiblcb=-0.225
+  drout=0.56
+  pscbe1=800000000.0
+  pscbe2=8.860770435e-09 lpscbe2=2.402531188e-14
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=-6.686266667e-11 lalpha0=1.338825943e-15
+  alpha1=-6.686266667e-11 lalpha1=1.338825943e-15
+  beta0=4.805292000e+01 lbeta0=-3.614830047e-4
* Gidl Induced Drain Leakage Model Parameters
+  agidl=1.354378090e-10 lagidl=-8.225743918e-16
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.443915098e-01 lkt1=1.229746438e-7
+  kt2=-6.522345350e-02 lkt2=1.337061237e-07 wkt2=-5.551115123e-23
+  at=7.716025872e+04 lat=-1.235502988e-1
+  ute=5.623649524e-01 lute=-1.292207756e-05 wute=-1.110223025e-22 pute=-3.552713679e-27
+  ua1=3.775543044e-09 lua1=-3.374650014e-14 wua1=1.654361225e-30
+  ub1=-2.648919653e-18 lub1=2.843379192e-23
+  uc1=-9.445040192e-11 luc1=1.294748875e-15 wuc1=2.584939414e-32
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.164 pmos
* Model Flag Parameters
+  lmin=4.0e-06 lmax=8.0e-06 wmin=5.5e-07 wmax=6.3e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.036424065e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-2.719534781e-7
+  k1=4.604103273e-01 lk1=-5.535191579e-8
+  k2=3.111376993e-02 lk2=-4.835272375e-8
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-1.903188674e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-1.051285932e-7
+  nfactor={7.782034620e-01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=5.692502402e-6
+  eta0=0.08
+  etab=-0.07
+  u0=5.374816804e-03 lu0=2.117898927e-8
+  ua=-5.231013447e-10 lua=1.676518894e-16
+  ub=-7.890771535e-20 lub=3.589066086e-24 pub=-1.540743956e-45
+  uc=-1.070071013e-10 luc=-1.329647545e-18
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=6.344101412e+04 lvsat=-1.907198821e-2
+  a0=1.169202877e+00 la0=4.149589883e-7
+  ags=4.476786908e-02 lags=5.563441444e-7
+  a1=0.0
+  a2=0.8
+  b0=1.333762438e-07 lb0=-8.183849488e-13 wb0=5.293955920e-29
+  b1=-1.241682582e-09 lb1=1.232920225e-14 wb1=-4.135903063e-31 pb1=1.654361225e-36
+  keta=7.540400483e-03 lketa=-3.290158170e-9
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-4.109336388e-01 lpclm=4.428121465e-6
+  pdiblc1=0.39
+  pdiblc2=2.318653116e-04 lpdiblc2=7.971988815e-10
+  pdiblcb=-0.225
+  drout=0.56
+  pscbe1=800000000.0
+  pscbe2=1.463489899e-08 lpscbe2=-2.230352405e-14
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=2.005880000e-10 lalpha0=-8.070698298e-16
+  alpha1=2.005880000e-10 lalpha1=-8.070698298e-16
+  beta0=-2.415876000e+01 lbeta0=2.179088540e-04 wbeta0=3.552713679e-21 pbeta0=2.842170943e-26
* Gidl Induced Drain Leakage Model Parameters
+  agidl=4.884466474e-11 lagidl=-1.277925667e-16
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.137901907e-01 lkt1=-1.225556520e-7
+  kt2=-3.851363950e-02 lkt2=-8.060060310e-8
+  at=2.230282385e+04 lat=3.165994270e-1
+  ute=-1.918426857e+00 lute=6.982605139e-6
+  ua1=-2.965829131e-09 lua1=2.034303433e-14 wua1=4.135903063e-31 pua1=-4.963083675e-36
+  ub1=2.930570959e-18 lub1=-1.633336259e-23
+  uc1=5.548297096e-10 luc1=-3.914763086e-15 puc1=1.240770919e-36
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.165 pmos
* Model Flag Parameters
+  lmin=2.0e-06 lmax=4.0e-06 wmin=5.5e-07 wmax=6.3e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.106065230e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=8.249143277e-9
+  k1=3.853412315e-01 lk1=2.466900923e-7
+  k2=4.064949326e-02 lk2=-8.671989728e-8
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=8.635279899e-01 ldsub=-1.221250938e-6
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.223718520e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=2.383723148e-8
+  nfactor={2.270962668e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-3.136441188e-7
+  eta0=1.604349200e-01 leta0=-3.236315093e-7
+  etab=-1.403173200e-01 letab=2.829231434e-7
+  u0=1.211265930e-02 lu0=-5.930854756e-9
+  ua=-1.308633256e-10 lua=-1.410525625e-15
+  ub=6.187485939e-19 lub=7.820319721e-25
+  uc=-1.338088641e-10 luc=1.065077811e-16
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=8.388955365e+04 lvsat=-1.013470960e-1
+  a0=1.400765170e+00 la0=-5.167365282e-7
+  ags=-4.432097709e-02 lags=9.147948988e-7
+  a1=0.0
+  a2=0.8
+  b0=-1.003353178e-07 lb0=1.219581936e-13
+  b1=1.451284080e-09 lb1=1.493997030e-15
+  keta=2.281093733e-02 lketa=-6.473146857e-08 wketa=-6.938893904e-24 pketa=2.775557562e-29
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=6.059902523e-01 lpclm=3.365078504e-7
+  pdiblc1=0.39
+  pdiblc2=4.185431636e-04 lpdiblc2=4.609681023e-11
+  pdiblcb=-4.273520000e-01 lpdiblcb=8.141673190e-7
+  drout=0.56
+  pscbe1=800000000.0
+  pscbe2=8.712478508e-09 lpscbe2=1.525453199e-15
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=-1.011760000e-10 lalpha0=4.070836595e-16
+  alpha1=-1.011760000e-10 lalpha1=4.070836595e-16
+  beta0=5.471942625e+01 lbeta0=-9.945910591e-05 wbeta0=2.842170943e-20
* Gidl Induced Drain Leakage Model Parameters
+  agidl=1.634728531e-11 lagidl=2.961289373e-18
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.355286288e-01 lkt1=-3.509061145e-8
+  kt2=-6.321122536e-02 lkt2=1.877062754e-8
+  at=1.626547485e+05 lat=-2.481093488e-1
+  ute=-9.154724880e-02 lute=-3.678815031e-7
+  ua1=2.886961000e-09 lua1=-3.205783819e-15
+  ub1=-1.904818744e-18 lub1=3.121924585e-24
+  uc1=-8.771411122e-10 luc1=1.846800155e-15
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.166 pmos
* Model Flag Parameters
+  lmin=1.0e-06 lmax=2.0e-06 wmin=5.5e-07 wmax=6.3e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.118108631e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=3.261920430e-8
+  k1=5.064652470e-01 lk1=1.593224533e-9
+  k2=-2.759691298e-03 lk2=1.119455858e-9
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=2.600000202e-01 ldsub=-2.071113236e-14
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.052413704e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-1.082664065e-8
+  nfactor={2.508128773e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-7.935544749e-7
+  eta0=-5.005130400e-01 leta0=1.013809907e-06 weta0=-1.552577511e-22 peta0=-2.151057110e-28
+  etab=2.645421120e-04 letab=-1.547066255e-9
+  u0=1.145910416e-02 lu0=-4.608372862e-9
+  ua=-3.318390994e-10 lua=-1.003847127e-15
+  ub=7.130469709e-19 lub=5.912173203e-25
+  uc=-1.196469642e-10 luc=7.785089353e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=1.537394825e+04 lvsat=3.729560184e-2
+  a0=1.030938530e+00 la0=2.316150734e-7
+  ags=2.475687006e-01 lags=3.241502982e-7
+  a1=0.0
+  a2=0.8
+  b0=2.062768896e-08 lb0=-1.228128700e-13 pb0=5.293955920e-35
+  b1=-2.754611245e-08 lb1=6.017080885e-14 wb1=6.617444900e-30 pb1=-9.926167351e-36
+  keta=-1.751182380e-02 lketa=1.686244502e-8
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=9.199174115e-01 lpclm=-2.987300348e-7
+  pdiblc1=3.957940034e-01 lpdiblc1=-1.172428182e-8
+  pdiblc2=4.529136727e-04 lpdiblc2=-2.345260230e-11
+  pdiblcb=1.797040000e-01 lpdiblcb=-4.142226381e-07 ppdiblcb=8.326672685e-29
+  drout=3.794864141e-01 ldrout=3.652728512e-7
+  pscbe1=800000000.0
+  pscbe2=9.769526283e-09 lpscbe2=-6.135041137e-16
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=4.643241089e+00 lbeta0=1.871056290e-6
* Gidl Induced Drain Leakage Model Parameters
+  agidl=2.528734937e-11 lagidl=-1.512910906e-17
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.260591597e-01 lkt1=-5.425227153e-8
+  kt2=-5.943725826e-02 lkt2=1.113392964e-8
+  at=2.804660864e+04 lat=2.427291432e-2
+  ute=5.196833265e-01 lute=-1.604718797e-06 pute=-4.440892099e-28
+  ua1=3.076566596e-09 lua1=-3.589454534e-15
+  ub1=-1.607506698e-18 lub1=2.520307714e-24 wub1=3.851859889e-40
+  uc1=3.394859767e-12 luc1=6.501800488e-17
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=2.75e-6
+  sbref=2.74e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.167 pmos
* Model Flag Parameters
+  lmin=5.0e-07 lmax=1.0e-06 wmin=5.5e-07 wmax=6.3e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.104135008e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=1.831692178e-8
+  k1=5.845342661e-01 lk1=-7.831197791e-8
+  k2=-3.521780815e-02 lk2=3.434098762e-08 wk2=8.673617380e-24 pk2=4.336808690e-30
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=-5.148096000e-01 ldsub=7.930331218e-7
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.286451354e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=1.312758095e-8
+  nfactor={5.348218125e-01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.226164665e-6
+  eta0=9.944947238e-01 leta0=-5.163604397e-7
+  etab=-1.505565344e-03 letab=2.646741292e-10
+  u0=5.252885488e-03 lu0=1.743816071e-9
+  ua=-1.855248330e-09 lua=5.553926879e-16
+  ub=1.646936524e-18 lub=-3.646373153e-25
+  uc=-3.861426543e-11 luc=-5.087694348e-18
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=5.284690706e+03 lvsat=4.762215872e-2
+  a0=1.406885884e+00 la0=-1.531745618e-7
+  ags=-1.537163707e-01 lags=7.348735944e-7
+  a1=0.0
+  a2=1.122324950e+00 la2=-3.299060332e-7
+  b0=-2.034000355e-07 lb0=1.064839866e-13
+  b1=6.395362368e-08 lb1=-3.348100107e-14
+  keta=4.345618449e-02 lketa=-4.553953082e-08 wketa=1.214306433e-23 pketa=5.204170428e-30
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=8.327961674e-01 lpclm=-2.095596990e-7
+  pdiblc1=7.135984939e-01 lpdiblc1=-3.370035339e-7
+  pdiblc2=3.879409928e-05 lpdiblc2=4.004070635e-10
+  pdiblcb=-0.225
+  drout=9.713112154e-01 ldrout=-2.404716693e-7
+  pscbe1=1.492842356e+09 lpscbe1=-7.091380085e+2
+  pscbe2=-6.308059837e-08 lpscbe2=7.395005547e-14 wpscbe2=-1.323488980e-29 ppscbe2=-1.985233470e-35
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=4.407774865e+00 lbeta0=2.112060679e-6
* Gidl Induced Drain Leakage Model Parameters
+  agidl=2.547348960e-12 lagidl=8.145736160e-18
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.740229702e-01 lkt1=-5.160352257e-9
+  kt2=-3.705763611e-02 lkt2=-1.177206122e-8
+  at=2.219515839e+04 lat=3.026199068e-2
+  ute=-1.895801293e+00 lute=8.675780209e-7
+  ua1=-2.625004008e-09 lua1=2.246217010e-15 pua1=-8.271806126e-37
+  ub1=2.657182254e-18 lub1=-1.844686722e-24 pub1=7.703719778e-46
+  uc1=2.075025205e-10 luc1=-1.438902680e-16
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.75e-6
+  sbref=1.74e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.168 pmos
* Model Flag Parameters
+  lmin=2.5e-07 lmax=5.0e-07 wmin=5.5e-07 wmax=6.3e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.083600825e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=7.566866302e-9
+  k1=2.785842657e-01 lk1=8.185896632e-8
+  k2=9.078834505e-02 lk2=-3.162575371e-8
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=1.235674842e+00 ldsub=-1.233804932e-7
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={8.554790169e-02+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-1.513587578e-7
+  nfactor={3.380644558e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-2.636804585e-7
+  eta0=-5.189894481e-01 leta0=2.759787940e-07 weta0=-6.938893904e-23 peta0=9.367506770e-29
+  etab=-2.015517863e-03 letab=5.316444720e-10
+  u0=1.182344359e-02 lu0=-1.696002504e-9
+  ua=-2.127182843e-10 lua=-3.045046414e-16
+  ub=5.497105694e-19 lub=2.097824166e-25
+  uc=-1.001292182e-10 luc=2.711661375e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=3.158190353e+04 lvsat=3.385504186e-2
+  a0=1.660440134e+00 la0=-2.859152828e-7
+  ags=9.698322770e-01 lags=1.466734064e-7
+  a1=0.0
+  a2=1.597024138e-01 la2=1.740461171e-7
+  b0=0.0
+  b1=0.0
+  keta=-5.647214109e-02 lketa=6.774946183e-9
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=2.085539131e-01 lpclm=1.172436059e-7
+  pdiblc1=-2.963791728e-01 lpdiblc1=1.917399742e-07 ppdiblc1=2.775557562e-29
+  pdiblc2=-7.700523841e-03 lpdiblc2=4.452094792e-09 wpdiblc2=-2.602085214e-24 ppdiblc2=-4.336808690e-31
+  pdiblcb=-1.560512404e-01 lpdiblcb=-3.609605461e-8
+  drout=4.936971948e-01 ldrout=9.568822735e-9
+  pscbe1=-5.856554958e+08 lpscbe1=3.789971870e+2
+  pscbe2=1.540275727e-07 lpscbe2=-3.971041422e-14
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=7.930281860e+00 lbeta0=2.679578173e-7
* Gidl Induced Drain Leakage Model Parameters
+  agidl=3.791729715e-11 lagidl=-1.037113912e-17
+  bgidl=7.372237654e+08 lbgidl=1.375686143e+2
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.00074326333
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.5407449e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.413228120e-01 lkt1=-2.227953908e-8
+  kt2=-6.690804875e-02 lkt2=3.855226801e-9
+  at=9.325182934e+04 lat=-6.937597694e-3
+  ute=4.134590933e-01 lute=-3.413659765e-7
+  ua1=3.165106439e-09 lua1=-7.850216110e-16
+  ub1=-1.629143462e-18 lub1=3.992905164e-25
+  uc1=-3.393906100e-11 luc1=-1.749077126e-17
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.1e-6
+  sbref=1.1e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.169 pmos
* Model Flag Parameters
+  lmin=1.8e-07 lmax=2.5e-07 wmin=5.5e-07 wmax=6.3e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.012266656e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-1.194445551e-8
+  k1=-8.579247482e-01 lk1=3.927169118e-7
+  k2=5.167953973e-01 lk2=-1.481472026e-07 wk2=-2.220446049e-22 pk2=4.163336342e-29
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=1.803960266e+00 ldsub=-2.788179225e-7
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-7.309221625e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=7.196213411e-8
+  nfactor={2.983359543e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.550150614e-7
+  eta0=4.900000008e-01 leta0=-7.095968257e-17
+  etab=2.195759126e-03 letab=-6.202240101e-10 wetab=2.168404345e-25 petab=-2.710505431e-32
+  u0=1.425126466e-02 lu0=-2.360060124e-9
+  ua=1.721124685e-09 lua=-8.334493704e-16
+  ub=-8.156452782e-19 lub=5.832345480e-25
+  uc=3.489543344e-11 luc=-9.815328983e-18 wuc=-3.231174268e-33 puc=-1.211690350e-39
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=3.617753405e+05 lvsat=-5.645946701e-2
+  a0=-1.466462483e-01 la0=2.083589844e-7
+  ags=2.250598986e+00 lags=-2.036419039e-7
+  a1=0.0
+  a2=9.336249622e-01 la2=-3.763717830e-8
+  b0=0.0
+  b1=0.0
+  keta=-8.737025015e-02 lketa=1.522619697e-8
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=6.849679741e-01 lpclm=-1.306516802e-8
+  pdiblc1=5.487137542e-01 lpdiblc1=-3.940984321e-8
+  pdiblc2=2.991525761e-02 lpdiblc2=-5.836573751e-9
+  pdiblcb=2.186325871e+00 lpdiblcb=-6.767830420e-07 wpdiblcb=-8.881784197e-22 ppdiblcb=-2.220446049e-28
+  drout=-8.416446543e-01 ldrout=3.748115253e-7
+  pscbe1=7.998956542e+08 lpscbe1=2.123647450e-2
+  pscbe2=1.957358274e-08 lpscbe2=-2.934558902e-15
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=1.052647787e+01 lbeta0=-4.421537155e-7
* Gidl Induced Drain Leakage Model Parameters
+  agidl=9.578483481e-15 lagidl=-2.619906802e-21
+  bgidl=1.938486425e+09 lbgidl=-1.910007484e+2
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.00074326333
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.5407449e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=2.438598179e-01 lkt1=-2.096906920e-7
+  kt2=-5.870698811e-02 lkt2=1.612072696e-9
+  at=2.121185134e+05 lat=-3.945001311e-2
+  ute=-1.856079955e+00 lute=2.793983441e-7
+  ua1=1.352904843e-10 lua1=4.369364895e-17
+  ub1=-3.305422621e-19 lub1=4.409711620e-26
+  uc1=-2.972920545e-10 luc1=5.454153952e-17
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.1e-6
+  sbref=1.1e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.170 pmos
* Model Flag Parameters
+  lmin=1.5e-07 lmax=1.8e-07 wmin=5.5e-07 wmax=6.3e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-2.026e-8
+  vth0={-1.378297177e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=6.777487612e-08 wvth0=1.642973108e-07 pvth0=-3.623084298e-14
+  k1=2.666255684e-01 lk1=1.775346702e-07 wk1=5.001690085e-07 pk1=-1.102972697e-13
+  k2=3.635604738e-01 lk2=-1.267305545e-07 wk2=-2.880318992e-07 pk2=6.351679442e-14
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=-5.155565835e+00 ldsub=1.232607147e-06 wdsub=3.472629596e-06 pdsub=-7.657842784e-13
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-3.651044768e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=7.219185591e-07 wvoff=1.681786844e-06 pvoff=-3.708676349e-13
+  nfactor={-5.199573980e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.195602754e-05 wnfactor=2.916468220e-05 pnfactor=-6.431395718e-12
+  eta0=-1.093665135e+01 leta0=2.519805157e-06 weta0=7.099058531e-06 peta0=-1.565484387e-12
+  etab=-6.496891861e-01 letab=1.430816369e-07 wetab=4.031045078e-07 petab=-8.889260606e-14
+  u0=3.313310763e-02 lu0=-6.721019662e-09 wu0=-1.805435160e-08 pu0=3.981345614e-15
+  ua=4.539381566e-09 lua=-1.524549299e-15 wua=-4.295119858e-15 pua=9.471598310e-22
+  ub=-2.519914808e-19 lub=5.076551211e-25 wub=1.430219136e-24 pub=-3.153919238e-31
+  uc=4.871909543e-10 luc=-1.103754104e-16 wuc=-3.109611408e-16 puc=6.857315077e-23
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=-1.316505234e+06 lvsat=3.089189131e-01 wvsat=7.121391582e-01 pvsat=-1.570409272e-7
+  a0=5.978140941e+00 la0=-1.124874887e-06 wa0=-3.169114315e-06 pa0=6.988530888e-13
+  ags=1.250000062e+00 lags=-1.188502452e-14 wags=2.786819664e-16 pags=-6.145484122e-23
+  a1=0.0
+  a2=8.547183572e+00 la2=-1.719722952e-06 wa2=-4.844983266e-06 pa2=1.068415710e-12
+  b0=0.0
+  b1=0.0
+  keta=1.996439835e+00 lketa=-4.430237606e-07 wketa=-1.248132844e-06 pketa=2.752382547e-13
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=6.633270275e-01 lpclm=-9.384238313e-09 wpclm=-2.643824375e-08 ppclm=5.830161512e-15
+  pdiblc1=-6.508220570e+00 lpdiblc1=1.513493415e-06 wpdiblc1=4.263972132e-06 ppdiblc1=-9.402911346e-13
+  pdiblc2=3.424790847e-02 lpdiblc2=-7.279538190e-09 wpdiblc2=-2.050868045e-08 ppdiblc2=4.522574214e-15
+  pdiblcb=3.875064748e+01 lpdiblcb=-8.796478846e-06 wpdiblcb=-2.478235988e-05 ppdiblcb=5.465006000e-12
+  drout=1.000000208e+00 ldrout=-4.006034438e-14 wdrout=-9.140411095e-15 pdrout=2.015642764e-21
+  pscbe1=7.861074015e+07 lpscbe1=1.590807596e+02 wpscbe1=4.481789490e+02 ppscbe1=-9.883242183e-5
+  pscbe2=1.562207629e-07 lpscbe2=-3.331311841e-14 wpscbe2=-9.385320288e-14 ppscbe2=2.069650830e-20
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=-5.199898492e+00 lbeta0=2.988893756e-06 wbeta0=8.420623412e-06 pbeta0=-1.856915875e-12
* Gidl Induced Drain Leakage Model Parameters
+  agidl=-2.421667034e-14 lagidl=4.613760032e-21
+  bgidl=1.000000307e+09 lbgidl=-5.816053009e-05 wbgidl=7.092559814e-06 pbgidl=-1.564051628e-12
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-1.106e-8
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-6.047618253e+00 lkt1=1.160190615e-06 wkt1=2.435073798e-06 pkt1=-5.369824740e-13
+  kt2=-1.639495540e+00 lkt2=3.503422204e-07 wkt2=9.870206023e-07 pkt2=-2.176577832e-13
+  at=1.423147570e+06 lat=-3.098013954e-01 wat=-8.728048606e-01 pat=1.924709279e-7
+  ute=1.151482466e+01 lute=-2.645815434e-06 wute=-7.454068023e-06 pute=1.643771080e-12
+  ua1=1.510530841e-08 lua1=-3.253844978e-15 wua1=-9.167071482e-15 pua1=2.021522603e-21
+  ub1=-2.011491045e-17 lub1=4.410629417e-24 wub1=1.242608594e-23 pub1=-2.740200472e-30
+  uc1=-4.826449106e-10 luc1=9.997139928e-17 wuc1=2.816498803e-16 puc1=-6.210943161e-23
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.04e-6
+  sbref=1.04e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.171 pmos
* Model Flag Parameters
+  lmin=2.0e-05 lmax=0.0001 wmin=5.4e-07 wmax=5.5e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.126311+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+  k1=0.43165561
+  k2=0.026980026
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=3.2465718e-7
+  voff={-0.23051772+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.8768912+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+  eta0=0.08
+  etab=-0.07
+  u0=0.0095864
+  ua=-7.4757916e-10
+  ub=9.5046395e-19
+  uc=-1.0566299e-10
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=80156.0
+  a0=1.464
+  ags=0.11329
+  a1=0.0
+  a2=0.97
+  b0=-8.9873e-8
+  b1=3.3859e-9
+  keta=0.023361259
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=0.015
+  pdiblc1=0.39
+  pdiblc2=0.0012771588
+  pdiblcb=-0.225
+  drout=0.56
+  pscbe1=800000000.0
+  pscbe2=1.0060625e-8
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=0.0
+  alpha1=0.0
+  beta0=30.0
* Gidl Induced Drain Leakage Model Parameters
+  agidl=9.43573999999999e-11
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-0.43825
+  kt2=-0.058546
+  at=70990.0
+  ute=-0.08298
+  ua1=2.0902e-9
+  ub1=-1.2289e-18
+  uc1=-2.9789e-11
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.172 pmos
* Model Flag Parameters
+  lmin=8.0e-06 lmax=2.0e-05 wmin=5.4e-07 wmax=5.5e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.163749012e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=7.496407775e-7
+  k1=4.170420989e-01 lk1=2.926139320e-7
+  k2=2.824548822e-02 lk2=-2.533900806e-8
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=-6.144535039e-06 lcit=1.295359998e-10 wcit=5.082197684e-27 pcit=2.710505431e-32
+  voff={-2.486350287e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=3.627722941e-7
+  nfactor={2.137127920e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-5.210855164e-6
+  eta0=0.08
+  etab=-0.07
+  u0=1.063746106e-02 lu0=-2.104594218e-8
+  ua=-9.116420042e-10 lua=3.285115641e-15
+  ub=1.339640455e-18 lub=-7.792683529e-24
+  uc=-1.046534774e-10 luc=-2.021399574e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=9.292141765e+04 lvsat=-2.556085955e-1
+  a0=1.626529302e+00 la0=-3.254408731e-6
+  ags=1.127437120e-01 lags=1.093860960e-8
+  a1=0.0
+  a2=1.083666533e+00 la2=-2.276004104e-6
+  b0=-1.709446520e-07 lb0=1.623339844e-12
+  b1=5.452591595e-09 lb1=-4.138244049e-14 pb1=2.117582368e-34
+  keta=3.421368674e-02 lketa=-2.173038039e-7
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-6.921953293e-02 lpclm=1.686371502e-06 wpclm=-1.110223025e-22 ppclm=1.776356839e-27
+  pdiblc1=0.39
+  pdiblc2=1.909636661e-03 lpdiblc2=-1.266443309e-8
+  pdiblcb=-0.225
+  drout=0.56
+  pscbe1=800000000.0
+  pscbe2=8.860770435e-09 lpscbe2=2.402531188e-14 wpscbe2=-5.293955920e-29
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=-6.686266667e-11 lalpha0=1.338825943e-15
+  alpha1=-6.686266667e-11 lalpha1=1.338825943e-15
+  beta0=4.805292000e+01 lbeta0=-3.614830047e-4
* Gidl Induced Drain Leakage Model Parameters
+  agidl=1.354378090e-10 lagidl=-8.225743918e-16 wagidl=8.271806126e-31
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.443915098e-01 lkt1=1.229746438e-7
+  kt2=-6.522345350e-02 lkt2=1.337061237e-7
+  at=7.716025872e+04 lat=-1.235502988e-1
+  ute=5.623649524e-01 lute=-1.292207756e-05 pute=-1.421085472e-26
+  ua1=3.775543044e-09 lua1=-3.374650014e-14
+  ub1=-2.648919653e-18 lub1=2.843379192e-23 wub1=-1.232595164e-38
+  uc1=-9.445040192e-11 luc1=1.294748875e-15
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.173 pmos
* Model Flag Parameters
+  lmin=4.0e-06 lmax=8.0e-06 wmin=5.4e-07 wmax=5.5e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.036424065e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-2.719534781e-7
+  k1=4.604103273e-01 lk1=-5.535191579e-8
+  k2=3.111376993e-02 lk2=-4.835272375e-8
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-1.903188674e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-1.051285932e-7
+  nfactor={7.782034620e-01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=5.692502402e-6
+  eta0=0.08
+  etab=-0.07
+  u0=5.374816804e-03 lu0=2.117898927e-8
+  ua=-5.231013447e-10 lua=1.676518894e-16
+  ub=-7.890771535e-20 lub=3.589066086e-24
+  uc=-1.070071013e-10 luc=-1.329647545e-18
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=6.344101412e+04 lvsat=-1.907198821e-2
+  a0=1.169202877e+00 la0=4.149589883e-7
+  ags=4.476786908e-02 lags=5.563441444e-7
+  a1=0.0
+  a2=0.8
+  b0=1.333762438e-07 lb0=-8.183849488e-13 wb0=2.117582368e-28 pb0=-8.470329473e-34
+  b1=-1.241682582e-09 lb1=1.232920225e-14
+  keta=7.540400483e-03 lketa=-3.290158170e-9
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-4.109336388e-01 lpclm=4.428121465e-06 wpclm=-8.881784197e-22 ppclm=-3.552713679e-27
+  pdiblc1=0.39
+  pdiblc2=2.318653116e-04 lpdiblc2=7.971988815e-10
+  pdiblcb=-0.225
+  drout=0.56
+  pscbe1=800000000.0
+  pscbe2=1.463489899e-08 lpscbe2=-2.230352405e-14
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=2.005880000e-10 lalpha0=-8.070698298e-16
+  alpha1=2.005880000e-10 lalpha1=-8.070698298e-16
+  beta0=-2.415876000e+01 lbeta0=2.179088540e-04 pbeta0=-3.410605132e-25
* Gidl Induced Drain Leakage Model Parameters
+  agidl=4.884466474e-11 lagidl=-1.277925667e-16 wagidl=-2.067951531e-31
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.137901907e-01 lkt1=-1.225556520e-7
+  kt2=-3.851363950e-02 lkt2=-8.060060310e-8
+  at=2.230282385e+04 lat=3.165994270e-1
+  ute=-1.918426857e+00 lute=6.982605139e-6
+  ua1=-2.965829131e-09 lua1=2.034303433e-14 wua1=3.308722450e-30 pua1=-3.970466940e-35
+  ub1=2.930570959e-18 lub1=-1.633336259e-23 wub1=6.162975822e-39
+  uc1=5.548297096e-10 luc1=-3.914763086e-15 puc1=-3.308722450e-36
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.174 pmos
* Model Flag Parameters
+  lmin=2.0e-06 lmax=4.0e-06 wmin=5.4e-07 wmax=5.5e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.106065230e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=8.249143277e-9
+  k1=3.853412315e-01 lk1=2.466900923e-7
+  k2=4.064949326e-02 lk2=-8.671989728e-8
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=8.635279899e-01 ldsub=-1.221250938e-6
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.223718520e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=2.383723148e-8
+  nfactor={2.270962668e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-3.136441188e-7
+  eta0=1.604349200e-01 leta0=-3.236315093e-7
+  etab=-1.403173200e-01 letab=2.829231434e-7
+  u0=1.211265930e-02 lu0=-5.930854756e-9
+  ua=-1.308633256e-10 lua=-1.410525625e-15
+  ub=6.187485939e-19 lub=7.820319721e-25
+  uc=-1.338088641e-10 luc=1.065077811e-16
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=8.388955365e+04 lvsat=-1.013470960e-1
+  a0=1.400765170e+00 la0=-5.167365282e-7
+  ags=-4.432097709e-02 lags=9.147948988e-7
+  a1=0.0
+  a2=0.8
+  b0=-1.003353178e-07 lb0=1.219581936e-13
+  b1=1.451284080e-09 lb1=1.493997030e-15
+  keta=2.281093733e-02 lketa=-6.473146857e-08 wketa=-5.551115123e-23
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=6.059902523e-01 lpclm=3.365078504e-7
+  pdiblc1=0.39
+  pdiblc2=4.185431636e-04 lpdiblc2=4.609681023e-11
+  pdiblcb=-4.273520000e-01 lpdiblcb=8.141673190e-7
+  drout=0.56
+  pscbe1=800000000.0
+  pscbe2=8.712478508e-09 lpscbe2=1.525453199e-15
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=-1.011760000e-10 lalpha0=4.070836595e-16
+  alpha1=-1.011760000e-10 lalpha1=4.070836595e-16
+  beta0=5.471942625e+01 lbeta0=-9.945910591e-05 pbeta0=4.547473509e-25
* Gidl Induced Drain Leakage Model Parameters
+  agidl=1.634728531e-11 lagidl=2.961289373e-18
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.355286288e-01 lkt1=-3.509061145e-8
+  kt2=-6.321122536e-02 lkt2=1.877062754e-8
+  at=1.626547485e+05 lat=-2.481093488e-1
+  ute=-9.154724880e-02 lute=-3.678815031e-7
+  ua1=2.886961000e-09 lua1=-3.205783819e-15
+  ub1=-1.904818744e-18 lub1=3.121924585e-24
+  uc1=-8.771411122e-10 luc1=1.846800155e-15
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.175 pmos
* Model Flag Parameters
+  lmin=1.0e-06 lmax=2.0e-06 wmin=5.4e-07 wmax=5.5e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.118108631e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=3.261920430e-8
+  k1=5.064652470e-01 lk1=1.593224533e-9
+  k2=-2.759691298e-03 lk2=1.119455858e-9
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=2.600000202e-01 ldsub=-2.071113059e-14
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.052413704e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-1.082664065e-8
+  nfactor={2.508128773e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-7.935544749e-07 wnfactor=1.421085472e-20
+  eta0=-5.005130400e-01 leta0=1.013809907e-06 weta0=7.355227538e-22 peta0=-4.163336342e-28
+  etab=2.645421120e-04 letab=-1.547066255e-9
+  u0=1.145910416e-02 lu0=-4.608372862e-9
+  ua=-3.318390994e-10 lua=-1.003847127e-15
+  ub=7.130469709e-19 lub=5.912173203e-25
+  uc=-1.196469642e-10 luc=7.785089353e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=1.537394825e+04 lvsat=3.729560184e-2
+  a0=1.030938530e+00 la0=2.316150734e-7
+  ags=2.475687006e-01 lags=3.241502982e-7
+  a1=0.0
+  a2=0.8
+  b0=2.062768896e-08 lb0=-1.228128700e-13
+  b1=-2.754611245e-08 lb1=6.017080885e-14 wb1=5.293955920e-29 pb1=2.646977960e-35
+  keta=-1.751182380e-02 lketa=1.686244502e-8
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=9.199174115e-01 lpclm=-2.987300348e-7
+  pdiblc1=3.957940034e-01 lpdiblc1=-1.172428182e-8
+  pdiblc2=4.529136727e-04 lpdiblc2=-2.345260230e-11
+  pdiblcb=1.797040000e-01 lpdiblcb=-4.142226381e-07 wpdiblcb=-2.220446049e-22 ppdiblcb=-6.661338148e-28
+  drout=3.794864141e-01 ldrout=3.652728512e-7
+  pscbe1=800000000.0
+  pscbe2=9.769526283e-09 lpscbe2=-6.135041137e-16
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=4.643241089e+00 lbeta0=1.871056290e-6
* Gidl Induced Drain Leakage Model Parameters
+  agidl=2.528734937e-11 lagidl=-1.512910906e-17
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.260591597e-01 lkt1=-5.425227153e-8
+  kt2=-5.943725826e-02 lkt2=1.113392964e-8
+  at=2.804660864e+04 lat=2.427291432e-2
+  ute=5.196833265e-01 lute=-1.604718797e-06 pute=-1.776356839e-27
+  ua1=3.076566596e-09 lua1=-3.589454534e-15
+  ub1=-1.607506698e-18 lub1=2.520307714e-24 pub1=6.162975822e-45
+  uc1=3.394859767e-12 luc1=6.501800488e-17
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=2.75e-6
+  sbref=2.74e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.176 pmos
* Model Flag Parameters
+  lmin=5.0e-07 lmax=1.0e-06 wmin=5.4e-07 wmax=5.5e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.104135008e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=1.831692178e-8
+  k1=5.845342661e-01 lk1=-7.831197791e-8
+  k2=-3.521780815e-02 lk2=3.434098762e-08 wk2=1.387778781e-23 pk2=3.469446952e-29
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=-5.148096000e-01 ldsub=7.930331218e-07 pdsub=-8.881784197e-28
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.286451354e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=1.312758095e-8
+  nfactor={5.348218125e-01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.226164665e-6
+  eta0=9.944947238e-01 leta0=-5.163604397e-7
+  etab=-1.505565344e-03 letab=2.646741292e-10
+  u0=5.252885488e-03 lu0=1.743816071e-9
+  ua=-1.855248330e-09 lua=5.553926879e-16
+  ub=1.646936524e-18 lub=-3.646373153e-25
+  uc=-3.861426543e-11 luc=-5.087694348e-18
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=5.284690706e+03 lvsat=4.762215872e-2
+  a0=1.406885884e+00 la0=-1.531745618e-7
+  ags=-1.537163707e-01 lags=7.348735944e-7
+  a1=0.0
+  a2=1.122324950e+00 la2=-3.299060332e-7
+  b0=-2.034000355e-07 lb0=1.064839866e-13
+  b1=6.395362368e-08 lb1=-3.348100107e-14
+  keta=4.345618449e-02 lketa=-4.553953082e-08 wketa=-9.714451465e-23 pketa=-2.775557562e-29
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=8.327961674e-01 lpclm=-2.095596990e-7
+  pdiblc1=7.135984939e-01 lpdiblc1=-3.370035339e-7
+  pdiblc2=3.879409928e-05 lpdiblc2=4.004070635e-10
+  pdiblcb=-0.225
+  drout=9.713112154e-01 ldrout=-2.404716693e-7
+  pscbe1=1.492842356e+09 lpscbe1=-7.091380085e+2
+  pscbe2=-6.308059837e-08 lpscbe2=7.395005547e-14 wpscbe2=-1.058791184e-28 ppscbe2=-1.058791184e-34
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=4.407774865e+00 lbeta0=2.112060679e-6
* Gidl Induced Drain Leakage Model Parameters
+  agidl=2.547348960e-12 lagidl=8.145736160e-18
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.740229702e-01 lkt1=-5.160352257e-9
+  kt2=-3.705763611e-02 lkt2=-1.177206122e-8
+  at=2.219515839e+04 lat=3.026199068e-2
+  ute=-1.895801293e+00 lute=8.675780209e-7
+  ua1=-2.625004008e-09 lua1=2.246217010e-15
+  ub1=2.657182254e-18 lub1=-1.844686722e-24 pub1=3.081487911e-45
+  uc1=2.075025205e-10 luc1=-1.438902680e-16 wuc1=8.271806126e-31 puc1=4.135903063e-37
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.75e-6
+  sbref=1.74e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.177 pmos
* Model Flag Parameters
+  lmin=2.5e-07 lmax=5.0e-07 wmin=5.4e-07 wmax=5.5e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.083600825e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=7.566866302e-9
+  k1=2.785842657e-01 lk1=8.185896632e-8
+  k2=9.078834505e-02 lk2=-3.162575371e-08 wk2=2.220446049e-22 pk2=5.551115123e-29
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=1.235674842e+00 ldsub=-1.233804932e-7
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={8.554790169e-02+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-1.513587578e-7
+  nfactor={3.380644558e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-2.636804585e-7
+  eta0=-5.189894481e-01 leta0=2.759787940e-07 weta0=-3.885780586e-22
+  etab=-2.015517863e-03 letab=5.316444720e-10
+  u0=1.182344359e-02 lu0=-1.696002504e-9
+  ua=-2.127182843e-10 lua=-3.045046414e-16
+  ub=5.497105694e-19 lub=2.097824166e-25
+  uc=-1.001292182e-10 luc=2.711661375e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=3.158190353e+04 lvsat=3.385504186e-2
+  a0=1.660440134e+00 la0=-2.859152828e-7
+  ags=9.698322770e-01 lags=1.466734064e-7
+  a1=0.0
+  a2=1.597024138e-01 la2=1.740461171e-7
+  b0=0.0
+  b1=0.0
+  keta=-5.647214109e-02 lketa=6.774946183e-9
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=2.085539131e-01 lpclm=1.172436059e-7
+  pdiblc1=-2.963791728e-01 lpdiblc1=1.917399742e-07 ppdiblc1=-2.220446049e-28
+  pdiblc2=-7.700523841e-03 lpdiblc2=4.452094792e-09 wpdiblc2=-6.938893904e-24 ppdiblc2=-5.204170428e-30
+  pdiblcb=-1.560512404e-01 lpdiblcb=-3.609605461e-8
+  drout=4.936971948e-01 ldrout=9.568822735e-9
+  pscbe1=-5.856554958e+08 lpscbe1=3.789971870e+02 ppscbe1=-9.536743164e-19
+  pscbe2=1.540275727e-07 lpscbe2=-3.971041422e-14
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=7.930281860e+00 lbeta0=2.679578173e-7
* Gidl Induced Drain Leakage Model Parameters
+  agidl=3.791729715e-11 lagidl=-1.037113912e-17
+  bgidl=7.372237654e+08 lbgidl=1.375686143e+2
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.00074326333
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.5407449e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.413228120e-01 lkt1=-2.227953908e-8
+  kt2=-6.690804875e-02 lkt2=3.855226801e-9
+  at=9.325182934e+04 lat=-6.937597694e-3
+  ute=4.134590933e-01 lute=-3.413659765e-07 pute=-4.440892099e-28
+  ua1=3.165106439e-09 lua1=-7.850216110e-16 pua1=3.308722450e-36
+  ub1=-1.629143462e-18 lub1=3.992905164e-25
+  uc1=-3.393906100e-11 luc1=-1.749077126e-17
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.1e-6
+  sbref=1.1e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.178 pmos
* Model Flag Parameters
+  lmin=1.8e-07 lmax=2.5e-07 wmin=5.4e-07 wmax=5.5e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.012266656e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-1.194445551e-8
+  k1=-8.579247482e-01 lk1=3.927169118e-7
+  k2=5.167953973e-01 lk2=-1.481472026e-7
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=1.803960266e+00 ldsub=-2.788179225e-7
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-7.309221625e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=7.196213411e-8
+  nfactor={2.983359543e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.550150614e-7
+  eta0=4.900000008e-01 leta0=-7.095835031e-17
+  etab=2.195759126e-03 letab=-6.202240101e-10 wetab=-3.469446952e-24 petab=-8.673617380e-31
+  u0=1.425126466e-02 lu0=-2.360060124e-9
+  ua=1.721124685e-09 lua=-8.334493704e-16
+  ub=-8.156452782e-19 lub=5.832345480e-25
+  uc=3.489543344e-11 luc=-9.815328983e-18 wuc=1.033975766e-31 puc=3.231174268e-39
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=3.617753405e+05 lvsat=-5.645946701e-2
+  a0=-1.466462483e-01 la0=2.083589844e-7
+  ags=2.250598986e+00 lags=-2.036419039e-7
+  a1=0.0
+  a2=9.336249622e-01 la2=-3.763717830e-8
+  b0=0.0
+  b1=0.0
+  keta=-8.737025015e-02 lketa=1.522619697e-8
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=6.849679741e-01 lpclm=-1.306516802e-8
+  pdiblc1=5.487137542e-01 lpdiblc1=-3.940984321e-8
+  pdiblc2=2.991525761e-02 lpdiblc2=-5.836573751e-9
+  pdiblcb=2.186325871e+00 lpdiblcb=-6.767830420e-7
+  drout=-8.416446543e-01 ldrout=3.748115253e-7
+  pscbe1=7.998956542e+08 lpscbe1=2.123647450e-2
+  pscbe2=1.957358274e-08 lpscbe2=-2.934558902e-15
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=1.052647787e+01 lbeta0=-4.421537155e-7
* Gidl Induced Drain Leakage Model Parameters
+  agidl=9.578483481e-15 lagidl=-2.619906802e-21
+  bgidl=1.938486425e+09 lbgidl=-1.910007484e+2
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.00074326333
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.5407449e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=2.438598179e-01 lkt1=-2.096906920e-7
+  kt2=-5.870698811e-02 lkt2=1.612072696e-9
+  at=2.121185134e+05 lat=-3.945001311e-2
+  ute=-1.856079955e+00 lute=2.793983441e-7
+  ua1=1.352904843e-10 lua1=4.369364895e-17
+  ub1=-3.305422621e-19 lub1=4.409711620e-26
+  uc1=-2.972920545e-10 luc1=5.454153952e-17
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.1e-6
+  sbref=1.1e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.179 pmos
* Model Flag Parameters
+  lmin=1.5e-07 lmax=1.8e-07 wmin=5.4e-07 wmax=5.5e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-2.026e-8
+  vth0={-6.474804959e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-9.338481841e-08 wvth0=-2.239651290e-07 pvth0=4.938879025e-14
+  k1=-3.250646473e-01 lk1=3.080141966e-07 wk1=8.145174527e-07 pk1=-1.796173887e-13
+  k2=-4.644389098e+00 lk2=9.776224850e-07 wk2=2.372551486e-06 pk2=-5.231950536e-13
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=5.340755379e+00 ldsub=-1.082041607e-06 wdsub=-2.103771968e-06 pdsub=4.639237944e-13
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={2.086293325e+01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-4.683903874e-06 wvoff=-1.134180329e-05 pvoff=2.501094461e-12
+  nfactor={3.464133704e+02+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-7.590114944e-05 wnfactor=-1.824989226e-04 pnfactor=4.024466241e-11
+  eta0=8.400759025e+00 leta0=-1.744480580e-06 weta0=-3.174366156e-06 peta0=7.000112247e-13
+  etab=4.527875495e-01 letab=-1.000365329e-07 wetab=-1.826105125e-07 petab=4.026927022e-14
+  u0=-5.075344287e-02 lu0=1.177764246e-08 wu0=2.651222386e-08 pu0=-5.846475606e-15
+  ua=-1.410045817e-09 lua=-2.125815723e-16 wua=-1.134355673e-15 pua=2.501481130e-22
+  ub=4.322556075e-19 lub=3.567649531e-25 wub=1.066697816e-24 pub=-2.352282025e-31
+  uc=-4.741072290e-10 luc=1.016100649e-16 wuc=1.997496677e-16 puc=-4.404879671e-23
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=2.641562598e+07 lvsat=-5.806570662e+00 wvsat=-1.402116566e+01 pvsat=3.091947450e-6
+  a0=-1.481837813e-01 la0=2.261022409e-07 wa0=8.563047240e-08 pa0=-1.888323177e-14
+  ags=1.249999924e+00 lags=1.854238008e-14 wags=7.358374887e-14 pags=-1.622668577e-20
+  a1=0.0
+  a2=-6.896131828e+00 la2=1.685836960e-06 wa2=3.359617793e-06 pa2=-7.408629158e-13
+  b0=0.0
+  b1=0.0
+  keta=-1.495159598e+00 lketa=3.269437463e-07 wketa=6.068561700e-07 pketa=-1.338239226e-13
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=6.657885017e-01 lpclm=-9.927042615e-09 wpclm=-2.774595610e-08 ppclm=6.118538239e-15
+  pdiblc1=1.346265424e+00 lpdiblc1=-2.185778367e-07 wpdiblc1=9.110364911e-08 ppdiblc1=-2.009017670e-14
+  pdiblc2=2.677645271e-02 lpdiblc2=-5.631932766e-09 wpdiblc2=-1.653930521e-08 ppdiblc2=3.647247585e-15
+  pdiblcb=-1.635021505e+01 lpdiblcb=3.354363360e-06 wpdiblcb=4.491185563e-06 ppdiblcb=-9.903962403e-13
+  drout=1.000000049e+00 ldrout=-5.076614684e-15 wdrout=7.514165645e-14 pdrout=-1.657023319e-20
+  pscbe1=1.299415028e+09 lpscbe1=-1.101310020e+02 wpscbe1=-2.004001866e+02 ppscbe1=4.419224916e-5
+  pscbe2=-1.480246716e-08 lpscbe2=4.400924285e-15 wpscbe2=-2.993349406e-15 ppscbe2=6.600934111e-22
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=1.828631003e+01 lbeta0=-2.190284947e-06 wbeta0=-4.056941559e-06 pbeta0=8.946367526e-13
* Gidl Induced Drain Leakage Model Parameters
+  agidl=-2.421667034e-14 lagidl=4.613760032e-21
+  bgidl=1.000000417e+09 lbgidl=-8.236108398e-05 wbgidl=-5.121087646e-05 pbgidl=1.129302216e-11
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-1.106e-8
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=3.511144361e+01 lkt1=-7.916205708e-06 wkt1=-1.943158332e-05 pkt1=4.285052753e-12
+  kt2=1.088471149e+00 lkt2=-2.512289938e-07 wkt2=-4.622717166e-07 pkt2=1.019401589e-13
+  at=-5.844186240e+05 lat=1.329071018e-01 wat=1.937588465e-01 pat=-4.272770084e-8
+  ute=-2.515781046e+00 lute=4.482137372e-07 wute=-6.669249331e-14 pute=1.470703026e-20
+  ua1=-1.852592475e-10 lua1=1.180310008e-16 wua1=-1.043621023e-15 pua1=2.301393080e-22
+  ub1=3.625483948e-18 lub1=-8.246023570e-25 wub1=-1.865208737e-25 pub1=4.113158307e-32
+  uc1=-7.639541558e-10 luc1=1.620057140e-16 wuc1=4.311016057e-16 puc1=-9.506652608e-23
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.04e-6
+  sbref=1.04e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.180 pmos
* Model Flag Parameters
+  lmin=2.0e-05 lmax=0.0001 wmin=4.2e-07 wmax=5.4e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.126311+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+  k1=0.43165561
+  k2=0.026980026
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=3.2465718e-7
+  voff={-0.23051772+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.8768912+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+  eta0=0.08
+  etab=-0.07
+  u0=0.0095864
+  ua=-7.4757916e-10
+  ub=9.5046395e-19
+  uc=-1.0566299e-10
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=80156.0
+  a0=1.464
+  ags=0.11329
+  a1=0.0
+  a2=0.97
+  b0=-8.9873e-8
+  b1=3.3859e-9
+  keta=0.023361259
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=0.015
+  pdiblc1=0.39
+  pdiblc2=0.0012771588
+  pdiblcb=-0.225
+  drout=0.56
+  pscbe1=800000000.0
+  pscbe2=1.0060625e-8
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=0.0
+  alpha1=0.0
+  beta0=30.0
* Gidl Induced Drain Leakage Model Parameters
+  agidl=9.43573999999999e-11
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-0.43825
+  kt2=-0.058546
+  at=70990.0
+  ute=-0.08298
+  ua1=2.0902e-9
+  ub1=-1.2289e-18
+  uc1=-2.9789e-11
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.181 pmos
* Model Flag Parameters
+  lmin=8.0e-06 lmax=2.0e-05 wmin=4.2e-07 wmax=5.4e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.219037832e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=1.856717570e-06 wvth0=2.882051378e-08 pvth0=-5.770881340e-13
+  k1=3.678002281e-01 lk1=1.278609517e-06 wk1=2.566840848e-08 pk1=-5.139718907e-13
+  k2=4.347795566e-02 lk2=-3.303466245e-07 wk2=-7.940258768e-09 pk2=1.589919303e-13
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=-6.144535039e-06 lcit=1.295359998e-10 wcit=-7.411538288e-28 pcit=4.235164736e-33
+  voff={-2.256707971e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-9.705245752e-08 wvoff=-1.197061096e-08 pvoff=2.396937679e-13
+  nfactor={4.813889219e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-5.880903857e-05 wnfactor=-1.395320716e-06 pnfactor=2.793923226e-11
+  eta0=0.08
+  etab=-0.07
+  u0=1.154013795e-02 lu0=-3.912071101e-08 wu0=-4.705401897e-10 pu0=9.421870900e-15
+  ua=-1.049188830e-09 lua=6.039287251e-15 wua=7.169930877e-17 pua=-1.435672543e-21
+  ub=1.521699024e-18 lub=-1.143813693e-23 wub=-9.490203445e-26 pub=1.900272785e-30
+  uc=-1.107681726e-10 luc=1.022237264e-16 wuc=3.187419409e-18 puc=-6.382335628e-23
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=1.356081232e+05 lvsat=-1.110346698e+00 wvsat=-2.225138439e-02 pvsat=4.455510404e-7
+  a0=2.018426298e+00 la0=-1.110156606e-05 wa0=-2.042849307e-07 pa0=4.090503396e-12
+  ags=1.385966975e-01 lags=-5.067291629e-07 wags=-1.347643746e-08 pags=2.698457151e-13
+  a1=0.0
+  a2=1.463759843e+00 la2=-9.886810092e-06 wa2=-1.981319997e-07 pa2=3.967300059e-12
+  b0=-2.850240693e-07 lb0=3.907611338e-12 wb0=5.946640601e-14 pb0=-1.190726770e-18
+  b1=6.534851399e-09 lb1=-6.305309131e-14 wb1=-5.641517322e-16 pb1=1.129630349e-20
+  keta=7.278892008e-02 lketa=-9.897157602e-07 wketa=-2.010818903e-08 pketa=4.026367253e-13
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-3.454727724e-01 lpclm=7.217933768e-06 wpclm=1.440030787e-07 ppclm=-2.883448525e-12
+  pdiblc1=0.39
+  pdiblc2=8.070424772e-03 lpdiblc2=-1.360250970e-07 wpdiblc2=-3.211446340e-09 ppdiblc2=6.430446002e-14
+  pdiblcb=-0.225
+  drout=0.56
+  pscbe1=4.870921626e+08 lpscbe1=6.265516340e+03 wpscbe1=1.631100942e+02 ppscbe1=-3.266038234e-3
+  pscbe2=4.060809250e-09 lpscbe2=1.201374307e-13 wpscbe2=2.502085367e-15 ppscbe2=-5.010055639e-20
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=-2.904469665e-10 lalpha0=5.815770642e-15 walpha0=1.165482351e-16 palpha0=-2.333705917e-21
+  alpha1=-2.904469665e-10 lalpha1=5.815770642e-15 walpha1=1.165482351e-16 palpha1=-2.333705917e-21
+  beta0=1.084206810e+02 lbeta0=-1.570258073e-03 wbeta0=-3.146802349e-05 pbeta0=6.301005977e-10
* Gidl Induced Drain Leakage Model Parameters
+  agidl=1.355639553e-10 lagidl=-8.251002840e-16 wagidl=-6.575651426e-20 pagidl=1.316676879e-24
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-6.164961059e-01 lkt1=3.569114466e-06 wkt1=8.971330702e-08 pkt1=-1.796376197e-12
+  kt2=-7.343082846e-02 lkt2=2.980466603e-07 wkt2=4.278274760e-09 pkt2=-8.566612021e-14
+  at=-3.857087195e+04 lat=2.193794311e+00 wat=6.032739794e-02 pat=-1.207966859e-6
+  ute=5.897759404e-01 lute=-1.347094203e-05 wute=-1.428858053e-08 pute=2.861076780e-13
+  ua1=5.823763019e-09 lua1=-7.475907378e-14 wua1=-1.067679723e-15 pua1=2.137870628e-20
+  ub1=-5.258272633e-18 lub1=8.068222350e-23 wub1=1.360182647e-24 pub1=-2.723564443e-29
+  uc1=-1.274889665e-10 luc1=1.956297233e-15 wuc1=1.722207863e-17 puc1=-3.448466359e-22
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.182 pmos
* Model Flag Parameters
+  lmin=4.0e-06 lmax=8.0e-06 wmin=4.2e-07 wmax=5.4e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-9.385022375e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-3.941653806e-07 wvth0=-5.104390693e-08 pvth0=6.370564283e-14
+  k1=5.245517312e-01 lk1=2.091069709e-08 wk1=-3.343511789e-08 pk1=-3.975356474e-14
+  k2=1.825892600e-02 lk2=-1.280012357e-07 wk2=6.700870205e-09 pk2=4.151853911e-14
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.939243404e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=4.505812123e-07 wvoff=5.400663215e-08 pvoff=-2.896759617e-13
+  nfactor={-8.135979557e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=4.509449255e-05 wnfactor=4.646714010e-06 pnfactor=-2.053915421e-11
+  eta0=0.08
+  etab=-0.07
+  u0=2.602979050e-03 lu0=3.258676221e-08 wu0=1.444881410e-09 pu0=-5.946552613e-15
+  ua=-4.660448638e-10 lua=1.360419979e-15 wua=-2.974194591e-17 pua=-6.217566074e-22
+  ub=-4.727047021e-19 lub=4.564001255e-24 wub=2.052753429e-25 pub=-5.082064058e-31
+  uc=-8.792147730e-11 luc=-8.108719050e-17 wuc=-9.948801378e-18 puc=4.157537393e-23
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=-7.769950388e+04 lvsat=6.011313138e-01 wvsat=7.357260010e-02 pvsat=-3.232946157e-7
+  a0=-4.988320312e-02 la0=5.493556585e-06 wa0=6.354754391e-07 pa0=-2.647330726e-12
+  ags=1.001309988e-03 lags=5.972701805e-07 wags=2.281428179e-08 pags=-2.133359666e-14
+  a1=0.0
+  a2=-3.402799291e-01 la2=4.587939100e-06 wa2=5.943959992e-07 pa2=-2.391564191e-12
+  b0=5.364888499e-07 lb0=-2.683813999e-12 wb0=-2.101313144e-13 pb0=9.723959319e-19
+  b1=-4.270837353e-09 lb1=2.364656850e-14 wb1=1.579013566e-15 pb1=-5.899426137e-21
+  keta=-8.490294513e-02 lketa=2.755280741e-07 wketa=4.818812765e-08 pketa=-1.453401376e-13
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-7.479194529e-01 lpclm=1.044697276e-05 wpclm=1.756612693e-07 ppclm=-3.137458651e-12
+  pdiblc1=0.39
+  pdiblc2=-1.775084640e-02 lpdiblc2=7.115238866e-08 wpdiblc2=9.373884102e-09 ppdiblc2=-3.667419049e-14
+  pdiblcb=-0.225
+  drout=0.56
+  pscbe1=1.738723512e+09 lpscbe1=-3.776972826e+03 wpscbe1=-4.893302827e+02 ppscbe1=1.968830179e-3
+  pscbe2=3.058199753e-08 lpscbe2=-9.265585393e-14 wpscbe2=-8.312775951e-15 ppscbe2=3.667269970e-20
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=8.713408995e-10 lalpha0=-3.505857536e-15 walpha0=-3.496447054e-16 palpha0=1.406802465e-21
+  alpha1=8.713408995e-10 lalpha1=-3.505857536e-15 walpha1=-3.496447054e-16 palpha1=1.406802465e-21
+  beta0=-2.052620429e+02 lbeta0=9.465815347e-04 wbeta0=9.440407046e-05 pbeta0=-3.798366656e-10
* Gidl Induced Drain Leakage Model Parameters
+  agidl=6.219379984e-11 lagidl=-2.364133743e-16 wagidl=-6.958530351e-18 pagidl=5.662098562e-23
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=1.899770848e-01 lkt1=-2.901639309e-06 wkt1=-3.147269752e-07 pkt1=1.448658496e-12
+  kt2=-1.389151463e-02 lkt2=-1.796682150e-07 wkt2=-1.283482428e-08 pkt2=5.164117218e-14
+  at=2.685883460e+05 lat=-2.707038177e-01 wat=-1.283817467e-01 pat=3.061447370e-7
+  ute=-1.798844082e+00 lute=5.694198491e-06 wute=-6.233515266e-08 pute=6.716103105e-13
+  ua1=-9.110489056e-09 lua1=4.506619643e-14 wua1=3.203039168e-15 pua1=-1.288749215e-20
+  ub1=1.075862990e-17 lub1=-4.782971430e-23 wub1=-4.080547940e-24 pub1=1.641816625e-29
+  uc1=1.960201142e-09 luc1=-1.479432611e-14 wuc1=-7.325807773e-16 puc1=5.671211575e-21
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.183 pmos
* Model Flag Parameters
+  lmin=2.0e-06 lmax=4.0e-06 wmin=4.2e-07 wmax=5.4e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-8.674727712e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-6.799538588e-07 wvth0=-1.243715684e-07 pvth0=3.587409553e-13
+  k1=4.326883529e-01 lk1=3.905248369e-07 wk1=-2.468072863e-08 pk1=-7.497702499e-14
+  k2=6.987632793e-02 lk2=-3.356848847e-07 wk2=-1.523513056e-08 pk2=1.297784769e-13
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=8.635279560e-01 ldsub=-1.221250802e-06 wdsub=1.763597646e-14 pdsub=-7.095870469e-20
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-1.799276959e-02+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-6.596349816e-07 wvoff=-1.065370930e-07 pvoff=3.562749274e-13
+  nfactor={6.734994912e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.473917064e-05 wnfactor=-2.326975016e-06 pnfactor=7.519623062e-12
+  eta0=1.604349200e-01 leta0=-3.236315093e-7
+  etab=-1.403173200e-01 letab=2.829231434e-7
+  u0=2.028548977e-03 lu0=3.489799309e-08 wu0=5.256564355e-09 pu0=-2.128293518e-14
+  ua=-2.130938621e-10 lua=3.426665642e-16 wua=4.286447621e-17 pua=-9.138899990e-22
+  ub=-6.852004360e-19 lub=5.418982091e-24 wub=6.797121187e-25 pub=-2.417112262e-30
+  uc=-9.429779189e-11 luc=-5.543196120e-17 wuc=-2.059601561e-17 puc=8.441465332e-23
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=1.672335230e+05 lvsat=-3.843616184e-01 wvsat=-4.344487758e-02 pvsat=1.475275461e-7
+  a0=1.772657770e+00 la0=-1.839473471e-06 wa0=-1.938571996e-07 pa0=6.895057318e-13
+  ags=-5.448374449e-01 lags=2.793463328e-06 wags=2.609052202e-07 pags=-9.792972492e-13
+  a1=0.0
+  a2=0.8
+  b0=3.750320935e-08 lb0=-6.761352945e-13 wb0=-7.185136475e-14 pb0=4.160237887e-19
+  b1=2.648032470e-07 lb1=-1.058978391e-12 wb1=-1.372780044e-13 pb1=5.527945629e-19
+  keta=3.671945602e-03 lketa=-8.085477023e-08 wketa=9.976620494e-09 pketa=8.404625702e-15
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=2.472467495e+00 lpclm=-2.510318534e-06 wpclm=-9.729423251e-07 ppclm=1.483970883e-12
+  pdiblc1=0.39
+  pdiblc2=-6.190729664e-04 lpdiblc2=2.222355596e-09 wpdiblc2=5.408802353e-10 ppdiblc2=-1.134422770e-15
+  pdiblcb=-1.104003598e+00 lpdiblcb=3.536688556e-06 wpdiblcb=3.527195317e-07 ppdiblcb=-1.419174090e-12
+  drout=0.56
+  pscbe1=800000000.0
+  pscbe2=5.319651270e-09 lpscbe2=8.987701501e-15 wpscbe2=1.768585840e-15 ppscbe2=-3.889861097e-21
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=-1.011760000e-10 lalpha0=4.070836595e-16
+  alpha1=-1.011760000e-10 lalpha1=4.070836595e-16
+  beta0=5.150479931e+01 lbeta0=-8.652499013e-05 wbeta0=1.675695013e-06 pbeta0=-6.742192400e-12
* Gidl Induced Drain Leakage Model Parameters
+  agidl=-3.023044261e-11 lagidl=1.354574137e-16 wagidl=2.427966539e-17 pagidl=-6.906651970e-23
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-8.918211702e-01 lkt1=1.450997606e-06 wkt1=2.378525256e-07 pkt1=-7.746561772e-13
+  kt2=-5.744277049e-02 lkt2=-4.438866005e-09 wkt2=-3.006934008e-09 pkt2=1.209845912e-14
+  at=2.628306516e+05 lat=-2.475376193e-01 wat=-5.221889339e-02 pat=-2.980265590e-10
+  ute=-3.176579848e+00 lute=1.123754590e-05 wute=1.608141113e-06 pute=-6.049584353e-12
+  ua1=2.127381787e-11 lua1=8.324365872e-15 wua1=1.493802489e-15 pua1=-6.010344190e-21
+  ub1=-1.600900679e-18 lub1=1.899104171e-24 wub1=-1.584239777e-25 pub1=6.374220426e-31
+  uc1=-3.433436375e-09 luc1=6.907082315e-15 wuc1=1.332525144e-15 puc1=-2.637783402e-21
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.184 pmos
* Model Flag Parameters
+  lmin=1.0e-06 lmax=2.0e-06 wmin=4.2e-07 wmax=5.4e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.413802750e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=4.255557794e-07 wvth0=1.541370649e-07 pvth0=-2.048268344e-13
+  k1=6.526904988e-01 lk1=-5.465390546e-08 wk1=-7.622312947e-08 pk1=2.932005394e-14
+  k2=-1.554261101e-01 lk2=1.202191047e-07 wk2=7.958072946e-08 pk2=-6.208331216e-14
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=2.792711245e+00 ldsub=-5.124991771e-06 wdsub=-1.320231446e-06 pdsub=2.671514700e-12
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-4.435697243e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=2.015284978e-07 wvoff=1.242338977e-07 pvoff=-1.106947877e-13
+  nfactor={4.981906464e-01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-2.118872476e-06 wnfactor=1.047724467e-06 pnfactor=6.908511650e-13
+  eta0=-1.424610354e+00 leta0=2.883739304e-06 weta0=4.817060552e-07 peta0=-9.747418368e-13
+  etab=-2.892223598e+00 letab=5.851460534e-06 wetab=1.507773078e-06 petab=-3.051008978e-12
+  u0=3.443501426e-02 lu0=-3.067713754e-08 wu0=-1.197669861e-08 pu0=1.358891710e-14
+  ua=1.503569224e-09 lua=-3.131035524e-15 wua=-9.567469677e-16 pua=1.108843750e-21
+  ub=2.581860102e-18 lub=-1.191980250e-24 wub=-9.741599586e-25 pub=9.295309638e-31
+  uc=-2.372030897e-10 luc=2.337397670e-16 wuc=6.127871664e-17 puc=-8.126050486e-23
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=-1.385557808e+05 lvsat=2.344091535e-01 wvsat=8.023925771e-02 pvsat=-1.027497753e-7
+  a0=2.390537165e-02 la0=1.699161982e-06 wa0=5.249381886e-07 pa0=-7.649911121e-13
+  ags=1.931257553e+00 lags=-2.216964424e-06 wags=-8.776598557e-07 pags=1.324611953e-12
+  a1=0.0
+  a2=0.8
+  b0=-3.788214190e-07 lb0=1.663059175e-13 wb0=2.082216354e-13 pb0=-1.507095286e-19
+  b1=-6.546755941e-07 lb1=8.016054331e-13 wb1=3.269050392e-13 pb1=-3.864891095e-19
+  keta=-1.163336882e-01 lketa=1.619790299e-07 wketa=5.151307091e-08 pketa=-7.564521245e-14
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=1.076016123e+00 lpclm=3.154287453e-07 wpclm=-8.136988773e-08 ppclm=-3.201437757e-13
+  pdiblc1=4.105462587e-01 lpdiblc1=-4.157576546e-08 wpdiblc1=-7.689937624e-09 ppdiblc1=1.556074258e-14
+  pdiblc2=5.295354667e-04 lpdiblc2=-1.018765409e-10 wpdiblc2=-3.994079580e-11 ppdiblc2=4.088020332e-17
+  pdiblcb=1.533007196e+00 lpdiblcb=-1.799355525e-06 wpdiblcb=-7.054390634e-07 ppdiblcb=7.220309902e-13
+  drout=7.504845501e-01 ldrout=-3.854492968e-07 wdrout=-1.933909403e-07 pdrout=3.913304356e-13
+  pscbe1=800000000.0
+  pscbe2=1.011067100e-08 lpscbe2=-7.070227457e-16 wpscbe2=-1.778291899e-16 ppscbe2=4.874864434e-23
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=2.091751448e-11 lalpha0=1.600249911e-16 walpha0=4.122348539e-17 palpha0=-8.341654716e-23
+  alpha1=-5.845165291e-10 lalpha1=1.385132887e-15 walpha1=3.568193001e-16 palpha1=-7.220309902e-22
+  beta0=1.035183562e+01 lbeta0=-3.251145041e-06 wbeta0=-2.975730489e-06 pbeta0=2.670060132e-12
* Gidl Induced Drain Leakage Model Parameters
+  agidl=5.067934279e-11 lagidl=-2.826515530e-17 wagidl=-1.323613520e-17 pagidl=6.847453099e-24
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=1.915921971e-01 lkt1=-7.413110111e-07 wkt1=-3.219643581e-07 pkt1=3.581444833e-13
+  kt2=-8.064576707e-02 lkt2=4.251286165e-08 wkt2=1.105540181e-08 pkt2=-1.635695865e-14
+  at=1.902595921e+05 lat=-1.006886290e-01 wat=-8.455708632e-02 pat=6.513895359e-8
+  ute=6.014459668e+00 lute=-7.360706380e-06 wute=-2.864273053e-06 pute=3.000435159e-12
+  ua1=8.200411971e-09 lua1=-8.226283763e-15 wua1=-2.670917126e-15 pua1=2.417049246e-21
+  ub1=-1.175855023e-18 lub1=1.039015785e-24 wub1=-2.250079321e-25 pub1=7.721560061e-31
+  uc1=2.855442131e-11 luc1=-9.832530060e-17 wuc1=-1.311497497e-17 puc1=8.514629154e-23
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=2.75e-6
+  sbref=2.74e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.185 pmos
* Model Flag Parameters
+  lmin=5.0e-07 lmax=1.0e-06 wmin=4.2e-07 wmax=5.4e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-9.944840031e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-3.625344272e-09 wvth0=-5.715799847e-08 pvth0=1.143788891e-14
+  k1=9.996026328e-01 lk1=-4.097254129e-07 wk1=-2.163635177e-07 pk1=1.727565441e-13
+  k2=-1.935714746e-01 lk2=1.592616482e-07 wk2=8.254533240e-08 pk2=-6.511764256e-14
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=-8.171143564e+00 ldsub=6.096732903e-06 wdsub=3.991032518e-06 pdsub=-2.764670192e-12
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.867046334e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=4.097393993e-08 wvoff=3.026479061e-08 pvoff=-1.451552724e-14
+  nfactor={-4.877113666e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=3.382858994e-06 wnfactor=2.821090431e-06 pnfactor=-1.124224366e-12
+  eta0=4.529686076e+00 leta0=-3.210602178e-06 weta0=-1.842796266e-06 peta0=1.404432779e-12
+  etab=5.786950059e+00 letab=-3.031847287e-06 wetab=-3.017359840e-06 petab=1.580555066e-12
+  u0=-9.274202173e-03 lu0=1.406011966e-08 wu0=7.572564040e-09 pu0=-6.420144206e-15
+  ua=-5.113614796e-09 lua=3.641784664e-15 wua=1.698495204e-15 pua=-1.608849718e-21
+  ub=3.700142673e-18 lub=-2.336564827e-24 wub=-1.070278876e-24 pub=1.027910598e-30
+  uc=1.403305441e-10 luc=-1.526734579e-16 wuc=-9.327891877e-17 puc=7.693232613e-23
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=1.525874702e+05 lvsat=-6.358178675e-02 wvsat=-7.678481449e-02 pvsat=5.796750307e-8
+  a0=1.328196563e+00 la0=3.641938621e-07 wa0=4.101853973e-08 pa0=-2.696896731e-13
+  ags=-1.789367385e+00 lags=1.591169613e-06 wags=8.526190754e-07 pags=-4.463631384e-13
+  a1=0.0
+  a2=2.795367529e+00 la2=-2.042298573e-06 wa2=-8.721102509e-07 pa2=8.926222840e-13
+  b0=-4.428507626e-07 lb0=2.318412312e-13 wb0=1.248189594e-13 pb0=-6.534522162e-20
+  b1=2.630637381e-07 lb1=-1.377191282e-13 wb1=-1.037905276e-13 pb1=5.433641699e-20
+  keta=1.816767316e-01 lketa=-1.430405949e-07 wketa=-7.205050102e-08 pketa=5.082457469e-14
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=1.002631546e+00 lpclm=3.905393281e-07 wpclm=-8.853042744e-08 ppclm=-3.128148201e-13
+  pdiblc1=4.850946201e-01 lpdiblc1=-1.178775043e-07 wpdiblc1=1.191126713e-07 ppdiblc1=-1.142242637e-13
+  pdiblc2=-2.680806485e-03 lpdiblc2=3.183972654e-09 wpdiblc2=1.417651636e-09 ppdiblc2=-1.450994802e-15
+  pdiblcb=2.123247738e-01 lpdiblcb=-4.476106525e-07 wpdiblcb=-2.279651595e-07 ppdiblcb=2.333269001e-13
+  drout=1.938003494e+00 ldrout=-1.600898687e-06 wdrout=-5.039096177e-07 pdrout=7.091525122e-13
+  pscbe1=3.809661006e+09 lpscbe1=-3.080448233e+03 wpscbe1=-1.207692691e+03 ppscbe1=1.236097623e-3
+  pscbe2=-3.042480798e-07 lpscbe2=3.210454458e-13 wpscbe2=1.257138554e-13 ppscbe2=-1.288039083e-19
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=2.581649710e-10 lalpha0=-8.280252564e-17 walpha0=-8.244697079e-17 palpha0=4.316263815e-23
+  alpha1=1.469033058e-09 lalpha1=-7.167161866e-16 walpha1=-7.136386003e-16 palpha1=3.736040800e-22
+  beta0=4.882723422e+00 lbeta0=2.346600676e-06 wbeta0=-2.475773844e-07 pbeta0=-1.222591332e-13
* Gidl Induced Drain Leakage Model Parameters
+  agidl=-1.101406921e-11 lagidl=3.487928576e-17 wagidl=7.069187574e-18 pagidl=-1.393545086e-23
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-6.538080550e-01 lkt1=1.239730549e-07 wkt1=9.371693074e-08 pkt1=-6.731362943e-14
+  kt2=-1.771443798e-02 lkt2=-2.189861231e-08 wkt2=-1.008306758e-08 pkt2=5.278687539e-15
+  at=1.043285375e+05 lat=-1.273647596e-02 wat=-4.281383080e-02 pat=2.241389670e-8
+  ute=-1.914663261e+00 lute=7.549095197e-07 wute=9.832215555e-09 pute=5.873093498e-14
+  ua1=-2.613319453e-09 lua1=2.841786624e-15 wua1=-6.090831250e-18 pua1=-3.104537637e-22
+  ub1=8.177959453e-19 lub1=-1.001525854e-24 wub1=9.588205798e-25 pub1=-4.395161524e-31
+  uc1=-6.768146163e-11 luc1=1.740503130e-19 wuc1=1.434457047e-16 puc1=-7.509669533e-23
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.75e-6
+  sbref=1.74e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.186 pmos
* Model Flag Parameters
+  lmin=2.5e-07 lmax=5.0e-07 wmin=4.2e-07 wmax=5.4e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-9.210736770e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-4.205711818e-08 wvth0=-8.472085133e-08 pvth0=2.586759364e-14
+  k1=8.237492375e-01 lk1=-3.176626434e-07 wk1=-2.841792352e-07 pk1=2.082594285e-13
+  k2=-1.419146917e-01 lk2=1.322182892e-07 wk2=1.213015774e-07 pk2=-8.540731193e-14
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=5.969492188e+00 ldsub=-1.306172726e-06 wdsub=-2.467606436e-06 pdsub=6.165564728e-13
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={3.841641620e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-3.102392918e-07 wvoff=-1.556602952e-07 pvoff=8.281997371e-14
+  nfactor={1.263844159e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.679447531e-07 wnfactor=1.103428777e-06 pnfactor=-2.249941373e-13
+  eta0=-3.892982897e+00 leta0=1.198833483e-06 weta0=1.758768313e-06 peta0=-4.810583092e-13
+  etab=-8.734375648e-03 letab=2.309428144e-09 wetab=3.502352435e-09 petab=-9.267088500e-16
+  u0=1.784056003e-02 lu0=-1.350006461e-10 wu0=-3.136554324e-09 pu0=-8.137065605e-16
+  ua=4.670154407e-10 lua=7.202131224e-16 wua=-3.543261583e-16 pua=-5.341566782e-22
+  ub=7.523483469e-19 lub=-7.933355413e-25 wub=-1.056293996e-25 pub=5.228973041e-31
+  uc=-3.111822620e-10 luc=8.370252639e-17 wuc=1.100160422e-16 puc=-2.949665186e-23
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=-5.770045568e+04 lvsat=4.650814822e-02 wvsat=4.654039395e-02 pvsat=-6.595710057e-9
+  a0=5.581686763e+00 la0=-1.862593327e-06 wa0=-2.044036073e-06 pa0=8.218781176e-13
+  ags=3.297008897e-02 lags=6.371394990e-07 wags=4.883600265e-07 pags=-2.556662411e-13
+  a1=0.0
+  a2=-4.443183087e+00 la2=1.747227446e-06 wa2=2.399355331e-06 pa2=-8.200553774e-13
+  b0=0.0
+  b1=0.0
+  keta=-1.442854522e-01 lketa=2.760712753e-08 wketa=4.577462033e-08 pketa=-1.085923283e-14
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=3.657737216e+00 lpclm=-9.994615926e-07 wpclm=-1.797962679e-06 ppclm=5.821071522e-13
+  pdiblc1=-6.917757901e-01 lpdiblc1=4.982376929e-07 wpdiblc1=2.061091855e-07 ppdiblc1=-1.597686788e-13
+  pdiblc2=-9.147055194e-03 lpdiblc2=6.569183178e-09 wpdiblc2=7.540362915e-10 ppdiblc2=-1.103578897e-15
+  pdiblcb=-8.001407327e-01 lpdiblcb=8.243528945e-08 wpdiblcb=3.357458178e-07 ppdiblcb=-6.178707078e-14
+  drout=-1.206281109e+00 ldrout=4.519718866e-08 wdrout=8.861510902e-07 pdrout=-1.857206956e-14
+  pscbe1=-5.219310158e+09 lpscbe1=1.646398751e+03 wpscbe1=2.415394433e+03 ppscbe1=-6.606609478e-4
+  pscbe2=6.391147549e-07 lpscbe2=-1.728238654e-13 wpscbe2=-2.528623657e-13 ppscbe2=6.938831490e-20
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=1.050424620e+01 lbeta0=-5.963789270e-07 wbeta0=-1.341735538e-06 pbeta0=4.505545433e-13
* Gidl Induced Drain Leakage Model Parameters
+  agidl=1.164528010e-10 lagidl=-3.185217012e-17 wagidl=-4.093835914e-17 pagidl=1.119745999e-23
+  bgidl=-1.414824446e+08 lbgidl=5.975888894e+02 wbgidl=4.580449435e+02 pbgidl=-2.397956888e-4
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-6.153156046e-01 lkt1=1.038214873e-07 wkt1=9.069757102e-08 pkt1=-6.573293423e-14
+  kt2=-2.856596699e-02 lkt2=-1.621761984e-08 wkt2=-1.998665364e-08 pkt2=1.046341291e-14
+  at=2.291783275e+05 lat=-7.809783800e-02 wat=-7.085467753e-02 pat=3.709384078e-8
+  ute=1.421668901e+00 lute=-9.917270933e-07 wute=-5.255515426e-07 pute=3.390150401e-13
+  ua1=5.565611091e-09 lua1=-1.440047095e-15 wua1=-1.251315861e-15 pua1=3.414464438e-22
+  ub1=-1.289193713e-18 lub1=1.015253722e-25 wub1=-1.772062858e-25 pub1=1.552166323e-31
+  uc1=1.107595423e-10 luc1=-9.324338408e-17 wuc1=-7.542733036e-17 puc1=3.948771599e-23
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.1e-6
+  sbref=1.1e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.187 pmos
* Model Flag Parameters
+  lmin=1.8e-07 lmax=2.5e-07 wmin=4.2e-07 wmax=5.4e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-8.851391922e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-5.188591846e-08 wvth0=-6.626798731e-08 pvth0=2.082036627e-14
+  k1=-6.574608203e+00 lk1=1.705936084e-06 wk1=2.979947018e-06 pk1=-6.845443842e-13
+  k2=2.694294218e+00 lk2=-6.435415718e-07 wk2=-1.135069165e-06 pk2=2.582352136e-13
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=5.622145527e+00 ldsub=-1.211166467e-06 wdsub=-1.990313067e-06 pdsub=4.860071907e-13
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-1.892956359e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=3.125987131e-07 wvoff=6.057358897e-07 pvoff=-1.254371108e-13
+  nfactor={4.339742980e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-6.733750923e-07 wnfactor=-7.070447069e-07 pnfactor=2.702065700e-13
+  eta0=4.900000034e-01 leta0=-3.082458733e-16 weta0=-1.384213189e-15 peta0=1.236903913e-22
+  etab=9.559130842e-03 letab=-2.694211752e-09 wetab=-3.838319501e-09 petab=1.081111738e-15
+  u0=5.482850678e-02 lu0=-1.025194384e-08 wu0=-2.115178015e-08 pu0=4.113818008e-15
+  ua=1.633664700e-08 lua=-3.620448502e-15 wua=-7.618662548e-15 pua=1.452784611e-21
+  ub=-1.141081170e-17 lub=2.533531994e-24 wub=5.522963590e-24 pub=-1.016635450e-30
+  uc=1.507205646e-10 luc=-4.263713475e-17 wuc=-6.037639777e-17 puc=1.710908833e-23
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=1.009001464e+06 lvsat=-2.452561607e-01 wvsat=-3.373808556e-01 pvsat=9.841443013e-8
+  a0=-4.537101132e+00 la0=9.050975375e-07 wa0=2.288621198e-06 pa0=-3.631902991e-13
+  ags=5.596535288e+00 lags=-8.846068543e-07 wags=-1.744142908e-06 pags=3.549679616e-13
+  a1=0.0
+  a2=2.542488304e+00 la2=-1.634933934e-07 wa2=-8.386554118e-07 pa2=6.560532094e-14
+  b0=0.0
+  b1=0.0
+  keta=-2.851689600e-01 lketa=6.614158458e-08 wketa=1.031069291e-07 pketa=-2.654076593e-14
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=2.111615595e-01 lpclm=-5.675421888e-08 wpclm=2.469820173e-07 ppclm=2.277387892e-14
+  pdiblc1=1.755692126e+00 lpdiblc1=-1.711937316e-07 wpdiblc1=-6.291640299e-07 ppdiblc1=6.869525106e-14
+  pdiblc2=1.075642290e-01 lpdiblc2=-2.535368727e-08 wpdiblc2=-4.047623460e-08 ppdiblc2=1.017372480e-14
+  pdiblcb=1.024963883e+01 lpdiblcb=-2.939900416e-06 wpdiblcb=-4.203179271e-06 ppdiblcb=1.179699720e-12
+  drout=-6.993642508e+00 ldrout=1.628156279e-06 wdrout=3.206864225e-06 pdrout=-6.533335262e-13
+  pscbe1=7.996518954e+08 lpscbe1=9.224982947e-02 wpscbe1=1.270646314e-01 ppscbe1=-3.701727357e-8
+  pscbe2=5.386929887e-08 lpscbe2=-1.274752823e-14 wpscbe2=-1.787739654e-14 ppscbe2=5.115226149e-21
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=1.534596650e+01 lbeta0=-1.920686263e-06 wbeta0=-2.512264475e-06 pbeta0=7.707176182e-13
* Gidl Induced Drain Leakage Model Parameters
+  agidl=4.160829368e-14 lagidl=-1.138070049e-20 wagidl=-1.669624322e-20 pagidl=4.566756445e-27
+  bgidl=5.076722465e+09 lbgidl=-8.296945176e+02 wbgidl=-1.635874577e+03 pbgidl=3.329331785e-4
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=3.094482121e+00 lkt1=-9.108823866e-07 wkt1=-1.485949589e-06 pkt1=3.655115970e-13
+  kt2=-1.134605128e-01 lkt2=7.002736321e-09 wkt2=2.854147930e-08 pkt2=-2.810002009e-15
+  at=5.701785796e+05 lat=-1.713682270e-01 wat=-1.866466868e-01 pat=6.876527117e-8
+  ute=-6.641415603e+00 lute=1.213687780e-06 wute=2.494461484e-06 pute=-4.870189229e-13
+  ua1=-3.931831201e-10 lua1=1.898022981e-16 wua1=2.754784927e-16 pua1=-7.616234778e-23
+  ub1=-1.618345368e-18 lub1=1.915549330e-25 wub1=6.712957006e-25 pub1=-7.686563106e-32
+  uc1=-1.096348514e-09 luc1=2.369248116e-16 wuc1=4.165257589e-16 puc1=-9.507129300e-23
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.1e-6
+  sbref=1.1e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.188 pmos
* Model Flag Parameters
+  lmin=1.5e-07 lmax=1.8e-07 wmin=4.2e-07 wmax=5.4e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-2.026e-8
+  vth0={-1.664536521e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=1.156527562e-07 wvth0=3.061976993e-07 pvth0=-5.957664437e-14
+  k1=5.083907541e+00 lk1=-7.225031816e-07 wk1=-2.005028298e-06 pk1=3.575624661e-13
+  k2=-1.385193918e+00 lk2=2.023122055e-07 wk2=6.736242960e-07 pk2=-1.190475136e-13
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=-2.672875551e-01 ldsub=-1.359726677e-08 wdsub=8.195437880e-07 pdsub=-9.302632354e-14
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.465724221e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=4.650168132e-07 wvoff=8.187726520e-07 pvoff=-1.828937237e-13
+  nfactor={-2.305959014e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=5.312478911e-06 wnfactor=1.009698649e-05 pnfactor=-2.089728068e-12
+  eta0=8.400758521e+00 leta0=-1.744480469e-06 weta0=-3.174365893e-06 peta0=7.000111666e-13
+  etab=4.320056556e-01 letab=-9.607716656e-08 wetab=-1.717774931e-07 petab=3.820536343e-14
+  u0=2.493779623e-02 lu0=-4.516787929e-09 wu0=-1.294349973e-08 pu0=2.647354709e-15
+  ua=5.363893492e-09 lua=-1.503152506e-15 wua=-4.665420564e-15 pua=9.228866047e-22
+  ub=-7.009096801e-18 lub=1.774491434e-24 wub=4.945666469e-24 pub=-9.742493206e-31
+  uc=-8.081621033e-10 luc=1.652541967e-16 wuc=3.738831201e-16 puc=-7.722470056e-23
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=-3.864694136e+06 lvsat=8.090049766e-01 wvsat=1.763117371e+00 pvsat=-3.565668939e-7
+  a0=-7.256387058e+00 la0=1.580357153e-06 wa0=3.790937811e-06 pa0=-7.248183985e-13
+  ags=1.250000285e+00 lags=-5.467549702e-14 wags=-1.144278841e-13 pags=2.193974602e-20
+  a1=0.0
+  a2=3.844541110e-01 la2=2.987397243e-07 wa2=-4.355478003e-07 pa2=-1.780796534e-14
+  b0=0.0
+  b1=0.0
+  keta=-1.110167005e+00 lketa=2.535949516e-07 wketa=4.061703108e-07 pketa=-9.558924971e-14
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-4.394951055e+00 lpclm=9.542450621e-07 wpclm=2.610275874e-06 ppclm=-4.964773831e-13
+  pdiblc1=5.458634989e+00 lpdiblc1=-1.002066483e-06 wpdiblc1=-2.052559459e-06 ppdiblc1=3.883205167e-13
+  pdiblc2=-1.073643652e-01 lpdiblc2=1.992457601e-08 wpdiblc2=5.338454722e-08 ppdiblc2=-9.674644857e-15
+  pdiblcb=-3.881799574e+01 lpdiblcb=7.634924848e-06 wpdiblcb=1.620301054e-05 ppdiblcb=-3.221733088e-12
+  drout=1.046597409e+00 ldrout=-8.877738664e-09 wdrout=-2.428982380e-08 pdrout=4.627697372e-15
+  pscbe1=1.300187946e+09 lpscbe1=-1.102782544e+02 wpscbe1=-2.008030871e+02 ppscbe1=4.426900774e-5
+  pscbe2=-1.171276176e-07 lpscbe2=2.389591237e-14 wpscbe2=5.034588644e-14 ppscbe2=-9.502098016e-21
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=3.116248542e-01 lbeta0=1.234252074e-06 wbeta0=5.312758529e-06 pbeta0=-8.904785090e-13
* Gidl Induced Drain Leakage Model Parameters
+  agidl=-1.051956015e-13 lagidl=2.004186600e-20 wagidl=4.221204940e-20 pagidl=-8.042239652e-27
+  bgidl=1.000001385e+09 lbgidl=-2.636625071e-04 wbgidl=-5.558318348e-04 pbgidl=1.058003817e-10
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-1.106e-8
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-1.269288625e+01 lkt1=2.494462196e-06 wkt1=5.487475320e-06 pkt1=-1.141736926e-12
+  kt2=8.806944199e-01 lkt2=-2.116433718e-07 wkt2=-3.539635255e-07 pkt2=8.130528254e-14
+  at=-2.717015847e+06 lat=5.392095215e-01 wat=1.305422066e+00 pat=-2.545217758e-7
+  ute=-3.946837913e+00 lute=7.208586955e-07 wute=7.459698082e-07 pute=-1.421221680e-13
+  ua1=1.207210285e-09 lua1=-1.472622934e-16 wua1=-1.769476401e-15 pua1=3.684292741e-22
+  ub1=-5.148958533e-19 lub1=-3.577719454e-26 wub1=1.971743186e-24 pub1=-3.700608870e-31
+  uc1=-5.029437159e-11 luc1=2.603925173e-17 wuc1=5.909074261e-17 puc1=-2.419101634e-23
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.04e-6
+  sbref=1.04e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.189 pmos
* Model Flag Parameters
+  lmin=2.0e-05 lmax=0.0001 wmin=3.6e-07 wmax=4.2e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.126311+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+  k1=0.43165561
+  k2=0.026980026
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=3.2465718e-7
+  voff={-0.23051772+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.8768912+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+  eta0=0.08
+  etab=-0.07
+  u0=0.0095864
+  ua=-7.4757916e-10
+  ub=9.5046395e-19
+  uc=-1.0566299e-10
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=80156.0
+  a0=1.464
+  ags=0.11329
+  a1=0.0
+  a2=0.97
+  b0=-8.9873e-8
+  b1=3.3859e-9
+  keta=0.023361259
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=0.015
+  pdiblc1=0.39
+  pdiblc2=0.0012771588
+  pdiblcb=-0.225
+  drout=0.56
+  pscbe1=800000000.0
+  pscbe2=1.0060625e-8
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=0.0
+  alpha1=0.0
+  beta0=30.0
* Gidl Induced Drain Leakage Model Parameters
+  agidl=9.43573999999999e-11
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-0.43825
+  kt2=-0.058546
+  at=70990.0
+  ute=-0.08298
+  ua1=2.0902e-9
+  ub1=-1.2289e-18
+  uc1=-2.9789e-11
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.190 pmos
* Model Flag Parameters
+  lmin=8.0e-06 lmax=2.0e-05 wmin=3.6e-07 wmax=4.2e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.147214944e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=4.185705429e-7
+  k1=4.317678323e-01 lk1=-2.247085463e-9
+  k2=2.369023370e-02 lk2=6.587322199e-8
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=-6.144535039e-06 lcit=1.295359998e-10 wcit=8.470329473e-28 pcit=-2.202285663e-32
+  voff={-2.555024598e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=5.002824373e-7
+  nfactor={1.336645066e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.081762928e-5
+  eta0=0.08
+  etab=-0.07
+  u0=1.036751642e-02 lu0=-1.564070020e-8
+  ua=-8.705087603e-10 lua=2.461483309e-15 wua=-4.135903063e-31
+  ub=1.285196017e-18 lub=-6.702514248e-24
+  uc=-1.028248838e-10 luc=-5.682887705e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=80156.0
+  a0=1.509332888e+00 la0=-9.077239895e-7
+  ags=1.050124019e-01 lags=1.657466518e-7
+  a1=0.0
+  a2=0.97
+  b0=-1.368293135e-07 lb0=9.402306834e-13
+  b1=5.128942857e-09 lb1=-3.490185351e-14 pb1=-1.323488980e-35
+  keta=2.267780086e-02 lketa=1.368523780e-8
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=1.339372874e-02 lpclm=3.216320472e-8
+  pdiblc1=0.39
+  pdiblc2=6.725898845e-05 lpdiblc2=2.422645307e-8
+  pdiblcb=-0.225
+  drout=0.56
+  pscbe1=8.935747834e+08 lpscbe1=-1.873696547e+3
+  pscbe2=1.029619414e-08 lpscbe2=-4.716923448e-15
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=0.0
+  alpha1=0.0
+  beta0=30.0
* Gidl Induced Drain Leakage Model Parameters
+  agidl=1.354000851e-10 lagidl=-8.218190262e-16
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-3.929237983e-01 lkt1=-9.075901069e-7
+  kt2=-6.276904603e-02 lkt2=8.456024658e-08 wkt2=-2.775557562e-23
+  at=1.117695404e+05 lat=-8.165499428e-1
+  ute=5.541677232e-01 lute=-1.275794018e-05 wute=-5.551115123e-23 pute=-4.440892099e-28
+  ua1=3.163024859e-09 lua1=-2.148173002e-14
+  ub1=-1.868595191e-18 lub1=1.280894945e-23
+  uc1=-8.457025143e-11 luc1=1.096913484e-15 wuc1=1.292469707e-32 puc1=1.033975766e-37
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.191 pmos
* Model Flag Parameters
+  lmin=4.0e-06 lmax=8.0e-06 wmin=3.6e-07 wmax=4.2e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.065707492e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-2.354061279e-7
+  k1=4.412289030e-01 lk1=-7.815817575e-8
+  k2=3.495799846e-02 lk2=-2.453391399e-8
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.56
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-1.593357517e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-2.713130682e-7
+  nfactor={3.443981194e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-6.090624299e-6
+  eta0=0.08
+  etab=-0.07
+  u0=6.203732179e-03 lu0=1.776750591e-8
+  ua=-5.401640296e-10 lua=-1.890442437e-16
+  ub=3.885688924e-20 lub=3.297512674e-24
+  uc=-1.127146385e-10 luc=2.252176784e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=1.056489483e+05 lvsat=-2.045431804e-1
+  a0=1.533769379e+00 la0=-1.103790667e-6
+  ags=5.785621586e-02 lags=5.441052533e-7
+  a1=0.0
+  a2=1.140999600e+00 la2=-1.372018711e-6
+  b0=1.282581228e-08 lb0=-2.605302117e-13 pb0=-5.293955920e-35
+  b1=-3.358168040e-10 lb1=8.944754923e-15 pb1=-1.654361225e-36
+  keta=3.518549277e-02 lketa=-8.667047844e-8
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-3.101583599e-01 lpclm=2.628189859e-06 ppclm=-1.110223025e-28
+  pdiblc1=0.39
+  pdiblc2=5.609577701e-03 lpdiblc2=-2.024245196e-8
+  pdiblcb=-0.225
+  drout=0.56
+  pscbe1=5.192756498e+08 lpscbe1=1.129500038e+3
+  pscbe2=9.865934732e-09 lpscbe2=-1.264728462e-15
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=0.0
+  alpha1=0.0
+  beta0=30.0
* Gidl Induced Drain Leakage Model Parameters
+  agidl=4.485261892e-11 lagidl=-9.530962023e-17
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-5.943462052e-01 lkt1=7.085266035e-7
+  kt2=-4.587686192e-02 lkt2=-5.097453045e-8
+  at=-5.134862120e+04 lat=4.922318892e-01 pat=2.910383046e-23
+  ute=-1.954187970e+00 lute=7.367901890e-6
+  ua1=-1.128274578e-09 lua1=1.294959683e-14 pua1=1.654361225e-36
+  ub1=5.895975724e-19 lub1=-6.914409353e-24
+  uc1=1.345547543e-10 luc1=-6.612403822e-16
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.192 pmos
* Model Flag Parameters
+  lmin=2.0e-06 lmax=4.0e-06 wmin=3.6e-07 wmax=4.2e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.177416073e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=2.140555794e-7
+  k1=3.711821211e-01 lk1=2.036764523e-7
+  k2=3.190923688e-02 lk2=-1.226716077e-8
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=8.635280000e-01 ldsub=-1.221250979e-6
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.834912171e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=2.282289298e-7
+  nfactor={9.359981820e-01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=4.000295510e-6
+  eta0=1.604349200e-01 leta0=-3.236315093e-7
+  etab=-1.403173200e-01 letab=2.829231434e-7
+  u0=1.512830265e-02 lu0=-1.814068186e-8
+  ua=-1.062723639e-10 lua=-1.934816038e-15
+  ub=1.008693279e-18 lub=-6.046434356e-25
+  uc=-1.456246116e-10 luc=1.549357029e-16
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=5.896562096e+04 lvsat=-1.671187928e-2
+  a0=1.289551051e+00 la0=-1.211733363e-7
+  ags=1.053579842e-01 lags=3.529809385e-7
+  a1=0.0
+  a2=0.8
+  b0=-1.415557949e-07 lb0=3.606272723e-13
+  b1=-7.730386343e-08 lb1=3.186272299e-13 wb1=-1.323488980e-29 pb1=9.926167351e-36
+  keta=2.853443412e-02 lketa=-5.990981094e-8
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=4.782205445e-02 lpclm=1.187848502e-6
+  pdiblc1=0.39
+  pdiblc2=7.288412547e-04 lpdiblc2=-6.047112557e-10
+  pdiblcb=-0.225
+  drout=0.56
+  pscbe1=800000000.0
+  pscbe2=9.727100183e-09 lpscbe2=-7.061248733e-16
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=-1.011760000e-10 lalpha0=4.070836595e-16
+  alpha1=-1.011760000e-10 lalpha1=4.070836595e-16
+  beta0=5.568075730e+01 lbeta0=-1.033270406e-4
* Gidl Induced Drain Leakage Model Parameters
+  agidl=3.027630938e-11 lagidl=-3.666154729e-17 wagidl=-1.292469707e-32
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-2.990747896e-01 lkt1=-4.795038425e-7
+  kt2=-6.493627616e-02 lkt2=2.571140394e-8
+  at=1.326972424e+05 lat=-2.482803239e-1
+  ute=8.310287392e-01 lute=-3.838473242e-06 wute=1.110223025e-22 pute=-4.440892099e-28
+  ua1=3.743941955e-09 lua1=-6.653863832e-15 pua1=-3.308722450e-36
+  ub1=-1.995705145e-18 lub1=3.487607836e-24
+  uc1=-1.126835086e-10 luc1=3.335277131e-16 wuc1=-2.584939414e-32
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.193 pmos
* Model Flag Parameters
+  lmin=1.0e-06 lmax=2.0e-06 wmin=3.6e-07 wmax=4.2e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.029681593e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-8.488809500e-8
+  k1=4.627367281e-01 lk1=1.841387386e-8
+  k2=4.289505226e-02 lk2=-3.449717790e-8
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=-4.974048000e-01 ldsub=1.532623761e-6
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-1.339695087e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-7.433123756e-8
+  nfactor={3.109198808e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-3.972194201e-7
+  eta0=-2.241626400e-01 leta0=4.546093453e-07 weta0=3.599551213e-23 peta0=6.331740687e-29
+  etab=8.652602975e-01 letab=-1.751883277e-06 wetab=7.502679034e-23 petab=-6.331740687e-29
+  u0=4.588180664e-03 lu0=3.187465775e-9
+  ua=-8.807161675e-10 lua=-3.677135132e-16
+  ub=1.541802277e-19 lub=1.124480813e-24
+  uc=-8.449191963e-11 luc=3.123247804e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=6.140648349e+04 lvsat=-2.165101343e-2
+  a0=1.332090813e+00 la0=-2.072533974e-7
+  ags=-2.559368078e-01 lags=1.084068176e-6
+  a1=0.0
+  a2=0.8
+  b0=1.400825549e-07 lb0=-2.092735612e-13 wb0=2.646977960e-29 pb0=-2.646977960e-35
+  b1=1.599963470e-07 lb1=-1.615544920e-13
+  keta=1.204075832e-02 lketa=-2.653452808e-08 wketa=-8.673617380e-25 pketa=3.469446952e-30
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=8.732362441e-01 lpclm=-4.823936187e-7
+  pdiblc1=3.913823559e-01 lpdiblc1=-2.797224764e-9
+  pdiblc2=0.00043
+  pdiblcb=-0.225
+  drout=2.685397836e-01 ldrout=5.897755770e-7
+  pscbe1=800000000.0
+  pscbe2=9.667507287e-09 lpscbe2=-5.855374581e-16
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.236495401e-10 lalpha0=-4.785531742e-17
+  alpha1=3.047040000e-10 lalpha1=-4.142226381e-16
+  beta0=2.936091465e+00 lbeta0=3.402845599e-6
* Gidl Induced Drain Leakage Model Parameters
+  agidl=1.769389851e-11 lagidl=-1.120078725e-17
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-6.107671952e-01 lkt1=1.512119740e-7
+  kt2=-5.309487440e-02 lkt2=1.750090646e-9
+  at=-2.046302576e+04 lat=6.164254189e-2
+  ute=-1.123524176e+00 lute=1.166036726e-7
+  ua1=1.544285637e-09 lua1=-2.202815278e-15
+  ub1=-1.736591710e-18 lub1=2.963286619e-24 wub1=1.925929944e-40 pub1=-3.851859889e-46
+  uc1=-4.129082560e-12 luc1=1.138656610e-16
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=2.75e-6
+  sbref=2.74e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.194 pmos
* Model Flag Parameters
+  lmin=5.0e-07 lmax=1.0e-06 wmin=3.6e-07 wmax=4.2e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.136926034e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=2.487873503e-8
+  k1=4.604084761e-01 lk1=2.079688639e-8
+  k2=1.213770125e-02 lk2=-3.016414004e-9
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=1.774809600e+00 ldsub=-7.930331218e-07 wdsub=8.881784197e-22
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-2.112824992e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=4.800154470e-9
+  nfactor={2.153255836e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=5.812073306e-7
+  eta0=-6.270080000e-02 leta0=2.893499228e-7
+  etab=-1.732537571e+00 letab=9.070147972e-7
+  u0=9.597196877e-03 lu0=-1.939362499e-9
+  ua=-8.808370178e-10 lua=-3.675898204e-16
+  ub=1.032927229e-18 lub=2.250656827e-25
+  uc=-9.212753610e-11 luc=3.904768421e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=-3.876606176e+04 lvsat=8.087759009e-02 pvsat=1.455191523e-23
+  a0=1.430417848e+00 la0=-3.078930841e-7
+  ags=3.354234688e-01 lags=4.787991056e-7
+  a1=0.0
+  a2=6.220032000e-01 la2=1.821832847e-7
+  b0=-1.317925293e-07 lb0=6.899602493e-14
+  b1=4.409938272e-09 lb1=-2.308690884e-15
+  keta=2.121464773e-03 lketa=-1.638193275e-8
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=7.820070632e-01 lpclm=-3.890187274e-07 ppclm=1.110223025e-28
+  pdiblc1=7.819323543e-01 lpdiblc1=-4.025329592e-7
+  pdiblc2=8.520880000e-04 lpdiblc2=-4.320155098e-10
+  pdiblcb=-3.557815468e-01 lpdiblcb=1.338575288e-7
+  drout=6.822228327e-01 ldrout=1.663627026e-7
+  pscbe1=800000000.0
+  pscbe2=9.040301580e-09 lpscbe2=5.642012712e-17
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=5.270091976e-11 lalpha0=2.476201449e-17
+  alpha1=-3.094080000e-10 lalpha1=2.143332762e-16 walpha1=1.033975766e-31
+  beta0=4.265741962e+00 lbeta0=2.041921722e-6
* Gidl Induced Drain Leakage Model Parameters
+  agidl=6.602877830e-12 lagidl=1.510942430e-19
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-4.202584160e-01 lkt1=-4.377757166e-8
+  kt2=-4.284220064e-02 lkt2=-8.743726001e-9
+  at=-2.366748480e+03 lat=4.312064016e-2
+  ute=-1.890160640e+00 lute=9.012714263e-7
+  ua1=-2.628498262e-09 lua1=2.068112498e-15 wua1=-4.135903063e-31 pua1=2.067951531e-37
+  ub1=3.207248934e-18 lub1=-2.096833157e-24 wub1=7.703719778e-40 pub1=3.851859889e-46
+  uc1=2.897960218e-10 luc1=-1.869725618e-16 wuc1=1.033975766e-31
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.75e-6
+  sbref=1.74e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.195 pmos
* Model Flag Parameters
+  lmin=2.5e-07 lmax=5.0e-07 wmin=3.6e-07 wmax=4.2e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.132204410e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=2.240687043e-8
+  k1=1.155532129e-01 lk1=2.013355138e-7
+  k2=1.603779611e-01 lk2=-8.062315484e-08 pk2=6.938893904e-30
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=-1.799686157e-01 ldsub=2.303323697e-7
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-3.752999542e-03+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-1.038456892e-7
+  nfactor={4.013671651e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-3.927575568e-7
+  eta0=0.49
+  etab=-6.25e-6
+  u0=1.002403078e-02 lu0=-2.162818586e-9
+  ua=-4.159919914e-10 lua=-6.109454887e-16
+  ub=4.891119397e-19 lub=5.097638630e-25
+  uc=-3.701401147e-11 luc=1.019465179e-17
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=5.828170592e+04 lvsat=3.007114276e-2
+  a0=4.877951562e-01 la0=1.855887477e-7
+  ags=1.25
+  a1=0.0
+  a2=1.536190831e+00 la2=-2.964122239e-7
+  b0=0.0
+  b1=0.0
+  keta=-3.021165609e-02 lketa=5.451026823e-10
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=-8.229209877e-01 lpclm=4.511932058e-07 ppclm=4.163336342e-29
+  pdiblc1=-1.781362003e-01 lpdiblc1=1.000821305e-07 ppdiblc1=1.040834086e-29
+  pdiblc2=-7.267940052e-03 lpdiblc2=3.818981576e-09 wpdiblc2=9.215718466e-25 ppdiblc2=4.607859233e-31
+  pdiblcb=3.656309366e-02 lpdiblcb=-7.154273738e-8
+  drout=1.002074047e+00 ldrout=-1.085805324e-9
+  pscbe1=8.000344088e+08 lpscbe1=-1.801370335e-2
+  pscbe2=8.962724207e-09 lpscbe2=9.703343354e-17
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=7.160540337e+00 lbeta0=5.264368771e-7
* Gidl Induced Drain Leakage Model Parameters
+  agidl=1.443133138e-11 lagidl=-3.947257759e-18
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-3.892904371e-01 lkt1=-5.998992796e-8
+  kt2=-7.837421088e-02 lkt2=9.857992000e-9
+  at=5.260314272e+04 lat=1.434280272e-2
+  ute=1.119549344e-01 lute=-1.468761193e-07 pute=-2.775557562e-29
+  ua1=2.447237866e-09 lua1=-5.891368794e-16
+  ub1=-1.730805103e-18 lub1=4.883368922e-25
+  uc1=-7.721103712e-11 luc1=5.162973673e-18
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.1e-6
+  sbref=1.1e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.196 pmos
* Model Flag Parameters
+  lmin=1.8e-07 lmax=2.5e-07 wmin=3.6e-07 wmax=4.2e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-1.176e-8
+  vth0={-1.050284+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+  k1=0.85164386
+  k2=-0.1343835
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=0.66213569
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={-0.38341697+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+  nfactor={2.5777344+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+  eta0=0.49
+  etab=-6.25e-6
+  u0=0.00211668
+  ua=-2.649633e-9
+  ub=2.3528289e-18
+  uc=2.58041e-13
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=168223.0
+  a0=1.166315
+  ags=1.25
+  a1=0.0
+  a2=0.45249595
+  b0=0.0
+  b1=0.0
+  keta=-0.028218739
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=0.82665932
+  pdiblc1=0.18776805
+  pdiblc2=0.0066944085
+  pdiblcb=-0.225
+  drout=0.9981043
+  pscbe1=799968550.0
+  pscbe2=9.3174823e-9
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=9.0852145
* Gidl Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=1000000000.0
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-2.56e-9
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=-0.608616
+  kt2=-0.042333
+  at=105041.0
+  ute=-0.42503
+  ua1=2.9333e-10
+  ub1=5.4574e-20
+  uc1=-5.8335e-11
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.1e-6
+  sbref=1.1e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.197 pmos
* Model Flag Parameters
+  lmin=1.5e-07 lmax=1.8e-07 wmin=3.6e-07 wmax=4.2e-7
+  level=54.0
+  version=4.5
+  binunit=2.0
+  mobmod=0.0
+  capmod=2.0
+  igcmod=0.0
+  igbmod=0.0
+  geomod=0.0
+  diomod=1.0
+  rdsmod=0.0
+  rbodymod=1.0
+  rgatemod=0.0
+  permod=1.0
+  acnqsmod=0.0
+  trnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  tempmod=0.0
* Process Parameters
+  toxe={4.23e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*1.0*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+  toxm=4.23e-9
+  dtox=0.0
+  epsrox=3.9
+  xj=1.5e-7
+  ngate=1.0e+23
+  ndep=1.7e+17
+  nsd=1.0e+20
+  rsh=1.0
+  rshg=0.1
* Basic Model Parameters
+  wint=9.364e-9
+  lint=-2.026e-8
+  vth0={-2.280380644e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0=-1.813216737e-07 wvth0=-2.702289094e-07 pvth0=5.959087909e-14
+  k1=-1.942612612e+00 lk1=6.161894372e-07 wk1=8.145174970e-07 pk1=-1.796173984e-13
+  k2=-8.663270902e-02 lk2=-1.053000443e-08 wk2=1.525480424e-07 pk2=-3.363989431e-14
+  k3=-13.778
+  k3b=2.0
+  w0=0.0
+  dvt0=4.05
+  dvt1=0.3
+  dvt2=0.03
+  dvt0w=-4.254
+  dvt1w=1147200.0
+  dvt2w=-0.00896
+  dsub=7.017835139e+00 ldsub=-1.401558843e-06 wdsub=-2.103771966e-06 pdsub=4.639237939e-13
+  minv=0.0
+  voffl=0.0
+  lpe0=0.0
+  lpeb=0.0
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
+  phin=0.0
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  cit=1.0e-5
+  voff={6.584120060e-02+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff=-9.907041178e-08 wvoff=-1.970736678e-07 pvoff=4.345868523e-14
+  nfactor={1.712485402e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor=-3.207930818e-06 wnfactor=-6.027905788e-06 pnfactor=1.329273784e-12
+  eta0=8.400758601e+00 leta0=-1.744480487e-06 weta0=-3.174365925e-06 peta0=7.000111738e-13
+  etab=4.590023598e-01 letab=-1.012205786e-07 wetab=-1.826105146e-07 petab=4.026927068e-14
+  u0=-3.433624693e-03 lu0=1.223953191e-09 wu0=-1.558842911e-09 pu0=3.437560387e-16
+  ua=-3.435785141e-09 lua=1.733622700e-16 wua=-1.134355920e-15 pua=2.501481675e-22
+  ub=2.657584049e-18 lub=-6.720460536e-26 wub=1.066698111e-24 pub=-2.352282675e-31
+  uc=-3.742083373e-10 luc=8.257732575e-17 wuc=1.997496245e-16 puc=-4.404878720e-23
+  ud=0.0
+  up=0.0
+  lp=1.0
+  eu=1.67
+  vtl=0.0
+  xn=3.0
+  vsat=3.929098756e+06 lvsat=-8.293483216e-01 wvsat=-1.364313490e+00 pvsat=3.008584108e-7
+  a0=1.977516561e+00 la0=-1.788861682e-07 wa0=8.563083787e-08 pa0=-1.888331237e-14
+  ags=1.249999985e+00 lags=3.332713661e-15 wags=6.064414748e-15 pags=-1.337324473e-21
+  a1=0.0
+  a2=-9.073383837e+00 la2=2.100647011e-06 wa2=3.359617749e-06 pa2=-7.408629060e-13
+  b0=0.0
+  b1=0.0
+  keta=-1.610291043e+00 lketa=3.488785845e-07 wketa=6.068560841e-07 pketa=-1.338239037e-13
+  dwg=-5.722e-9
+  dwb=-1.7864e-8
+  pclm=2.179197569e+00 lpclm=-2.982617346e-07 wpclm=-2.774589244e-08 ppclm=6.118524200e-15
+  pdiblc1=1.164651831e-01 lpdiblc1=1.572370822e-08 wpdiblc1=9.110370374e-08 ppdiblc1=-2.009018875e-14
+  pdiblc2=6.689112786e-02 lpdiblc2=-1.327458055e-08 wpdiblc2=-1.653930299e-08 ppdiblc2=3.647247095e-15
+  pdiblcb=-9.631244073e+00 lpdiblcb=2.074264943e-06 wpdiblcb=4.491184323e-06 ppdiblcb=-9.903959668e-13
+  drout=9.860653258e-01 ldrout=2.654834583e-09 wdrout=6.165500110e-15 pdrout=-1.359615975e-21
+  pscbe1=1.299183743e+09 lpscbe1=-1.100869344e+02 wpscbe1=-2.004001287e+02 ppscbe1=4.419223639e-5
+  pscbe2=1.579775404e-08 lpscbe2=-1.429029524e-15 wpscbe2=-2.993343308e-15 ppscbe2=6.600920663e-22
+  pvag=0.0
+  delta=0.01
+  fprout=0.0
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
+  lambda=0.0
+  lc=5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+  rdsw=531.92
+  rsw=0.0
+  rdw=0.0
+  rdswmin=0.0
+  rdwmin=0.0
+  rswmin=0.0
+  prwb=-0.32348
+  prwg=0.02
+  wr=1.0
* Impact Ionization Current Model Parameters
+  alpha0=1.0e-10
+  alpha1=1.0e-10
+  beta0=2.366162204e+01 lbeta0=-3.214389391e-06 wbeta0=-4.056941542e-06 pbeta0=8.946367488e-13
* Gidl Induced Drain Leakage Model Parameters
+  agidl=0.0
+  bgidl=1.000000011e+09 lbgidl=-2.319414139e-06 wbgidl=-4.220550537e-06 pbgidl=9.307160378e-13
+  cgidl=300.0
+  egidl=0.1
* Gate Dielectric Tunneling Current Model Parameters
+  toxref=4.23e-9
+  dlcig=0.0
+  aigbacc=0.43
+  bigbacc=0.054
+  cigbacc=0.075
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  nigc=1.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  vfbsdoff=0.0
* Charge AND Capacitance Model Parameters
+  dlc=-1.106e-8
+  dwc=0.0
+  xpart=0.0
+  cgso=5.93202e-11
+  cgdo=5.93202e-11
+  cgbo=0.0
+  cgdl=7.513892e-12
+  cgsl=7.513892e-12
+  clc=1.0e-7
+  cle=0.6
+  cf=1.2e-11
+  ckappas=0.6
+  vfbcv=-0.1446893
+  acde=0.552
+  moin=14.504
+  noff=4.0
+  voffcv=-0.1375
* High-Speed/RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* Flicker AND Thermal Noise Model Parameters
+  ef=0.88
+  noia=1.2e+41
+  noib=2.0e+25
+  noic=0.0
+  em=41000000.0
+  ntnoi=1.0
+  lintnoi=-6.0e-8
+  af=1.0
+  kf=0.0
+  tnoia=1.5
+  tnoib=3.5
+  rnoia=0.577
+  rnoib=0.37
* Layout-Dependent Parasitics Model Parameters
+  xl=0.0
+  xw=0.0
+  dmcg=0.0
+  dmdg=0.0
+  dmcgt=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+  jss=2.17e-5
+  jsws=8.2e-10
+  ijthsfwd=0.1
+  ijthsrev=0.1
+  bvs=12.8
+  xjbvs=1.0
+  pbs=0.6587
+  cjs=0.0007432633326
+  mjs=0.34629
+  pbsws=0.7418
+  cjsws=9.5078641e-11
+  mjsws=0.26859
+  pbswgs=1.3925
+  cjswgs=2.54074486e-10
+  mjswgs=0.70393
* Temperature Dependence Parameters
+  tnom=30.0
+  kt1=1.445498355e+01 lkt1=-3.321824974e-06 wkt1=-5.406204692e-06 pkt1=1.192176259e-12
+  kt2=1.150606588e+00 lkt2=-2.630670379e-07 wkt2=-4.622717210e-07 pkt2=1.019401599e-13
+  at=5.333259814e+04 lat=1.140273678e-02 wat=1.937588049e-01 pat=-4.272769165e-8
+  ute=-2.087825043e+00 lute=3.666795630e-07 wute=-3.973519291e-15 pute=8.762401915e-22
+  ua1=-6.016759380e-10 lua1=1.973667094e-16 wua1=-1.043621009e-15 pua1=2.301393049e-22
+  ub1=4.863660387e-18 lub1=-1.060499730e-24 wub1=-1.865208340e-25 pub1=4.113157431e-32
+  uc1=-9.773734095e-10 luc1=2.026663501e-16 wuc1=4.311016023e-16 puc1=-9.506652534e-23
+  kt1l=0.0
+  prt=0.0
+  tvoff=0.0
+  njs=1.2556
+  tpb=0.0019551
+  tcj=0.0012407
+  tpbsw=0.00014242
+  tcjsw=0.0
+  tpbswg=0.0
+  tcjswg=2.0e-12
+  xtis=2.0
+  tvfbsdoff=0.0
* DW AND DL Parameters
+  ll=0.0
+  wl=0.0
+  lln=1.0
+  wln=1.0
+  lw=0.0
+  ww=0.0
+  lwn=1.0
+  wwn=1.0
+  lwl=0.0
+  wwl=0.0
+  llc=0.0
+  wlc=0.0
+  lwc=0.0
+  wwc=0.0
+  lwlc=0.0
+  wwlc=0.0
* Stress Parameters
+  saref=1.04e-6
+  sbref=1.04e-6
+  kvth0=2.65e-8
+  lkvth0=0.0
+  wkvth0=2.5e-7
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  wlod=0.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0=4.5e-8
+  lku0=0.0
+  wku0=2.5e-7
+  pku0=0.0
+  tku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat=0.4
+  steta0=0.0
.ends sky130_fd_pr__pfet_01v8_hvt
* Well Proximity Effect Parameters
