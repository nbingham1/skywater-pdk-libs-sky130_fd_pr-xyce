* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param sky130_fd_pr__cap_vpp_04p4x04p6_l1m1m2_shieldpo_floatm3__slope=0.0
* statistics {
*   mismatch {
*     vary  sky130_fd_pr__cap_vpp_04p4x04p6_l1m1m2_shieldpo_floatm3__slope dist=gauss std=0.00731
*   }
* }
.subckt sky130_fd_pr__cap_vpp_04p4x04p6_l1m1m2_shieldpo_floatm3 c0 c1 b m3
.param mult=1.0
+  ctot_a={9.766e-15*sky130_fd_pr__cap_vpp_04p4x04p6_l1m1m2_shieldpo_floatm3__cor+1.15082/sqrt(mult/0.31785)*sky130_fd_pr__cap_vpp_04p4x04p6_l1m1m2_shieldpo_floatm3__slope*9.766e-15*sky130_fd_pr__cap_vpp_04p4x04p6_l1m1m2_shieldpo_floatm3__cor}
+  cm3_c0={1.386e-15*cm3m2_vpp}
+  cm3_c1={0.745e-15*cm3m2_vpp}
+  cpl2s={2.838e-15*cpl2s_vpp}
+  rat_m2=0.300
+  rat_m1=0.385
+  rat_li=0.280
+  rat_li2p=0.035
+  cap_m2={rat_m2*ctot_a}
+  cap_m1={rat_m1*ctot_a}
+  cap_li={rat_li*ctot_a}
+  cap_li2p={rat_li2p*ctot_a}
+  lm2=1.585
+  wm2=0.140
+  nfm2=24.0
+  nvia_c0=40.0
+  nvia_c1=18.0
+  lm1=1.665
+  wm1=0.140
+  nfm1=20.0
+  ncon_c0=42.0
+  ncon_c1=8.0
+  ll1=1.555
+  wl1=0.170
+  nfl1=20.0
+  nlicon=44.0
ccmvpp4p4x4p6_m3shield m3 c0 c={cm3_c0}
cm3_1 m3 c1 c={cm3_c1}
rm21 c0 a1 r={rm2*lm2/wm2*(1/3)*(1/nfm2)}
cm2 a1 c1 c={cap_m2}
rvia1 c0 d0 r={rcvia/nvia_c0}
rvia2 c1 d1 r={rcvia/nvia_c1}
rm11 d0 b1 r={rm1*lm1/wm1*(1/3)*(1/nfm1)}
cm1 b1 d1 c={cap_m1}
rcon1 d0 e0 r={rcl1/ncon_c0}
rcon2 d1 e1 r={rcl1/ncon_c1}
rli1 e0 f1 r={rl1*ll1/wl1*(1/3)*(1/nfl1)}
cli f1 e1 c={cap_li}
rlicon e0 g0 r={rcp1/nlicon}
rpoly g0 h0 r={rp1}
cpl2b h0 b c={cpl2s}
cl12p e1 h0 c={cap_li2p}
.ends sky130_fd_pr__cap_vpp_04p4x04p6_l1m1m2_shieldpo_floatm3
