* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 63
.param
+  sky130_fd_pr__nfet_01v8__toxe_mult=0.948
+  sky130_fd_pr__nfet_01v8__rshn_mult=1.0
+  sky130_fd_pr__nfet_01v8__overlap_mult=0.94816
+  sky130_fd_pr__nfet_01v8__lint_diff=1.21275e-8
+  sky130_fd_pr__nfet_01v8__wint_diff=-3.2175e-8
+  sky130_fd_pr__nfet_01v8__dlc_diff=12.773e-9
+  sky130_fd_pr__nfet_01v8__dwc_diff=-3.2175e-8
*
* sky130_fd_pr__nfet_01v8, Bin 000, W = 1.26, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__voff_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_0=-1.1625e-19
+  sky130_fd_pr__nfet_01v8__pditsd_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_0=5.3075e-11
+  sky130_fd_pr__nfet_01v8__vsat_diff_0=-35091.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_0=0.040393
+  sky130_fd_pr__nfet_01v8__vth0_diff_0=-0.10867
+  sky130_fd_pr__nfet_01v8__nfactor_diff_0=0.99193
+  sky130_fd_pr__nfet_01v8__u0_diff_0=-0.006001
+  sky130_fd_pr__nfet_01v8__eta0_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_0=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 001, W = 1.68, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__eta0_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_1=-5.7353e-20
+  sky130_fd_pr__nfet_01v8__pditsd_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_1=3.1406e-11
+  sky130_fd_pr__nfet_01v8__vsat_diff_1=-27431.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_1=0.037642
+  sky130_fd_pr__nfet_01v8__vth0_diff_1=-0.078099
+  sky130_fd_pr__nfet_01v8__nfactor_diff_1=1.041
+  sky130_fd_pr__nfet_01v8__u0_diff_1=-0.0051246
*
* sky130_fd_pr__nfet_01v8, Bin 002, W = 1.0, L = 1.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__nfactor_diff_2=1.2221
+  sky130_fd_pr__nfet_01v8__u0_diff_2=0.00091513
+  sky130_fd_pr__nfet_01v8__vth0_diff_2=-0.0069074
+  sky130_fd_pr__nfet_01v8__eta0_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_2=2.7806e-19
+  sky130_fd_pr__nfet_01v8__kt1_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_2=2.1701e-12
+  sky130_fd_pr__nfet_01v8__vsat_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_2=-0.18927
+  sky130_fd_pr__nfet_01v8__a0_diff_2=0.4
+  sky130_fd_pr__nfet_01v8__b0_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_2=-0.0045103
*
* sky130_fd_pr__nfet_01v8, Bin 003, W = 1.0, L = 2.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__keta_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_3=-0.0040338
+  sky130_fd_pr__nfet_01v8__nfactor_diff_3=0.90771
+  sky130_fd_pr__nfet_01v8__u0_diff_3=0.00015125
+  sky130_fd_pr__nfet_01v8__vth0_diff_3=-0.013159
+  sky130_fd_pr__nfet_01v8__eta0_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_3=2.5047e-19
+  sky130_fd_pr__nfet_01v8__kt1_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_3=-3.3276e-13
+  sky130_fd_pr__nfet_01v8__vsat_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_3=-0.070457
+  sky130_fd_pr__nfet_01v8__a0_diff_3=0.13825
+  sky130_fd_pr__nfet_01v8__b0_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_3=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 004, W = 1.0, L = 4.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__pdits_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_4=0.0042246
+  sky130_fd_pr__nfet_01v8__nfactor_diff_4=1.0788
+  sky130_fd_pr__nfet_01v8__u0_diff_4=-0.0015927
+  sky130_fd_pr__nfet_01v8__vth0_diff_4=-0.015085
+  sky130_fd_pr__nfet_01v8__eta0_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_4=1.1584e-19
+  sky130_fd_pr__nfet_01v8__kt1_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_4=6.7133e-12
+  sky130_fd_pr__nfet_01v8__vsat_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_4=-0.028272
+  sky130_fd_pr__nfet_01v8__a0_diff_4=0.060814
+  sky130_fd_pr__nfet_01v8__b0_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_4=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 005, W = 1.0, L = 8.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__pdits_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_5=0.0056805
+  sky130_fd_pr__nfet_01v8__nfactor_diff_5=0.83107
+  sky130_fd_pr__nfet_01v8__u0_diff_5=-0.0016848
+  sky130_fd_pr__nfet_01v8__vth0_diff_5=-0.010908
+  sky130_fd_pr__nfet_01v8__eta0_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_5=1.177e-19
+  sky130_fd_pr__nfet_01v8__kt1_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_5=7.1008e-12
+  sky130_fd_pr__nfet_01v8__vsat_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_5=-0.034049
+  sky130_fd_pr__nfet_01v8__a0_diff_5=0.059073
+  sky130_fd_pr__nfet_01v8__b0_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_5=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 006, W = 1.0, L = 0.15
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__pclm_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_6=0.038669
+  sky130_fd_pr__nfet_01v8__nfactor_diff_6=1.492
+  sky130_fd_pr__nfet_01v8__u0_diff_6=-0.0061621
+  sky130_fd_pr__nfet_01v8__vth0_diff_6=-0.091488
+  sky130_fd_pr__nfet_01v8__eta0_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_6=-1.6835e-19
+  sky130_fd_pr__nfet_01v8__kt1_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_6=4.536e-11
+  sky130_fd_pr__nfet_01v8__vsat_diff_6=-36968.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_6=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 007, W = 1.0, L = 0.18
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__tvoff_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_7=0.021665
+  sky130_fd_pr__nfet_01v8__nfactor_diff_7=0.84742
+  sky130_fd_pr__nfet_01v8__u0_diff_7=-0.0034651
+  sky130_fd_pr__nfet_01v8__vth0_diff_7=-0.067997
+  sky130_fd_pr__nfet_01v8__eta0_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_7=7.5328e-20
+  sky130_fd_pr__nfet_01v8__kt1_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_7=2.1924e-11
+  sky130_fd_pr__nfet_01v8__vsat_diff_7=-35764.0
+  sky130_fd_pr__nfet_01v8__a0_diff_7=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 008, W = 1.0, L = 0.25
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__a0_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_8=1.028e-11
+  sky130_fd_pr__nfet_01v8__tvoff_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_8=0.0075414
+  sky130_fd_pr__nfet_01v8__nfactor_diff_8=1.5686
+  sky130_fd_pr__nfet_01v8__u0_diff_8=-0.0013777
+  sky130_fd_pr__nfet_01v8__vth0_diff_8=-0.043813
+  sky130_fd_pr__nfet_01v8__eta0_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_8=3.8454e-19
+  sky130_fd_pr__nfet_01v8__kt1_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_8=-37066.0
*
* sky130_fd_pr__nfet_01v8, Bin 009, W = 1.0, L = 0.5
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__kt1_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_9=-1.3217e-20
+  sky130_fd_pr__nfet_01v8__vsat_diff_9=-23454.0
+  sky130_fd_pr__nfet_01v8__a0_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_9=1.0588e-11
+  sky130_fd_pr__nfet_01v8__tvoff_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_9=0.0058993
+  sky130_fd_pr__nfet_01v8__nfactor_diff_9=1.5632
+  sky130_fd_pr__nfet_01v8__u0_diff_9=-0.0025729
+  sky130_fd_pr__nfet_01v8__vth0_diff_9=-0.011525
+  sky130_fd_pr__nfet_01v8__eta0_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_9=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 010, W = 2.0, L = 0.15
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__ags_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_10=0.041517
+  sky130_fd_pr__nfet_01v8__ua_diff_10=2.7907e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_10=-7.431e-20
+  sky130_fd_pr__nfet_01v8__tvoff_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_10=-31379.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_10=-0.069966
+  sky130_fd_pr__nfet_01v8__pdits_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_10=1.0586
+  sky130_fd_pr__nfet_01v8__u0_diff_10=-0.004511
*
* sky130_fd_pr__nfet_01v8, Bin 011, W = 3.0, L = 1.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__pclm_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_11=0.90844
+  sky130_fd_pr__nfet_01v8__u0_diff_11=-8.1412e-5
+  sky130_fd_pr__nfet_01v8__ags_diff_11=-0.16008
+  sky130_fd_pr__nfet_01v8__keta_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_11=-0.0012493
+  sky130_fd_pr__nfet_01v8__ua_diff_11=3.3022e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_11=1.3668e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_11=0.025831
+  sky130_fd_pr__nfet_01v8__rdsw_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_11=0.0012222
+  sky130_fd_pr__nfet_01v8__pdits_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_11=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 012, W = 3.0, L = 2.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__pditsd_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_12=1.0714
+  sky130_fd_pr__nfet_01v8__u0_diff_12=-0.0028219
+  sky130_fd_pr__nfet_01v8__ags_diff_12=-0.023677
+  sky130_fd_pr__nfet_01v8__keta_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_12=0.0029922
+  sky130_fd_pr__nfet_01v8__ua_diff_12=1.1894e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_12=-8.5344e-20
+  sky130_fd_pr__nfet_01v8__tvoff_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_12=0.03384
+  sky130_fd_pr__nfet_01v8__rdsw_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_12=-0.011332
+  sky130_fd_pr__nfet_01v8__pdits_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_12=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 013, W = 3.0, L = 4.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__pdits_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_13=1.4703
+  sky130_fd_pr__nfet_01v8__u0_diff_13=-0.0040635
+  sky130_fd_pr__nfet_01v8__ags_diff_13=0.011298
+  sky130_fd_pr__nfet_01v8__keta_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_13=0.0052932
+  sky130_fd_pr__nfet_01v8__ua_diff_13=1.5958e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_13=-1.9512e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_13=0.014103
+  sky130_fd_pr__nfet_01v8__rdsw_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_13=-0.014516
+  sky130_fd_pr__nfet_01v8__b0_diff_13=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 014, W = 3.0, L = 8.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__b0_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_14=1.1989
+  sky130_fd_pr__nfet_01v8__u0_diff_14=-0.0029321
+  sky130_fd_pr__nfet_01v8__ags_diff_14=-0.0095841
+  sky130_fd_pr__nfet_01v8__keta_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_14=0.0064914
+  sky130_fd_pr__nfet_01v8__ua_diff_14=1.1147e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_14=-1.3332e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_14=0.035541
+  sky130_fd_pr__nfet_01v8__rdsw_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_14=-0.0089431
*
* sky130_fd_pr__nfet_01v8, Bin 015, W = 3.0, L = 0.15
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__kt1_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_15=-26551.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_15=-0.090092
+  sky130_fd_pr__nfet_01v8__b0_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_15=1.1928
+  sky130_fd_pr__nfet_01v8__u0_diff_15=-0.0073153
+  sky130_fd_pr__nfet_01v8__ags_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_15=0.047342
+  sky130_fd_pr__nfet_01v8__ua_diff_15=4.014e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_15=-4.9615e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_15=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 016, W = 3.0, L = 0.18
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__a0_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_16=-24194.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_16=-0.045047
+  sky130_fd_pr__nfet_01v8__b0_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_16=0.54872
+  sky130_fd_pr__nfet_01v8__u0_diff_16=-0.0031346
+  sky130_fd_pr__nfet_01v8__ags_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_16=0.033945
+  sky130_fd_pr__nfet_01v8__ua_diff_16=1.9692e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_16=4.519e-20
+  sky130_fd_pr__nfet_01v8__tvoff_diff_16=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 017, W = 3.0, L = 0.25
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__tvoff_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_17=-23827.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_17=-0.035942
+  sky130_fd_pr__nfet_01v8__pdits_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_17=1.25
+  sky130_fd_pr__nfet_01v8__u0_diff_17=-0.00047656
+  sky130_fd_pr__nfet_01v8__ags_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_17=0.016135
+  sky130_fd_pr__nfet_01v8__ua_diff_17=3.0188e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_17=1.7684e-19
*
* sky130_fd_pr__nfet_01v8, Bin 018, W = 3.0, L = 0.5
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__ub_diff_18=1.0996e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_18=-9502.5
+  sky130_fd_pr__nfet_01v8__vth0_diff_18=-0.01712
+  sky130_fd_pr__nfet_01v8__pdits_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_18=0.93684
+  sky130_fd_pr__nfet_01v8__u0_diff_18=-0.0013645
+  sky130_fd_pr__nfet_01v8__ags_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_18=0.0045237
+  sky130_fd_pr__nfet_01v8__ua_diff_18=6.0012e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_18=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 019, W = 5.0, L = 1.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__eta0_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_19=1.0534e-12
+  sky130_fd_pr__nfet_01v8__ub_diff_19=1.1911e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_19=0.01338
+  sky130_fd_pr__nfet_01v8__rdsw_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_19=0.0027696
+  sky130_fd_pr__nfet_01v8__pdits_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_19=0.86302
+  sky130_fd_pr__nfet_01v8__u0_diff_19=-0.00044898
+  sky130_fd_pr__nfet_01v8__ags_diff_19=-0.0031687
+  sky130_fd_pr__nfet_01v8__keta_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_19=0.004879
*
* sky130_fd_pr__nfet_01v8, Bin 020, W = 5.0, L = 2.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__ua_diff_20=1.7846e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_20=-2.4238e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_20=0.031901
+  sky130_fd_pr__nfet_01v8__rdsw_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_20=-0.015969
+  sky130_fd_pr__nfet_01v8__pdits_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_20=1.0179
+  sky130_fd_pr__nfet_01v8__u0_diff_20=-0.0040411
+  sky130_fd_pr__nfet_01v8__ags_diff_20=-0.011538
+  sky130_fd_pr__nfet_01v8__keta_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_20=0.0029706
*
* sky130_fd_pr__nfet_01v8, Bin 021, W = 5.0, L = 4.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__ags_diff_21=-0.034012
+  sky130_fd_pr__nfet_01v8__keta_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_21=0.0024091
+  sky130_fd_pr__nfet_01v8__ua_diff_21=1.1125e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_21=-1.5169e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_21=0.050141
+  sky130_fd_pr__nfet_01v8__rdsw_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_21=-0.010686
+  sky130_fd_pr__nfet_01v8__pdits_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_21=0.81902
+  sky130_fd_pr__nfet_01v8__u0_diff_21=-0.0026598
*
* sky130_fd_pr__nfet_01v8, Bin 022, W = 5.0, L = 8.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__pclm_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_22=1.1736
+  sky130_fd_pr__nfet_01v8__u0_diff_22=-0.0021258
+  sky130_fd_pr__nfet_01v8__ags_diff_22=0.017294
+  sky130_fd_pr__nfet_01v8__keta_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_22=0.0068712
+  sky130_fd_pr__nfet_01v8__ua_diff_22=8.0644e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_22=-6.0978e-20
+  sky130_fd_pr__nfet_01v8__tvoff_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_22=0.0028956
+  sky130_fd_pr__nfet_01v8__rdsw_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_22=-0.0065592
+  sky130_fd_pr__nfet_01v8__pdits_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_22=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 023, W = 5.0, L = 0.15
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__pditsd_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_23=1.5918
+  sky130_fd_pr__nfet_01v8__u0_diff_23=-0.0025309
+  sky130_fd_pr__nfet_01v8__ags_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_23=0.038594
+  sky130_fd_pr__nfet_01v8__ua_diff_23=1.3169e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_23=-8.3378e-20
+  sky130_fd_pr__nfet_01v8__tvoff_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_23=-19734.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_23=-0.071485
+  sky130_fd_pr__nfet_01v8__pdits_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_23=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 024, W = 5.0, L = 0.18
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__pdits_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_24=1.5765
+  sky130_fd_pr__nfet_01v8__u0_diff_24=-0.0098305
+  sky130_fd_pr__nfet_01v8__ags_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_24=0.031749
+  sky130_fd_pr__nfet_01v8__ua_diff_24=5.3365e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_24=-4.9047e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_24=-18507.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_24=-0.061419
+  sky130_fd_pr__nfet_01v8__b0_diff_24=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 025, W = 5.0, L = 0.25
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__b0_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_25=0.99413
+  sky130_fd_pr__nfet_01v8__u0_diff_25=-0.00035965
+  sky130_fd_pr__nfet_01v8__ags_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_25=0.014701
+  sky130_fd_pr__nfet_01v8__ua_diff_25=2.2831e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_25=1.9499e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_25=-19710.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_25=-0.017685
*
* sky130_fd_pr__nfet_01v8, Bin 026, W = 5.0, L = 0.5
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__kt1_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_26=-11407.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_26=-0.013166
+  sky130_fd_pr__nfet_01v8__b0_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_26=1.1139
+  sky130_fd_pr__nfet_01v8__u0_diff_26=-0.0010353
+  sky130_fd_pr__nfet_01v8__ags_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_26=0.0022571
+  sky130_fd_pr__nfet_01v8__ua_diff_26=3.58e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_26=3.3057e-20
+  sky130_fd_pr__nfet_01v8__tvoff_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_26=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 027, W = 7.0, L = 1.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__a0_diff_27=0.084507
+  sky130_fd_pr__nfet_01v8__rdsw_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_27=-0.013193
+  sky130_fd_pr__nfet_01v8__b0_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_27=0.95703
+  sky130_fd_pr__nfet_01v8__u0_diff_27=-0.001564
+  sky130_fd_pr__nfet_01v8__ags_diff_27=-0.075834
+  sky130_fd_pr__nfet_01v8__keta_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_27=0.003712
+  sky130_fd_pr__nfet_01v8__ua_diff_27=7.7409e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_27=3.1147e-20
+  sky130_fd_pr__nfet_01v8__tvoff_diff_27=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 028, W = 7.0, L = 2.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__tvoff_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_28=0.005117
+  sky130_fd_pr__nfet_01v8__rdsw_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_28=-0.0059123
+  sky130_fd_pr__nfet_01v8__pdits_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_28=0.9391
+  sky130_fd_pr__nfet_01v8__u0_diff_28=-0.0015284
+  sky130_fd_pr__nfet_01v8__ags_diff_28=0.0069276
+  sky130_fd_pr__nfet_01v8__keta_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_28=0.0043703
+  sky130_fd_pr__nfet_01v8__ua_diff_28=6.5911e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_28=1.4716e-20
*
* sky130_fd_pr__nfet_01v8, Bin 029, W = 7.0, L = 4.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__ub_diff_29=5.7406e-20
+  sky130_fd_pr__nfet_01v8__tvoff_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_29=-0.031005
+  sky130_fd_pr__nfet_01v8__rdsw_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_29=-0.0089838
+  sky130_fd_pr__nfet_01v8__pdits_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_29=0.84229
+  sky130_fd_pr__nfet_01v8__u0_diff_29=-0.0011415
+  sky130_fd_pr__nfet_01v8__ags_diff_29=0.030935
+  sky130_fd_pr__nfet_01v8__keta_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_29=0.0021451
+  sky130_fd_pr__nfet_01v8__ua_diff_29=4.9559e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_29=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 030, W = 7.0, L = 8.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__eta0_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_30=-2.815e-21
+  sky130_fd_pr__nfet_01v8__tvoff_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_30=-0.005506
+  sky130_fd_pr__nfet_01v8__rdsw_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_30=9.4355e-5
+  sky130_fd_pr__nfet_01v8__pdits_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_30=0.7784
+  sky130_fd_pr__nfet_01v8__u0_diff_30=-0.0010835
+  sky130_fd_pr__nfet_01v8__ags_diff_30=0.018208
+  sky130_fd_pr__nfet_01v8__keta_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_30=0.0043056
+  sky130_fd_pr__nfet_01v8__ua_diff_30=4.0515e-12
*
* sky130_fd_pr__nfet_01v8, Bin 031, W = 7.0, L = 0.15
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__ua_diff_31=1.7239e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_31=1.8943e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_31=-14812.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_31=-0.048201
+  sky130_fd_pr__nfet_01v8__pdits_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_31=-0.058235
+  sky130_fd_pr__nfet_01v8__u0_diff_31=0.00031791
+  sky130_fd_pr__nfet_01v8__ags_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_31=0.032412
*
* sky130_fd_pr__nfet_01v8, Bin 032, W = 7.0, L = 0.18
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__ags_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_32=0.030209
+  sky130_fd_pr__nfet_01v8__ua_diff_32=4.6597e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_32=-3.6939e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_32=-17879.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_32=-0.051364
+  sky130_fd_pr__nfet_01v8__pdits_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_32=1.4588
+  sky130_fd_pr__nfet_01v8__u0_diff_32=-0.0082299
*
* sky130_fd_pr__nfet_01v8, Bin 033, W = 7.0, L = 0.25
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__pclm_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_33=0.69099
+  sky130_fd_pr__nfet_01v8__u0_diff_33=-0.000468
+  sky130_fd_pr__nfet_01v8__ags_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_33=0.01592
+  sky130_fd_pr__nfet_01v8__ua_diff_33=3.2229e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_33=1.4018e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_33=-20786.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_33=-0.01658
+  sky130_fd_pr__nfet_01v8__pdits_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_33=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 034, W = 7.0, L = 0.5
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__pditsd_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_34=1.0312
+  sky130_fd_pr__nfet_01v8__u0_diff_34=-0.0010308
+  sky130_fd_pr__nfet_01v8__ags_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_34=0.0023487
+  sky130_fd_pr__nfet_01v8__ua_diff_34=3.7206e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_34=2.9272e-20
+  sky130_fd_pr__nfet_01v8__tvoff_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_34=-8888.2
+  sky130_fd_pr__nfet_01v8__kt1_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_34=-0.015053
+  sky130_fd_pr__nfet_01v8__pdits_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_34=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 035, W = 0.42, L = 1.0
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__pdits_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_35=9.7159e-9
+  sky130_fd_pr__nfet_01v8__pditsd_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_35=2.515
+  sky130_fd_pr__nfet_01v8__u0_diff_35=-0.003834
+  sky130_fd_pr__nfet_01v8__ags_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_35=0.0033794
+  sky130_fd_pr__nfet_01v8__ua_diff_35=1.5064e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_35=9.0683e-20
+  sky130_fd_pr__nfet_01v8__tvoff_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_35=-0.047761
+  sky130_fd_pr__nfet_01v8__b0_diff_35=1.8786e-8
*
* sky130_fd_pr__nfet_01v8, Bin 036, W = 0.42, L = 20.0
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__b0_diff_36=9.1484e-8
+  sky130_fd_pr__nfet_01v8__pdits_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_36=1.6098e-9
+  sky130_fd_pr__nfet_01v8__pditsd_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_36=0.98042
+  sky130_fd_pr__nfet_01v8__u0_diff_36=-0.002233
+  sky130_fd_pr__nfet_01v8__ags_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_36=0.0010001
+  sky130_fd_pr__nfet_01v8__ua_diff_36=8.3058e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_36=1.181e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_36=-0.0057401
*
* sky130_fd_pr__nfet_01v8, Bin 037, W = 0.42, L = 2.0
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__kt1_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_37=-0.066137
+  sky130_fd_pr__nfet_01v8__b0_diff_37=1.8557e-7
+  sky130_fd_pr__nfet_01v8__pdits_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_37=1.5528e-8
+  sky130_fd_pr__nfet_01v8__pditsd_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_37=1.8673
+  sky130_fd_pr__nfet_01v8__u0_diff_37=-0.0051091
+  sky130_fd_pr__nfet_01v8__ags_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_37=0.0048975
+  sky130_fd_pr__nfet_01v8__ua_diff_37=2.335e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_37=-2.9837e-20
+  sky130_fd_pr__nfet_01v8__tvoff_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_37=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 038, W = 0.42, L = 4.0
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__a0_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_38=-0.041505
+  sky130_fd_pr__nfet_01v8__b0_diff_38=9.9093e-8
+  sky130_fd_pr__nfet_01v8__pdits_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_38=1.362e-9
+  sky130_fd_pr__nfet_01v8__pditsd_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_38=1.4073
+  sky130_fd_pr__nfet_01v8__u0_diff_38=-0.0036085
+  sky130_fd_pr__nfet_01v8__ags_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_38=0.0098745
+  sky130_fd_pr__nfet_01v8__ua_diff_38=1.4848e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_38=1.0787e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_38=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 039, W = 0.42, L = 8.0
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__tvoff_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_39=-0.0082635
+  sky130_fd_pr__nfet_01v8__pdits_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_39=1.1142e-7
+  sky130_fd_pr__nfet_01v8__b1_diff_39=1.5277e-9
+  sky130_fd_pr__nfet_01v8__pditsd_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_39=0.9461
+  sky130_fd_pr__nfet_01v8__u0_diff_39=-0.0027345
+  sky130_fd_pr__nfet_01v8__ags_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_39=-0.0017247
+  sky130_fd_pr__nfet_01v8__ua_diff_39=1.0828e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_39=7.0155e-20
*
* sky130_fd_pr__nfet_01v8, Bin 040, W = 0.42, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__tvoff_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_40=-57437.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_40=-0.14897
+  sky130_fd_pr__nfet_01v8__pdits_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_40=-2.5003e-7
+  sky130_fd_pr__nfet_01v8__voff_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_40=2.2838e-8
+  sky130_fd_pr__nfet_01v8__pditsd_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_40=1.2701
+  sky130_fd_pr__nfet_01v8__u0_diff_40=-0.0010145
+  sky130_fd_pr__nfet_01v8__ags_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_40=0.033085
+  sky130_fd_pr__nfet_01v8__ua_diff_40=1.9284e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_40=8.61e-19
*
* sky130_fd_pr__nfet_01v8, Bin 041, W = 0.42, L = 0.18
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__eta0_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_41=2.6772e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_41=-9474.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_41=-0.13141
+  sky130_fd_pr__nfet_01v8__pdits_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_41=1.0704e-6
+  sky130_fd_pr__nfet_01v8__voff_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_41=1.6377e-8
+  sky130_fd_pr__nfet_01v8__pditsd_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_41=0.69719
+  sky130_fd_pr__nfet_01v8__u0_diff_41=-0.006133
+  sky130_fd_pr__nfet_01v8__ags_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_41=0.016032
+  sky130_fd_pr__nfet_01v8__ua_diff_41=4.4403e-11
*
* sky130_fd_pr__nfet_01v8, Bin 042, W = 0.42, L = 0.5
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__ua_diff_42=1.515e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_42=1.7745e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_42=6287.8
+  sky130_fd_pr__nfet_01v8__kt1_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_42=-0.045618
+  sky130_fd_pr__nfet_01v8__pdits_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_42=3.4771e-7
+  sky130_fd_pr__nfet_01v8__voff_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_42=5.442e-9
+  sky130_fd_pr__nfet_01v8__pditsd_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_42=1.724
+  sky130_fd_pr__nfet_01v8__u0_diff_42=-0.0033408
+  sky130_fd_pr__nfet_01v8__ags_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_42=0.0094315
*
* sky130_fd_pr__nfet_01v8, Bin 043, W = 0.55, L = 1.0
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__ags_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_43=0.011586
+  sky130_fd_pr__nfet_01v8__ua_diff_43=2.0363e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_43=2.8166e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_43=-0.025181
+  sky130_fd_pr__nfet_01v8__pdits_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_43=2.9678e-7
+  sky130_fd_pr__nfet_01v8__voff_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_43=7.2562e-9
+  sky130_fd_pr__nfet_01v8__pditsd_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_43=2.0375
+  sky130_fd_pr__nfet_01v8__u0_diff_43=-0.00084089
*
* sky130_fd_pr__nfet_01v8, Bin 044, W = 0.55, L = 2.0
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__pclm_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_44=1.5325
+  sky130_fd_pr__nfet_01v8__u0_diff_44=-0.0063868
+  sky130_fd_pr__nfet_01v8__ags_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_44=0.0039682
+  sky130_fd_pr__nfet_01v8__ua_diff_44=2.7076e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_44=-2.4014e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_44=-0.039391
+  sky130_fd_pr__nfet_01v8__pdits_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_44=2.0206e-7
+  sky130_fd_pr__nfet_01v8__voff_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_44=5.7041e-9
+  sky130_fd_pr__nfet_01v8__pditsd_diff_44=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 045, W = 0.55, L = 4.0
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__pditsd_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_45=1.49
+  sky130_fd_pr__nfet_01v8__u0_diff_45=-0.0039817
+  sky130_fd_pr__nfet_01v8__ags_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_45=0.0054607
+  sky130_fd_pr__nfet_01v8__ua_diff_45=1.6328e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_45=-3.3128e-20
+  sky130_fd_pr__nfet_01v8__tvoff_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_45=-0.022827
+  sky130_fd_pr__nfet_01v8__pdits_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_45=1.4014e-7
+  sky130_fd_pr__nfet_01v8__voff_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_45=3.2239e-9
*
* sky130_fd_pr__nfet_01v8, Bin 046, W = 0.55, L = 8.0
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__pdits_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_46=7.6808e-10
+  sky130_fd_pr__nfet_01v8__pditsd_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_46=0.64977
+  sky130_fd_pr__nfet_01v8__u0_diff_46=-0.0017403
+  sky130_fd_pr__nfet_01v8__ags_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_46=0.0020875
+  sky130_fd_pr__nfet_01v8__ua_diff_46=7.7949e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_46=1.8699e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_46=-0.0063547
+  sky130_fd_pr__nfet_01v8__b0_diff_46=9.4853e-8
*
* sky130_fd_pr__nfet_01v8, Bin 047, W = 0.55, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__b0_diff_47=4.5808e-7
+  sky130_fd_pr__nfet_01v8__pdits_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_47=1.6807e-8
+  sky130_fd_pr__nfet_01v8__pditsd_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_47=1.1215
+  sky130_fd_pr__nfet_01v8__u0_diff_47=-0.0059137
+  sky130_fd_pr__nfet_01v8__ags_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_47=0.035099
+  sky130_fd_pr__nfet_01v8__ua_diff_47=1.3878e-10
+  sky130_fd_pr__nfet_01v8__eta0_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_47=-1.9739e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_47=-47947.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_47=-0.15378
*
* sky130_fd_pr__nfet_01v8, Bin 048, W = 0.55, L = 0.5
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__kt1_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_48=-53290.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_48=-0.04144
+  sky130_fd_pr__nfet_01v8__b0_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_48=1.6886
+  sky130_fd_pr__nfet_01v8__u0_diff_48=-0.00069694
+  sky130_fd_pr__nfet_01v8__ags_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_48=0.0019981
+  sky130_fd_pr__nfet_01v8__ua_diff_48=6.8934e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_48=2.4766e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_48=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 049, W = 0.64, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__a0_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_49=-36934.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_49=-0.093996
+  sky130_fd_pr__nfet_01v8__b0_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_49=0.94211
+  sky130_fd_pr__nfet_01v8__u0_diff_49=-0.0040145
+  sky130_fd_pr__nfet_01v8__ags_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_49=0.03981
+  sky130_fd_pr__nfet_01v8__ua_diff_49=3.2111e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_49=2.0511e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_49=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 050, W = 0.84, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__tvoff_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_50=-31469.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_50=-0.12205
+  sky130_fd_pr__nfet_01v8__pdits_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_50=5.7064e-7
+  sky130_fd_pr__nfet_01v8__voff_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_50=-8.1551e-10
+  sky130_fd_pr__nfet_01v8__pditsd_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_50=0.571
+  sky130_fd_pr__nfet_01v8__u0_diff_50=-0.0053284
+  sky130_fd_pr__nfet_01v8__ags_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_50=0.035308
+  sky130_fd_pr__nfet_01v8__ua_diff_50=3.754e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_50=3.2112e-20
*
* sky130_fd_pr__nfet_01v8, Bin 051, W = 0.74, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__tvoff_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_51=-38324.63321946
+  sky130_fd_pr__nfet_01v8__kt1_diff_51=6.07518e-5
+  sky130_fd_pr__nfet_01v8__vth0_diff_51=-0.10491489
+  sky130_fd_pr__nfet_01v8__pdits_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_51=3.22831e-7
+  sky130_fd_pr__nfet_01v8__b1_diff_51=-4.61362e-10
+  sky130_fd_pr__nfet_01v8__voff_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_51=0.00033347
+  sky130_fd_pr__nfet_01v8__u0_diff_51=-0.0019502
+  sky130_fd_pr__nfet_01v8__nfactor_diff_51=0.34959259
+  sky130_fd_pr__nfet_01v8__keta_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_51=0.03502317
+  sky130_fd_pr__nfet_01v8__ua_diff_51=2.4186e-11
+  sky130_fd_pr__nfet_01v8__ub_diff_51=1.66053e-19
+  sky130_fd_pr__nfet_01v8__eta0_diff_51=-4.85723e-17
*
* sky130_fd_pr__nfet_01v8, Bin 052, W = 0.36, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__ub_diff_52=4.16095e-19
+  sky130_fd_pr__nfet_01v8__eta0_diff_52=3.2537e-5
+  sky130_fd_pr__nfet_01v8__tvoff_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_52=-65067.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_52=-0.12224
+  sky130_fd_pr__nfet_01v8__pdits_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_52=-7.39989e-7
+  sky130_fd_pr__nfet_01v8__b1_diff_52=2.7011e-8
+  sky130_fd_pr__nfet_01v8__voff_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_52=0.00091873
+  sky130_fd_pr__nfet_01v8__u0_diff_52=-0.0083504
+  sky130_fd_pr__nfet_01v8__nfactor_diff_52=0.5935569
+  sky130_fd_pr__nfet_01v8__keta_diff_52=0.00306555
+  sky130_fd_pr__nfet_01v8__ags_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_52=0.020341
+  sky130_fd_pr__nfet_01v8__ua_diff_52=-4.02468e-11
*
* sky130_fd_pr__nfet_01v8, Bin 053, W = 0.39, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__ua_diff_53=-4.99625e-12
+  sky130_fd_pr__nfet_01v8__ub_diff_53=3.05799e-19
+  sky130_fd_pr__nfet_01v8__eta0_diff_53=1.15988e-5
+  sky130_fd_pr__nfet_01v8__tvoff_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_53=-59191.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_53=-0.12953
+  sky130_fd_pr__nfet_01v8__pdits_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_53=-4.77112e-7
+  sky130_fd_pr__nfet_01v8__b1_diff_53=2.47721e-8
+  sky130_fd_pr__nfet_01v8__voff_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_53=0.00032751
+  sky130_fd_pr__nfet_01v8__u0_diff_53=-0.0072906
+  sky130_fd_pr__nfet_01v8__nfactor_diff_53=0.56383409
+  sky130_fd_pr__nfet_01v8__keta_diff_53=0.0010928
+  sky130_fd_pr__nfet_01v8__ags_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_53=0.022274
*
* sky130_fd_pr__nfet_01v8, Bin 054, W = 0.52, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__keta_diff_54=-0.00037717
+  sky130_fd_pr__nfet_01v8__ags_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_54=0.029985
+  sky130_fd_pr__nfet_01v8__ua_diff_54=1.04128e-10
+  sky130_fd_pr__nfet_01v8__ub_diff_54=-6.43431e-20
+  sky130_fd_pr__nfet_01v8__eta0_diff_54=-4.00316e-6
+  sky130_fd_pr__nfet_01v8__tvoff_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_54=-49054.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_54=-0.15398
+  sky130_fd_pr__nfet_01v8__pdits_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_54=3.24896e-7
+  sky130_fd_pr__nfet_01v8__b1_diff_54=1.79413e-8
+  sky130_fd_pr__nfet_01v8__voff_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_54=-0.00011304
+  sky130_fd_pr__nfet_01v8__u0_diff_54=-0.00048232
+  sky130_fd_pr__nfet_01v8__nfactor_diff_54=0.49466752
*
* sky130_fd_pr__nfet_01v8, Bin 055, W = 0.54, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__pclm_diff_55=-4.18441e-5
+  sky130_fd_pr__nfet_01v8__u0_diff_55=-0.00096228
+  sky130_fd_pr__nfet_01v8__nfactor_diff_55=0.48878058
+  sky130_fd_pr__nfet_01v8__keta_diff_55=-0.00013962
+  sky130_fd_pr__nfet_01v8__ags_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_55=0.031175
+  sky130_fd_pr__nfet_01v8__ua_diff_55=1.16564e-10
+  sky130_fd_pr__nfet_01v8__ub_diff_55=-1.09034e-19
+  sky130_fd_pr__nfet_01v8__eta0_diff_55=-1.48189e-6
+  sky130_fd_pr__nfet_01v8__tvoff_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_55=-47873.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_55=-0.14959
+  sky130_fd_pr__nfet_01v8__pdits_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_55=4.15269e-7
+  sky130_fd_pr__nfet_01v8__b1_diff_55=1.71716e-8
+  sky130_fd_pr__nfet_01v8__voff_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_55=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 056, W = 0.58, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__pditsd_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_56=-7.83128e-5
+  sky130_fd_pr__nfet_01v8__u0_diff_56=0.00065384
+  sky130_fd_pr__nfet_01v8__nfactor_diff_56=0.48174064
+  sky130_fd_pr__nfet_01v8__keta_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_56=0.030661
+  sky130_fd_pr__nfet_01v8__ua_diff_56=8.51462e-11
+  sky130_fd_pr__nfet_01v8__ub_diff_56=4.16055e-20
+  sky130_fd_pr__nfet_01v8__eta0_diff_56=2.77352e-6
+  sky130_fd_pr__nfet_01v8__tvoff_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_56=-48118.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_56=-3.99555e-5
+  sky130_fd_pr__nfet_01v8__vth0_diff_56=-0.14576
+  sky130_fd_pr__nfet_01v8__pdits_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_56=2.90133e-7
+  sky130_fd_pr__nfet_01v8__b1_diff_56=1.0645e-8
+  sky130_fd_pr__nfet_01v8__voff_diff_56=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 057, W = 0.6, L = 0.15
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__pdits_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_57=6.86799e-9
+  sky130_fd_pr__nfet_01v8__voff_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_57=-8.11826e-5
+  sky130_fd_pr__nfet_01v8__u0_diff_57=0.001579
+  sky130_fd_pr__nfet_01v8__nfactor_diff_57=0.47867486
+  sky130_fd_pr__nfet_01v8__keta_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_57=0.030486
+  sky130_fd_pr__nfet_01v8__ua_diff_57=6.22602e-11
+  sky130_fd_pr__nfet_01v8__ub_diff_57=1.46466e-19
+  sky130_fd_pr__nfet_01v8__eta0_diff_57=2.87515e-6
+  sky130_fd_pr__nfet_01v8__tvoff_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_57=-49294.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_57=-4.14197e-5
+  sky130_fd_pr__nfet_01v8__vth0_diff_57=-0.14144
+  sky130_fd_pr__nfet_01v8__b0_diff_57=1.87189e-7
*
* sky130_fd_pr__nfet_01v8, Bin 058, W = 0.61, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__b0_diff_58=1.38166e-7
+  sky130_fd_pr__nfet_01v8__pdits_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_58=5.06931e-9
+  sky130_fd_pr__nfet_01v8__voff_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_58=-7.0636e-5
+  sky130_fd_pr__nfet_01v8__u0_diff_58=0.0016663
+  sky130_fd_pr__nfet_01v8__nfactor_diff_58=0.47711421
+  sky130_fd_pr__nfet_01v8__keta_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_58=0.03038
+  sky130_fd_pr__nfet_01v8__ua_diff_58=5.13586e-11
+  sky130_fd_pr__nfet_01v8__ub_diff_58=1.96251e-19
+  sky130_fd_pr__nfet_01v8__eta0_diff_58=2.50164e-6
+  sky130_fd_pr__nfet_01v8__tvoff_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_58=-49772.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_58=-3.60388e-5
+  sky130_fd_pr__nfet_01v8__vth0_diff_58=-0.14016
*
* sky130_fd_pr__nfet_01v8, Bin 059, W = 0.65, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__kt1_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_59=-42486.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_59=-0.13818
+  sky130_fd_pr__nfet_01v8__b0_diff_59=3.66155e-8
+  sky130_fd_pr__nfet_01v8__pdits_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_59=-5.23278e-11
+  sky130_fd_pr__nfet_01v8__voff_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_59=8.25295e-5
+  sky130_fd_pr__nfet_01v8__u0_diff_59=0.0016984
+  sky130_fd_pr__nfet_01v8__nfactor_diff_59=0.45856873
+  sky130_fd_pr__nfet_01v8__keta_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_59=0.0299
+  sky130_fd_pr__nfet_01v8__ua_diff_59=2.10287e-11
+  sky130_fd_pr__nfet_01v8__ub_diff_59=3.16657e-19
+  sky130_fd_pr__nfet_01v8__eta0_diff_59=-4.84694e-17
+  sky130_fd_pr__nfet_01v8__tvoff_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_59=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 060, W = 0.65, L = 0.18
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__vsat_diff_60=-41425.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_60=-0.095911
+  sky130_fd_pr__nfet_01v8__pdits_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_60=3.66155e-8
+  sky130_fd_pr__nfet_01v8__voff_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_60=-5.23278e-11
+  sky130_fd_pr__nfet_01v8__pditsd_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_60=8.25291e-5
+  sky130_fd_pr__nfet_01v8__u0_diff_60=0.00078095
+  sky130_fd_pr__nfet_01v8__nfactor_diff_60=0.45856873
+  sky130_fd_pr__nfet_01v8__keta_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_60=0.012547
+  sky130_fd_pr__nfet_01v8__ua_diff_60=2.10287e-11
+  sky130_fd_pr__nfet_01v8__ub_diff_60=3.16657e-19
+  sky130_fd_pr__nfet_01v8__eta0_diff_60=-2.39546e-11
+  sky130_fd_pr__nfet_01v8__tvoff_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_60=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 061, W = 0.65, L = 0.25
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__tvoff_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_61=-37582.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_61=-0.047403
+  sky130_fd_pr__nfet_01v8__pdits_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_61=0.0030431
+  sky130_fd_pr__nfet_01v8__nfactor_diff_61=0.4633
+  sky130_fd_pr__nfet_01v8__keta_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_61=0.0058357
+  sky130_fd_pr__nfet_01v8__ua_diff_61=-9.108e-12
+  sky130_fd_pr__nfet_01v8__ub_diff_61=4.60449e-19
+  sky130_fd_pr__nfet_01v8__eta0_diff_61=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 062, W = 0.65, L = 0.5
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__tvoff_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_62=-49521.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_62=-0.037598
+  sky130_fd_pr__nfet_01v8__pdits_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_62=5.45502e-17
+  sky130_fd_pr__nfet_01v8__b1_diff_62=-2.18149e-18
+  sky130_fd_pr__nfet_01v8__voff_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_62=0.0014459
+  sky130_fd_pr__nfet_01v8__nfactor_diff_62=0.0317
+  sky130_fd_pr__nfet_01v8__keta_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_62=-0.0023861
+  sky130_fd_pr__nfet_01v8__ua_diff_62=2.9602e-12
+  sky130_fd_pr__nfet_01v8__ub_diff_62=2.5142e-19
+  sky130_fd_pr__nfet_01v8__eta0_diff_62=0.0
.include "sky130_fd_pr__nfet_01v8__sf.pm3.spice"
