* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param sky130_fd_pr__nfet_01v8__vth0_correldiff=0.0168
* Number of bins: 63
.param
+  sky130_fd_pr__nfet_01v8__toxe_mult=1.0
+  sky130_fd_pr__nfet_01v8__rshn_mult=1.0
+  sky130_fd_pr__nfet_01v8__overlap_mult=0.9642
+  sky130_fd_pr__nfet_01v8__lint_diff=0.0
+  sky130_fd_pr__nfet_01v8__wint_diff=0.0
+  sky130_fd_pr__nfet_01v8__dlc_diff=-.61492e-9
+  sky130_fd_pr__nfet_01v8__dwc_diff=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 000, W = 1.26, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__voff_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_0=-1.1675e-19
+  sky130_fd_pr__nfet_01v8__pditsd_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_0=1.3935e-11
+  sky130_fd_pr__nfet_01v8__vsat_diff_0=594.41
+  sky130_fd_pr__nfet_01v8__tvoff_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_0=0.0031843
+  sky130_fd_pr__nfet_01v8__vth0_diff_0=' -0.024441 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__nfactor_diff_0=0.37668
+  sky130_fd_pr__nfet_01v8__u0_diff_0=-0.0034894
+  sky130_fd_pr__nfet_01v8__eta0_diff_0=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_0=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 001, W = 1.68, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__eta0_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_1=-1.6979e-19
+  sky130_fd_pr__nfet_01v8__pditsd_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_1=1.0381e-11
+  sky130_fd_pr__nfet_01v8__vsat_diff_1=249.83
+  sky130_fd_pr__nfet_01v8__tvoff_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_1=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_1=0.0047171
+  sky130_fd_pr__nfet_01v8__vth0_diff_1=' 0.0064909 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__nfactor_diff_1=0.31936
+  sky130_fd_pr__nfet_01v8__u0_diff_1=-0.002698
*
* sky130_fd_pr__nfet_01v8, Bin 002, W = 1.0, L = 1.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__nfactor_diff_2=1.11
+  sky130_fd_pr__nfet_01v8__u0_diff_2=-9.2293e-5
+  sky130_fd_pr__nfet_01v8__vth0_diff_2=' 0.0065633 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__eta0_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_2=1.6548e-19
+  sky130_fd_pr__nfet_01v8__kt1_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_2=4.5462e-13
+  sky130_fd_pr__nfet_01v8__vsat_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_2=-0.052872
+  sky130_fd_pr__nfet_01v8__a0_diff_2=0.23412
+  sky130_fd_pr__nfet_01v8__b0_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_2=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_2=-0.0066238
*
* sky130_fd_pr__nfet_01v8, Bin 003, W = 1.0, L = 2.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__keta_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_3=-0.0052707
+  sky130_fd_pr__nfet_01v8__nfactor_diff_3=0.81272
+  sky130_fd_pr__nfet_01v8__u0_diff_3=-0.00043394
+  sky130_fd_pr__nfet_01v8__vth0_diff_3=' -0.0016362 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__eta0_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_3=9.8355e-20
+  sky130_fd_pr__nfet_01v8__kt1_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_3=5.2286e-13
+  sky130_fd_pr__nfet_01v8__vsat_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_3=-0.0086458
+  sky130_fd_pr__nfet_01v8__a0_diff_3=0.030693
+  sky130_fd_pr__nfet_01v8__b0_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_3=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_3=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 004, W = 1.0, L = 4.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__pdits_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_4=0.004486
+  sky130_fd_pr__nfet_01v8__nfactor_diff_4=1.0914
+  sky130_fd_pr__nfet_01v8__u0_diff_4=-0.0017527
+  sky130_fd_pr__nfet_01v8__vth0_diff_4=' -0.0082831 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__eta0_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_4=-1.6247e-20
+  sky130_fd_pr__nfet_01v8__kt1_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_4=4.1897e-12
+  sky130_fd_pr__nfet_01v8__vsat_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_4=-0.011391
+  sky130_fd_pr__nfet_01v8__a0_diff_4=0.034396
+  sky130_fd_pr__nfet_01v8__b0_diff_4=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_4=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 005, W = 1.0, L = 8.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__pdits_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_5=0.0066435
+  sky130_fd_pr__nfet_01v8__nfactor_diff_5=1.1205
+  sky130_fd_pr__nfet_01v8__u0_diff_5=-0.002135
+  sky130_fd_pr__nfet_01v8__vth0_diff_5=' -0.0094295 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__eta0_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_5=-2.1979e-20
+  sky130_fd_pr__nfet_01v8__kt1_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_5=5.0336e-12
+  sky130_fd_pr__nfet_01v8__vsat_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_5=-0.018373
+  sky130_fd_pr__nfet_01v8__a0_diff_5=0.043822
+  sky130_fd_pr__nfet_01v8__b0_diff_5=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_5=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 006, W = 1.0, L = 0.15
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__pclm_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_6=0.0010401
+  sky130_fd_pr__nfet_01v8__nfactor_diff_6=0.85366
+  sky130_fd_pr__nfet_01v8__u0_diff_6=-0.0039089
+  sky130_fd_pr__nfet_01v8__vth0_diff_6=' -0.0015129 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__eta0_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_6=-3.443e-19
+  sky130_fd_pr__nfet_01v8__kt1_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_6=1.4919e-11
+  sky130_fd_pr__nfet_01v8__vsat_diff_6=-2391.8
+  sky130_fd_pr__nfet_01v8__tvoff_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_6=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_6=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 007, W = 1.0, L = 0.18
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__tvoff_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_7=0.0026665
+  sky130_fd_pr__nfet_01v8__nfactor_diff_7=0.063918
+  sky130_fd_pr__nfet_01v8__u0_diff_7=-0.0037374
+  sky130_fd_pr__nfet_01v8__vth0_diff_7=' -0.012203 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__eta0_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_7=-2.5113e-19
+  sky130_fd_pr__nfet_01v8__kt1_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_7=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_7=1.4741e-11
+  sky130_fd_pr__nfet_01v8__vsat_diff_7=-5172.6
+  sky130_fd_pr__nfet_01v8__a0_diff_7=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 008, W = 1.0, L = 0.25
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__a0_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_8=1.9388e-11
+  sky130_fd_pr__nfet_01v8__tvoff_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_8=0.00033191
+  sky130_fd_pr__nfet_01v8__nfactor_diff_8=1.1053
+  sky130_fd_pr__nfet_01v8__u0_diff_8=-0.0052052
+  sky130_fd_pr__nfet_01v8__vth0_diff_8=' -0.010036 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__eta0_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_8=-7.5909e-20
+  sky130_fd_pr__nfet_01v8__kt1_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_8=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_8=-13673.0
*
* sky130_fd_pr__nfet_01v8, Bin 009, W = 1.0, L = 0.5
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__kt1_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_9=-1.1801e-19
+  sky130_fd_pr__nfet_01v8__vsat_diff_9=-6758.5
+  sky130_fd_pr__nfet_01v8__a0_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_9=6.0594e-12
+  sky130_fd_pr__nfet_01v8__tvoff_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_9=0.0048538
+  sky130_fd_pr__nfet_01v8__nfactor_diff_9=1.4173
+  sky130_fd_pr__nfet_01v8__u0_diff_9=-0.0025986
+  sky130_fd_pr__nfet_01v8__vth0_diff_9=' 0.001985 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__eta0_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_9=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_9=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 010, W = 2.0, L = 0.15
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__ags_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_10=0.0036033
+  sky130_fd_pr__nfet_01v8__ua_diff_10=6.5387e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_10=-1.6773e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_10=-3162.6
+  sky130_fd_pr__nfet_01v8__kt1_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_10=' 0.004973 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__pdits_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_10=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_10=0.58499
+  sky130_fd_pr__nfet_01v8__u0_diff_10=-0.0017828
*
* sky130_fd_pr__nfet_01v8, Bin 011, W = 3.0, L = 1.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__pclm_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_11=0.9632
+  sky130_fd_pr__nfet_01v8__u0_diff_11=-0.00030771
+  sky130_fd_pr__nfet_01v8__ags_diff_11=-0.029026
+  sky130_fd_pr__nfet_01v8__keta_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_11=-0.0031799
+  sky130_fd_pr__nfet_01v8__ua_diff_11=3.5948e-14
+  sky130_fd_pr__nfet_01v8__eta0_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_11=6.1194e-20
+  sky130_fd_pr__nfet_01v8__tvoff_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_11=0.016472
+  sky130_fd_pr__nfet_01v8__rdsw_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_11=' 0.0058576 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__pdits_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_11=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_11=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 012, W = 3.0, L = 2.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__pditsd_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_12=1.0173
+  sky130_fd_pr__nfet_01v8__u0_diff_12=-0.0031613
+  sky130_fd_pr__nfet_01v8__ags_diff_12=-0.037956
+  sky130_fd_pr__nfet_01v8__keta_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_12=0.003257
+  sky130_fd_pr__nfet_01v8__ua_diff_12=8.1792e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_12=-2.2603e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_12=0.044769
+  sky130_fd_pr__nfet_01v8__rdsw_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_12=' -0.010873 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__pdits_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_12=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_12=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 013, W = 3.0, L = 4.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__pdits_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_13=0.98167
+  sky130_fd_pr__nfet_01v8__u0_diff_13=-0.0031709
+  sky130_fd_pr__nfet_01v8__ags_diff_13=-0.0017409
+  sky130_fd_pr__nfet_01v8__keta_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_13=0.0033393
+  sky130_fd_pr__nfet_01v8__ua_diff_13=8.1683e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_13=-2.1077e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_13=0.021688
+  sky130_fd_pr__nfet_01v8__rdsw_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_13=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_13=' -0.0074909 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__b0_diff_13=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 014, W = 3.0, L = 8.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__b0_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_14=0.91425
+  sky130_fd_pr__nfet_01v8__u0_diff_14=-0.0024205
+  sky130_fd_pr__nfet_01v8__ags_diff_14=-0.022734
+  sky130_fd_pr__nfet_01v8__keta_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_14=0.0045599
+  sky130_fd_pr__nfet_01v8__ua_diff_14=5.8682e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_14=-1.7238e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_14=0.04225
+  sky130_fd_pr__nfet_01v8__rdsw_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_14=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_14=' -0.0073982 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
*
* sky130_fd_pr__nfet_01v8, Bin 015, W = 3.0, L = 0.15
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__kt1_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_15=-647.87
+  sky130_fd_pr__nfet_01v8__vth0_diff_15=' -0.018099 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__b0_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_15=1.0234
+  sky130_fd_pr__nfet_01v8__u0_diff_15=-0.0038701
+  sky130_fd_pr__nfet_01v8__ags_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_15=0.010464
+  sky130_fd_pr__nfet_01v8__ua_diff_15=1.3818e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_15=-3.6525e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_15=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_15=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 016, W = 3.0, L = 0.18
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__a0_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_16=-1586.1
+  sky130_fd_pr__nfet_01v8__vth0_diff_16=' -0.0039193 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__b0_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_16=0.63266
+  sky130_fd_pr__nfet_01v8__u0_diff_16=-0.0019616
+  sky130_fd_pr__nfet_01v8__ags_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_16=0.0098403
+  sky130_fd_pr__nfet_01v8__ua_diff_16=7.4303e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_16=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_16=-3.9342e-20
+  sky130_fd_pr__nfet_01v8__tvoff_diff_16=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 017, W = 3.0, L = 0.25
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__tvoff_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_17=-3384.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_17=' -0.018442 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__pdits_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_17=1.3587
+  sky130_fd_pr__nfet_01v8__u0_diff_17=-0.0013448
+  sky130_fd_pr__nfet_01v8__ags_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_17=0.0072332
+  sky130_fd_pr__nfet_01v8__ua_diff_17=3.3377e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_17=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_17=8.1803e-20
*
* sky130_fd_pr__nfet_01v8, Bin 018, W = 3.0, L = 0.5
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__ub_diff_18=5.989e-20
+  sky130_fd_pr__nfet_01v8__tvoff_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_18=2230.3
+  sky130_fd_pr__nfet_01v8__vth0_diff_18=' -0.0085702 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__pdits_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_18=0.98656
+  sky130_fd_pr__nfet_01v8__u0_diff_18=-0.0010556
+  sky130_fd_pr__nfet_01v8__ags_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_18=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_18=0.0032531
+  sky130_fd_pr__nfet_01v8__ua_diff_18=2.2684e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_18=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 019, W = 5.0, L = 1.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__eta0_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_19=4.4209e-13
+  sky130_fd_pr__nfet_01v8__ub_diff_19=8.0805e-20
+  sky130_fd_pr__nfet_01v8__tvoff_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_19=0.013728
+  sky130_fd_pr__nfet_01v8__rdsw_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_19=' 0.0022292 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__pdits_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_19=0.91555
+  sky130_fd_pr__nfet_01v8__u0_diff_19=-0.00035451
+  sky130_fd_pr__nfet_01v8__ags_diff_19=0.0044706
+  sky130_fd_pr__nfet_01v8__keta_diff_19=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_19=0.0051373
*
* sky130_fd_pr__nfet_01v8, Bin 020, W = 5.0, L = 2.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__ua_diff_20=1.2021e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_20=-3.4149e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_20=0.039045
+  sky130_fd_pr__nfet_01v8__rdsw_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_20=' -0.013628 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__pdits_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_20=0.98704
+  sky130_fd_pr__nfet_01v8__u0_diff_20=-0.0042881
+  sky130_fd_pr__nfet_01v8__ags_diff_20=-0.016925
+  sky130_fd_pr__nfet_01v8__keta_diff_20=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_20=0.0035839
*
* sky130_fd_pr__nfet_01v8, Bin 021, W = 5.0, L = 4.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__ags_diff_21=-0.047476
+  sky130_fd_pr__nfet_01v8__keta_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_21=0.0031859
+  sky130_fd_pr__nfet_01v8__ua_diff_21=7.4952e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_21=-2.4257e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_21=0.065845
+  sky130_fd_pr__nfet_01v8__rdsw_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_21=' -0.011082 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__pdits_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_21=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_21=0.87421
+  sky130_fd_pr__nfet_01v8__u0_diff_21=-0.0028759
*
* sky130_fd_pr__nfet_01v8, Bin 022, W = 5.0, L = 8.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__pclm_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_22=0.91257
+  sky130_fd_pr__nfet_01v8__u0_diff_22=-0.0016954
+  sky130_fd_pr__nfet_01v8__ags_diff_22=0.0065854
+  sky130_fd_pr__nfet_01v8__keta_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_22=0.0050836
+  sky130_fd_pr__nfet_01v8__ua_diff_22=4.0804e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_22=-8.907e-20
+  sky130_fd_pr__nfet_01v8__tvoff_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_22=0.0086619
+  sky130_fd_pr__nfet_01v8__rdsw_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_22=' -0.0040453 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__pdits_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_22=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_22=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 023, W = 5.0, L = 0.15
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__pditsd_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_23=1.3757
+  sky130_fd_pr__nfet_01v8__u0_diff_23=3.9678e-6
+  sky130_fd_pr__nfet_01v8__ags_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_23=0.0034222
+  sky130_fd_pr__nfet_01v8__ua_diff_23=-6.8599e-13
+  sky130_fd_pr__nfet_01v8__eta0_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_23=5.4464e-20
+  sky130_fd_pr__nfet_01v8__tvoff_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_23=4444.9
+  sky130_fd_pr__nfet_01v8__kt1_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_23=' -0.0038779 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__pdits_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_23=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_23=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 024, W = 5.0, L = 0.18
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__pdits_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_24=1.6087
+  sky130_fd_pr__nfet_01v8__u0_diff_24=-0.0073288
+  sky130_fd_pr__nfet_01v8__ags_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_24=0.0088478
+  sky130_fd_pr__nfet_01v8__ua_diff_24=2.5229e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_24=-4.484e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_24=-1451.2
+  sky130_fd_pr__nfet_01v8__kt1_diff_24=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_24=' -0.021745 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__b0_diff_24=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 025, W = 5.0, L = 0.25
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__b0_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_25=1.1914
+  sky130_fd_pr__nfet_01v8__u0_diff_25=-0.0010782
+  sky130_fd_pr__nfet_01v8__ags_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_25=0.0056373
+  sky130_fd_pr__nfet_01v8__ua_diff_25=2.7261e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_25=1.3675e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_25=-3533.5
+  sky130_fd_pr__nfet_01v8__kt1_diff_25=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_25=' -0.0035273 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
*
* sky130_fd_pr__nfet_01v8, Bin 026, W = 5.0, L = 0.5
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__kt1_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_26=-3043.1
+  sky130_fd_pr__nfet_01v8__vth0_diff_26=' -0.0034318 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__b0_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_26=1.1397
+  sky130_fd_pr__nfet_01v8__u0_diff_26=-0.00035449
+  sky130_fd_pr__nfet_01v8__ags_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_26=0.0023237
+  sky130_fd_pr__nfet_01v8__ua_diff_26=-1.4727e-13
+  sky130_fd_pr__nfet_01v8__eta0_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_26=3.1599e-20
+  sky130_fd_pr__nfet_01v8__tvoff_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_26=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_26=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 027, W = 7.0, L = 1.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__a0_diff_27=0.066133
+  sky130_fd_pr__nfet_01v8__rdsw_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_27=' -0.013324 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__b0_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_27=0.97611
+  sky130_fd_pr__nfet_01v8__u0_diff_27=-0.0014921
+  sky130_fd_pr__nfet_01v8__ags_diff_27=-0.056372
+  sky130_fd_pr__nfet_01v8__keta_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_27=0.0031651
+  sky130_fd_pr__nfet_01v8__ua_diff_27=4.6745e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_27=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_27=-1.0031e-20
+  sky130_fd_pr__nfet_01v8__tvoff_diff_27=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 028, W = 7.0, L = 2.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__tvoff_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_28=0.040647
+  sky130_fd_pr__nfet_01v8__rdsw_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_28=' -0.0068792 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__pdits_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_28=0.95569
+  sky130_fd_pr__nfet_01v8__u0_diff_28=-0.0017647
+  sky130_fd_pr__nfet_01v8__ags_diff_28=-0.024329
+  sky130_fd_pr__nfet_01v8__keta_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_28=0.0043246
+  sky130_fd_pr__nfet_01v8__ua_diff_28=4.7856e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_28=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_28=-7.3548e-20
*
* sky130_fd_pr__nfet_01v8, Bin 029, W = 7.0, L = 4.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__ub_diff_29=-4.1864e-20
+  sky130_fd_pr__nfet_01v8__tvoff_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_29=-0.021276
+  sky130_fd_pr__nfet_01v8__rdsw_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_29=' -0.0095112 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__pdits_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_29=0.87453
+  sky130_fd_pr__nfet_01v8__u0_diff_29=-0.0014569
+  sky130_fd_pr__nfet_01v8__ags_diff_29=0.022917
+  sky130_fd_pr__nfet_01v8__keta_diff_29=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_29=0.0026623
+  sky130_fd_pr__nfet_01v8__ua_diff_29=3.7953e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_29=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 030, W = 7.0, L = 8.0
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__eta0_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_30=-6.3508e-20
+  sky130_fd_pr__nfet_01v8__tvoff_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_30=0.014619
+  sky130_fd_pr__nfet_01v8__rdsw_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_30=' -0.0023907 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__pdits_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_30=0.83331
+  sky130_fd_pr__nfet_01v8__u0_diff_30=-0.0012126
+  sky130_fd_pr__nfet_01v8__ags_diff_30=-0.0001807
+  sky130_fd_pr__nfet_01v8__keta_diff_30=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_30=0.0043065
+  sky130_fd_pr__nfet_01v8__ua_diff_30=2.9064e-12
*
* sky130_fd_pr__nfet_01v8, Bin 031, W = 7.0, L = 0.15
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__ua_diff_31=-6.1562e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_31=2.6424e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_31=5596.7
+  sky130_fd_pr__nfet_01v8__kt1_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_31=' 0.0036689 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__pdits_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_31=-0.54209
+  sky130_fd_pr__nfet_01v8__u0_diff_31=0.0020466
+  sky130_fd_pr__nfet_01v8__ags_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_31=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_31=-0.0021477
*
* sky130_fd_pr__nfet_01v8, Bin 032, W = 7.0, L = 0.18
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__ags_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_32=0.0071845
+  sky130_fd_pr__nfet_01v8__ua_diff_32=2.0407e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_32=-3.0535e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_32=-360.04
+  sky130_fd_pr__nfet_01v8__kt1_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_32=' -0.019564 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__pdits_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_32=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_32=1.5101
+  sky130_fd_pr__nfet_01v8__u0_diff_32=-0.0057978
*
* sky130_fd_pr__nfet_01v8, Bin 033, W = 7.0, L = 0.25
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__pclm_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_33=1.0177
+  sky130_fd_pr__nfet_01v8__u0_diff_33=-0.0012465
+  sky130_fd_pr__nfet_01v8__ags_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_33=0.0060444
+  sky130_fd_pr__nfet_01v8__ua_diff_33=3.6045e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_33=9.6789e-20
+  sky130_fd_pr__nfet_01v8__tvoff_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_33=-3883.6
+  sky130_fd_pr__nfet_01v8__kt1_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_33=' -0.0060464 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__pdits_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_33=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_33=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 034, W = 7.0, L = 0.5
* ---------------------------------
+  sky130_fd_pr__nfet_01v8__pditsd_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_34=1.0862
+  sky130_fd_pr__nfet_01v8__u0_diff_34=-0.0003721
+  sky130_fd_pr__nfet_01v8__ags_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_34=0.0018509
+  sky130_fd_pr__nfet_01v8__ua_diff_34=3.6306e-15
+  sky130_fd_pr__nfet_01v8__eta0_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_34=2.1029e-20
+  sky130_fd_pr__nfet_01v8__tvoff_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_34=-1504.3
+  sky130_fd_pr__nfet_01v8__kt1_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_34=' -0.0060299 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__pdits_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_34=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_34=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 035, W = 0.42, L = 1.0
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__pdits_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_35=4.952e-9
+  sky130_fd_pr__nfet_01v8__pditsd_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_35=1.7654
+  sky130_fd_pr__nfet_01v8__u0_diff_35=-0.0051179
+  sky130_fd_pr__nfet_01v8__ags_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_35=0.0017141
+  sky130_fd_pr__nfet_01v8__ua_diff_35=1.4292e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_35=-1.067e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_35=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_35=' -0.010841 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__b0_diff_35=-1.4147e-7
*
* sky130_fd_pr__nfet_01v8, Bin 036, W = 0.42, L = 20.0
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__b0_diff_36=2.3328e-8
+  sky130_fd_pr__nfet_01v8__pdits_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_36=3.9114e-9
+  sky130_fd_pr__nfet_01v8__pditsd_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_36=1.5453
+  sky130_fd_pr__nfet_01v8__u0_diff_36=-0.0036019
+  sky130_fd_pr__nfet_01v8__ags_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_36=0.0051159
+  sky130_fd_pr__nfet_01v8__ua_diff_36=7.4306e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_36=-1.172e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_36=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_36=' -0.0082177 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
*
* sky130_fd_pr__nfet_01v8, Bin 037, W = 0.42, L = 2.0
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__kt1_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_37=' -0.039645 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__b0_diff_37=4.2553e-8
+  sky130_fd_pr__nfet_01v8__pdits_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_37=8.1602e-9
+  sky130_fd_pr__nfet_01v8__pditsd_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_37=1.4271
+  sky130_fd_pr__nfet_01v8__u0_diff_37=-0.0061353
+  sky130_fd_pr__nfet_01v8__ags_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_37=0.004022
+  sky130_fd_pr__nfet_01v8__ua_diff_37=1.7334e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_37=-2.4886e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_37=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_37=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 038, W = 0.42, L = 4.0
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__a0_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_38=' -0.02604 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__b0_diff_38=4.0509e-9
+  sky130_fd_pr__nfet_01v8__pdits_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_38=5.7829e-9
+  sky130_fd_pr__nfet_01v8__pditsd_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_38=1.2119
+  sky130_fd_pr__nfet_01v8__u0_diff_38=-0.0039583
+  sky130_fd_pr__nfet_01v8__ags_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_38=0.008427
+  sky130_fd_pr__nfet_01v8__ua_diff_38=1.0335e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_38=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_38=-1.0155e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_38=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 039, W = 0.42, L = 8.0
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__tvoff_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_39=' -0.0044661 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__pdits_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_39=3.9409e-8
+  sky130_fd_pr__nfet_01v8__b1_diff_39=3.4348e-9
+  sky130_fd_pr__nfet_01v8__pditsd_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_39=1.2957
+  sky130_fd_pr__nfet_01v8__u0_diff_39=-0.0037655
+  sky130_fd_pr__nfet_01v8__ags_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_39=-0.00018284
+  sky130_fd_pr__nfet_01v8__ua_diff_39=8.7608e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_39=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_39=-1.6334e-19
*
* sky130_fd_pr__nfet_01v8, Bin 040, W = 0.42, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__tvoff_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_40=-10.537
+  sky130_fd_pr__nfet_01v8__kt1_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_40=' -0.021136 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__pdits_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_40=0.72905
+  sky130_fd_pr__nfet_01v8__u0_diff_40=0.0019295
+  sky130_fd_pr__nfet_01v8__ags_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_40=0.0019759
+  sky130_fd_pr__nfet_01v8__ua_diff_40=-6.3825e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_40=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_40=6.55e-19
*
* sky130_fd_pr__nfet_01v8, Bin 041, W = 0.42, L = 0.18
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__eta0_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_41=-2.2736e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_41=-14544.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_41=' -0.039339 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__pdits_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_41=0.1923
+  sky130_fd_pr__nfet_01v8__u0_diff_41=-0.0066627
+  sky130_fd_pr__nfet_01v8__ags_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_41=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_41=-0.0033684
+  sky130_fd_pr__nfet_01v8__ua_diff_41=2.7564e-11
*
* sky130_fd_pr__nfet_01v8, Bin 042, W = 0.42, L = 0.5
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__ua_diff_42=1.5471e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_42=-1.3038e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_42=-14884.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_42=' -0.011611 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__pdits_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_42=1.7635
+  sky130_fd_pr__nfet_01v8__u0_diff_42=-0.005084
+  sky130_fd_pr__nfet_01v8__ags_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_42=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_42=0.010251
*
* sky130_fd_pr__nfet_01v8, Bin 043, W = 0.55, L = 1.0
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__ags_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_43=0.0063157
+  sky130_fd_pr__nfet_01v8__ua_diff_43=5.5055e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_43=5.3284e-20
+  sky130_fd_pr__nfet_01v8__tvoff_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_43=' 0.0027609 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__pdits_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_43=1.1418e-7
+  sky130_fd_pr__nfet_01v8__voff_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_43=2.2032e-9
+  sky130_fd_pr__nfet_01v8__pditsd_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_43=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_43=1.4822
+  sky130_fd_pr__nfet_01v8__u0_diff_43=-0.0023728
*
* sky130_fd_pr__nfet_01v8, Bin 044, W = 0.55, L = 2.0
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__pclm_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_44=1.4443
+  sky130_fd_pr__nfet_01v8__u0_diff_44=-0.0075566
+  sky130_fd_pr__nfet_01v8__ags_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_44=0.0055983
+  sky130_fd_pr__nfet_01v8__ua_diff_44=2.0025e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_44=-4.8209e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_44=' -0.022111 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__pdits_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_44=6.6128e-8
+  sky130_fd_pr__nfet_01v8__voff_diff_44=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_44=8.0499e-9
+  sky130_fd_pr__nfet_01v8__pditsd_diff_44=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 045, W = 0.55, L = 4.0
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__pditsd_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_45=1.116
+  sky130_fd_pr__nfet_01v8__u0_diff_45=-0.0043212
+  sky130_fd_pr__nfet_01v8__ags_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_45=0.0030788
+  sky130_fd_pr__nfet_01v8__ua_diff_45=1.1458e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_45=-1.9509e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_45=' -0.0093871 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__pdits_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_45=3.319e-8
+  sky130_fd_pr__nfet_01v8__voff_diff_45=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_45=3.3437e-9
*
* sky130_fd_pr__nfet_01v8, Bin 046, W = 0.55, L = 8.0
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__pdits_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_46=1.9669e-9
+  sky130_fd_pr__nfet_01v8__pditsd_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_46=1.063
+  sky130_fd_pr__nfet_01v8__u0_diff_46=-0.0026409
+  sky130_fd_pr__nfet_01v8__ags_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_46=0.0037614
+  sky130_fd_pr__nfet_01v8__ua_diff_46=6.4629e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_46=-7.4503e-22
+  sky130_fd_pr__nfet_01v8__tvoff_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_46=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_46=' -0.0024093 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__b0_diff_46=2.1974e-8
*
* sky130_fd_pr__nfet_01v8, Bin 047, W = 0.55, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__b0_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_47=0.63538
+  sky130_fd_pr__nfet_01v8__u0_diff_47=-0.0041087
+  sky130_fd_pr__nfet_01v8__ags_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_47=0.0015007
+  sky130_fd_pr__nfet_01v8__ua_diff_47=1.6315e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_47=-6.6985e-20
+  sky130_fd_pr__nfet_01v8__tvoff_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_47=-1436.9
+  sky130_fd_pr__nfet_01v8__kt1_diff_47=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_47=' -0.02218 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
*
* sky130_fd_pr__nfet_01v8, Bin 048, W = 0.55, L = 0.5
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__kt1_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_48=-12346.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_48=' -0.010226 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__b0_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_48=1.6569
+  sky130_fd_pr__nfet_01v8__u0_diff_48=-0.0021061
+  sky130_fd_pr__nfet_01v8__ags_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_48=0.0022728
+  sky130_fd_pr__nfet_01v8__ua_diff_48=3.9332e-12
+  sky130_fd_pr__nfet_01v8__eta0_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_48=-3.7598e-21
+  sky130_fd_pr__nfet_01v8__tvoff_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_48=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_48=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 049, W = 0.64, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__a0_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_49=2643.3
+  sky130_fd_pr__nfet_01v8__vth0_diff_49=' 0.011361 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__b0_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_49=0.46974
+  sky130_fd_pr__nfet_01v8__u0_diff_49=-0.0029103
+  sky130_fd_pr__nfet_01v8__ags_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_49=0.0040992
+  sky130_fd_pr__nfet_01v8__ua_diff_49=1.1487e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_49=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_49=-1.3093e-19
+  sky130_fd_pr__nfet_01v8__tvoff_diff_49=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 050, W = 0.84, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__tvoff_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_50=5763.7
+  sky130_fd_pr__nfet_01v8__kt1_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_50=' -0.017481 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__pdits_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_50=0.31729
+  sky130_fd_pr__nfet_01v8__u0_diff_50=-0.0027183
+  sky130_fd_pr__nfet_01v8__ags_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_50=0.00076174
+  sky130_fd_pr__nfet_01v8__ua_diff_50=1.0629e-11
+  sky130_fd_pr__nfet_01v8__eta0_diff_50=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_50=-4.8113e-21
*
* sky130_fd_pr__nfet_01v8, Bin 051, W = 0.74, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__tvoff_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_51=' 0.0 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__pdits_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_51=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_51=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 052, W = 0.36, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__ub_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_52=-2546.2
+  sky130_fd_pr__nfet_01v8__kt1_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_52=' 0.042004 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__pdits_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_52=-0.0031323
+  sky130_fd_pr__nfet_01v8__nfactor_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_52=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_52=0.011633
+  sky130_fd_pr__nfet_01v8__ua_diff_52=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 053, W = 0.39, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__ua_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_53=-1950.4
+  sky130_fd_pr__nfet_01v8__kt1_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_53=' 0.032109 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__pdits_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_53=-0.0029036
+  sky130_fd_pr__nfet_01v8__nfactor_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_53=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_53=0.0090649
*
* sky130_fd_pr__nfet_01v8, Bin 054, W = 0.52, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__keta_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_54=' 0.0 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__pdits_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_54=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_54=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 055, W = 0.54, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__pclm_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_55=' 0.0 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__pdits_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_55=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_55=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 056, W = 0.58, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__pditsd_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_56=' 0.0 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__pdits_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_56=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_56=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 057, W = 0.6, L = 0.15
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__pdits_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_57=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_57=' 0.0 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__b0_diff_57=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 058, W = 0.61, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__b0_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_58=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_58=' 0.0 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
*
* sky130_fd_pr__nfet_01v8, Bin 059, W = 0.65, L = 0.15
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__kt1_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_59=' 0.0 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__b0_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__pdits_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_59=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_59=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 060, W = 0.65, L = 0.18
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__vsat_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_60=' 0.0 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__pdits_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__tvoff_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_60=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_60=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 061, W = 0.65, L = 0.25
* -----------------------------------
+  sky130_fd_pr__nfet_01v8__tvoff_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_61=' 0.0 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__pdits_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_61=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_61=0.0
*
* sky130_fd_pr__nfet_01v8, Bin 062, W = 0.65, L = 0.5
* ----------------------------------
+  sky130_fd_pr__nfet_01v8__tvoff_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__rdsw_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__a0_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__vsat_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__kt1_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__vth0_diff_62=' 0.0 + sky130_fd_pr__nfet_01v8__vth0_correldiff'
+  sky130_fd_pr__nfet_01v8__pdits_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__b0_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__b1_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__voff_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__pditsd_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__pclm_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__u0_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__nfactor_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__keta_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__ags_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__k2_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__ua_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__ub_diff_62=0.0
+  sky130_fd_pr__nfet_01v8__eta0_diff_62=0.0
.include "sky130_fd_pr__nfet_01v8.pm3.spice"
