* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 18
.param
+  sky130_fd_pr__rf_nfet_01v8_lvt_b__toxe_mult=1.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_b__rbpb_mult=1.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_b__overlap_mult=9.2429e-1
+  sky130_fd_pr__rf_nfet_01v8_lvt_b__ajunction_mult=1.0004e+0
+  sky130_fd_pr__rf_nfet_01v8_lvt_b__pjunction_mult=8.9176e-1
+  sky130_fd_pr__rf_nfet_01v8_lvt_b__lint_diff=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_b__wint_diff=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_b__rshg_diff=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_b__dlc_diff=-1.3619e-9
+  sky130_fd_pr__rf_nfet_01v8_lvt_b__dwc_diff=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_b__xgw_diff=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt__aw_cap_mult_p42=1.0
+  sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_dist_mult_p42=1.0
+  sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_stub_mult_p42=1.0
+  sky130_fd_pr__rf_nfet_01v8_lvt__aw_cap_mult=1.0
+  sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_dist_mult=1.0
+  sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_stub_mult=1.0
+  sky130_fd_pr__rf_nfet_01v8_lvt__aw_rd_mult=1.0
+  sky130_fd_pr__rf_nfet_01v8_lvt__aw_rs_mult=1.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 000, W = 1.65, L = 0.15
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_0=-0.0019098
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ags_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_0=-0.00025989
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_0=-4140.2
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b1_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__voff_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b0_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ub_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ua_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__a0_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__pclm_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__kt1_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__nfactor_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__rdsw_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_0=-0.017838
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 001, W = 1.65, L = 0.18
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__kt1_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__nfactor_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__rdsw_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_1=-0.0088849
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_1=-0.002597
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ags_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_1=0.0006887
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_1=-1709.2
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b1_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__voff_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b0_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ub_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ua_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__a0_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__pclm_diff_1=0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 002, W = 1.65, L = 0.25
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__kt1_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__nfactor_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__rdsw_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_2=-0.0018947
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_2=-0.012344
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ags_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_2=0.00070107
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_2=-3891.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b1_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__voff_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b0_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ub_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ua_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__a0_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__pclm_diff_2=0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 003, W = 3.01, L = 0.15
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__pclm_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__kt1_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__nfactor_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__rdsw_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_3=-0.013074
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_3=-0.011262
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ags_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_3=-0.0041387
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_3=-6088.7
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b1_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__voff_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b0_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ub_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ua_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__a0_diff_3=0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 004, W = 3.01, L = 0.18
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__pclm_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__kt1_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__nfactor_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__rdsw_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_4=-0.008659
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_4=-0.020003
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ags_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_4=-0.0021579
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_4=-1519.6
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b1_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__voff_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b0_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ub_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ua_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__a0_diff_4=0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 005, W = 3.01, L = 0.25
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__a0_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__pclm_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__kt1_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__nfactor_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__rdsw_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_5=-0.0014917
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_5=-0.0074298
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ags_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_5=-0.0010425
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_5=-415.88
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b1_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__voff_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b0_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ub_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ua_diff_5=0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 006, W = 5.05, L = 0.15
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ua_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__a0_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__pclm_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__kt1_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__nfactor_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__rdsw_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_6=-0.020457
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_6=-0.010257
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ags_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_6=-0.008363
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_6=-5555.5
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b1_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__voff_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b0_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ub_diff_6=0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 007, W = 5.05, L = 0.18
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ub_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ua_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__a0_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__pclm_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__kt1_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__nfactor_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__rdsw_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_7=-0.0091424
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_7=-0.01706
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ags_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_7=-0.0042397
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_7=-790.25
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b1_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__voff_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b0_diff_7=0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 008, W = 5.05, L = 0.25
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__voff_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b0_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ub_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ua_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__a0_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__pclm_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__kt1_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__nfactor_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__rdsw_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_8=-0.0013518
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_8=-0.0069456
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ags_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_8=-0.0019193
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_8=-105.44
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b1_diff_8=0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 000, W = 1.65, L = 0.15
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ua_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__pclm_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__nfactor_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__a0_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__voff_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b0_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_0=-0.017526
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_0=-0.0051133
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_0=-0.0060348
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_0=145.4
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__kt1_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b1_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__rdsw_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ags_diff_0=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ub_diff_0=0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 001, W = 1.65, L = 0.18
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ags_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ub_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ua_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__pclm_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__nfactor_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__a0_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__voff_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b0_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_1=-0.0093978
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_1=-0.010042
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_1=-0.0028136
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_1=-1622.4
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__kt1_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b1_diff_1=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__rdsw_diff_1=0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 002, W = 1.65, L = 0.25
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ags_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ub_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ua_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__pclm_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__nfactor_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__a0_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__voff_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b0_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_2=-0.0023374
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_2=-0.017756
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_2=-0.0017253
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_2=2328.3
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__kt1_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b1_diff_2=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__rdsw_diff_2=0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 003, W = 3.01, L = 0.15
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__kt1_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b1_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__rdsw_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ags_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ub_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ua_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__pclm_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__nfactor_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__a0_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__voff_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b0_diff_3=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_3=-0.014282
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_3=-0.0085151
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_3=-0.0046757
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_3=-6719.9
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 004, W = 3.01, L = 0.18
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_4=-0.0069428
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_4=327.64
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__kt1_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b1_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__rdsw_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ags_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ub_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ua_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__pclm_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__nfactor_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__a0_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__voff_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b0_diff_4=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_4=-0.0096416
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_4=-0.017088
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 005, W = 3.01, L = 0.25
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_5=-0.019991
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_5=-0.0042474
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_5=9083.2
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__kt1_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b1_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__rdsw_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ags_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ub_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ua_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__pclm_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__nfactor_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__a0_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__voff_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b0_diff_5=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_5=-0.0027118
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 006, W = 5.05, L = 0.15
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__voff_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b0_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_6=-0.01916
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_6=-0.013021
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_6=-0.0061579
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_6=-6431.2
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__kt1_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b1_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__rdsw_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ags_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ub_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ua_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__pclm_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__nfactor_diff_6=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__a0_diff_6=0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 007, W = 5.05, L = 0.18
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__nfactor_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__a0_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__voff_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b0_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_7=-0.011438
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_7=-0.018674
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_7=-0.0084514
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_7=-2625.5
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__kt1_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b1_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__rdsw_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ags_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ub_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ua_diff_7=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__pclm_diff_7=0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 008, W = 5.05, L = 0.25
* ------------------------------------------------
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__pclm_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__nfactor_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__a0_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__voff_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b0_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_8=-0.0028374
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_8=-0.0065635
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_8=14190.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_8=-0.024019
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__kt1_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b1_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__rdsw_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ags_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ub_diff_8=0.0
+  sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ua_diff_8=0.0
.include "sky130_fd_pr__rf_nfet_01v8_lvt_b.pm3.spice"
