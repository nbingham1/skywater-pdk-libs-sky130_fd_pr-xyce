* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 68
.param
+  sky130_fd_pr__pfet_01v8_hvt__toxe_mult=1.0
+  sky130_fd_pr__pfet_01v8_hvt__rshp_mult=1.0
+  sky130_fd_pr__pfet_01v8_hvt__overlap_mult=1.0
+  sky130_fd_pr__pfet_01v8_hvt__lint_diff=0.0
+  sky130_fd_pr__pfet_01v8_hvt__wint_diff=0.0
+  sky130_fd_pr__pfet_01v8_hvt__dlc_diff=0.0
+  sky130_fd_pr__pfet_01v8_hvt__dwc_diff=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 000, W = 1.26, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_0=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_0=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 001, W = 1.68, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_1=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_1=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 002, W = 1.0, L = 1.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_2=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_2=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 003, W = 1.0, L = 2.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_3=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_3=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 004, W = 1.0, L = 4.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_4=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_4=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 005, W = 1.0, L = 8.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_5=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_5=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 006, W = 1.0, L = 0.15
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_6=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_6=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 007, W = 1.0, L = 0.18
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_7=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_7=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 008, W = 1.0, L = 0.25
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_8=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_8=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 009, W = 1.0, L = 0.5
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_9=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_9=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 010, W = 3.0, L = 1.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_10=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_10=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 011, W = 3.0, L = 2.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_11=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_11=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 012, W = 3.0, L = 4.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_12=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_12=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 013, W = 3.0, L = 8.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_13=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_13=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 014, W = 3.0, L = 0.15
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_14=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_14=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 015, W = 3.0, L = 0.18
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_15=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_15=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 016, W = 3.0, L = 0.25
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_16=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_16=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 017, W = 3.0, L = 0.5
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_17=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_17=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 018, W = 5.0, L = 1.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_18=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_18=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 019, W = 5.0, L = 2.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_19=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_19=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 020, W = 5.0, L = 4.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_20=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_20=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 021, W = 5.0, L = 8.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_21=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_21=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 022, W = 5.0, L = 0.15
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_22=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_22=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 023, W = 5.0, L = 0.18
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_23=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_23=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 024, W = 5.0, L = 0.25
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_24=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_24=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 025, W = 5.0, L = 0.5
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_25=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_25=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 026, W = 7.0, L = 1.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_26=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_26=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 027, W = 7.0, L = 2.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_27=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_27=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 028, W = 7.0, L = 4.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_28=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_28=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 029, W = 7.0, L = 8.0
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_29=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_29=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 030, W = 7.0, L = 0.15
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_30=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_30=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 031, W = 7.0, L = 0.18
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_31=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_31=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 032, W = 7.0, L = 0.25
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_32=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_32=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 033, W = 7.0, L = 0.5
* ----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_33=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_33=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 034, W = 0.42, L = 1.0
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_34=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_34=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 035, W = 0.42, L = 20.0
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_35=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_35=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 036, W = 0.42, L = 2.0
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_36=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_36=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 037, W = 0.42, L = 4.0
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_37=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_37=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 038, W = 0.42, L = 8.0
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_38=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_38=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 039, W = 0.42, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_39=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_39=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 040, W = 0.42, L = 0.18
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_40=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_40=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 041, W = 0.42, L = 0.5
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_41=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_41=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 042, W = 0.55, L = 1.0
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_42=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_42=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 043, W = 0.55, L = 2.0
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_43=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_43=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 044, W = 0.55, L = 4.0
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_44=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_44=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 045, W = 0.55, L = 8.0
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_45=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_45=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 046, W = 0.55, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_46=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_46=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 047, W = 0.55, L = 0.5
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_47=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_47=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 048, W = 0.64, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_48=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_48=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 049, W = 0.84, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_49=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_49=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 050, W = 0.64, L = 0.18
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_50=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_50=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 051, W = 2.0, L = 0.15
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_51=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_51=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 052, W = 1.12, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_52=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_52=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 053, W = 1.65, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_53=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_53=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 054, W = 0.84, L = 0.18
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_54=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_54=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 055, W = 1.68, L = 0.18
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_55=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_55=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 056, W = 0.36, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_56=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_56=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 057, W = 0.54, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_57=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_57=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 058, W = 0.63, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_58=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_58=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 059, W = 0.7, L = 0.15
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_59=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_59=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 060, W = 0.75, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_60=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_60=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 061, W = 0.79, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_61=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_61=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 062, W = 0.82, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_62=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_62=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 063, W = 0.82, L = 0.18
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_63=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_63=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 064, W = 0.82, L = 0.25
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_64=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_64=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 065, W = 0.82, L = 0.5
* -----------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_65=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_65=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 066, W = 0.86, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_66=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_66=0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 067, W = 0.94, L = 0.15
* ------------------------------------
+  sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__keta_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ua_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__eta0_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pclm_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ub_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__ags_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b0_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__b1_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__agidl_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__a0_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__u0_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__voff_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__k2_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__kt1_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pdits_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vsat_diff_67=0.0
+  sky130_fd_pr__pfet_01v8_hvt__vth0_diff_67=0.0
.include "sky130_fd_pr__pfet_01v8_hvt.pm3.spice"
