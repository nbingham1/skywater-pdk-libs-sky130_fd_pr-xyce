* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre=0.0
* statistics {
*   process {
*   }
*   mismatch {
*     vary sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre dist=gauss std = 1.0
*   }
* }
.subckt sky130_fd_pr__nfet_g5v0d10v5 d g s b
.param l=1 w=1 ad=0 as=0 pd=0 ps=0 nrd=0 nrs=0 sa=0 sb=0 sd=0 mult=1 nf=1.0
msky130_fd_pr__nfet_g5v0d10v5 d g s b sky130_fd_pr__nfet_g5v0d10v5__model l={l} w={w} ad={ad} as={as} pd={pd} ps={ps} nrd={nrd} nrs={nrs} sa={sa} sb={sb} sd={sd} nf={nf}
.model sky130_fd_pr__nfet_g5v0d10v5__model.0 nmos
* DC IV MOS Parameters
+  lmin=2.0e-05 lmax=1.0e-04 wmin=2.0e-05 wmax=1.0e-4
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.793111+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+  k1=0.88325
+  k2=-0.0384371
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=105660.0
+  ua=-5.84299e-11
+  ub=1.6951e-18
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0418565
+  a0=0.94501626
+  keta=-0.02132
+  a1=0.0
+  a2=0.65972622
+  ags=0.1410462
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.92473+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.33405
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.4467e-5
+  alpha1=0.0
+  beta0=24.0
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.40273
+  kt2=-0.019151
+  at=160000.0
+  ute=-1.2986
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.1 nmos
* DC IV MOS Parameters
+  lmin=8e-06 lmax=2.0e-05 wmin=2.0e-05 wmax=1.0e-4
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.793111+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+  k1=0.88325
+  k2=-0.0384371
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=105660.0
+  ua=-5.84299e-11
+  ub=1.6951e-18
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0418565
+  a0=0.94501626
+  keta=-0.02132
+  a1=0.0
+  a2=0.65972622
+  ags=0.1410462
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.92473+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.33405
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.4467e-5
+  alpha1=0.0
+  beta0=24.0
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.40273
+  kt2=-0.019151
+  at=160000.0
+  ute=-1.2986
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.2 nmos
* DC IV MOS Parameters
+  lmin=4e-06 lmax=8e-06 wmin=2.0e-05 wmax=1.0e-4
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.788258849356+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=3.79066311535435e-8
+  k1=0.88325
+  k2=-0.0396087261612 lk2=9.15313723768459e-9
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=110425.42 lvsat=-0.03722906222112
+  ua=-1.009810976472e-10 lua=3.32424253222336e-16
+  ub=1.84142698652e-18 lub=-1.14315558456171e-24
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0419580987544 lu0=-7.9372360655426e-10
+  a0=1.03070800431664 la0=-6.69452699027683e-7
+  keta=-0.017304657108 lketa=-3.13692078275157e-8
+  a1=0.0
+  a2=0.65972622
+  ags=0.1570791696648 lags=-1.25254946099225e-7
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.96233869464+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-2.93811759049081e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.26057675444 lpclm=5.73997681325229e-7
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.4467e-5
+  alpha1=0.0
+  beta0=21.5219816 lbeta0=1.93591123549824e-5
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.414167008 lkt1=8.93497493306873e-8
+  kt2=-0.019151
+  at=236246.72 lat=-0.59566499553792
+  ute=-1.33672336 lute=2.97832497768961e-7
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.3 nmos
* DC IV MOS Parameters
+  lmin=2e-06 lmax=4e-06 wmin=2.0e-05 wmax=1.0e-4
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.805263767224+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-2.69218294116754e-8
+  k1=0.88325
+  k2=-0.0416511041712 lk2=1.6939368450816e-08 wk2=-2.11758236813575e-22
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=93909.0484 lvsat=0.0257368958189376
+  ua=1.047175735464e-10 lua=-4.51768196121188e-16 wua=9.86076131526265e-32 pua=3.76158192263132e-37
+  ub=1.49940600296e-18 lub=1.60743323819486e-25
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0422586227152 lu0=-1.93942192117469e-9
+  a0=0.4891605022816 la0=1.39510833869057e-6
+  keta=-0.039010436664 lketa=5.13805169818871e-8
+  a1=0.0
+  a2=0.65972622
+  ags=0.112641360624 lags=4.41569130681423e-8
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.92460675288+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.49964919127528e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.59742095576 lpclm=-7.10165593758256e-7
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.4467e-5
+  alpha1=0.0
+  beta0=23.910493376 lbeta0=1.02533029249137e-5
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.407041024 lkt1=6.21831039920641e-8
+  kt2=-0.019151
+  at=137994.752 lat=-0.221095480860672
+  ute=-1.22235328 lute=-1.3818467553792e-7
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.4 nmos
* DC IV MOS Parameters
+  lmin=1e-06 lmax=2e-06 wmin=2.0e-05 wmax=1.0e-4
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.788685223008+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=3.12406309857321e-9
+  k1=0.88325
+  k2=-0.0396502732144 lk2=1.33131904778928e-8
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=119403.907408 lvsat=-0.0204683549761851
+  ua=-1.4015488735776e-10 lua=-7.97701981598668e-18
+  ub=1.694312932e-18 lub=-1.92493520329152e-25
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.039851394944 lu0=2.42328362877081e-09 wu0=-2.11758236813575e-22
+  a0=1.6443791171696 la0=-6.98535944941084e-07 wa0=6.7762635780344e-21
+  keta=0.00275004268800001 lketa=-2.43035031249992e-8
+  a1=0.0
+  a2=0.65972622
+  ags=0.186902926464 lags=-9.04299961200599e-8
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.90605891408+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.16350003148091e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.10120107072 lpclm=1.89151567815598e-7
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.4467e-5
+  alpha1=0.0
+  beta0=27.186230848 lbeta0=4.31656597785907e-6
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.38085336 lkt1=1.472225776896e-8
+  kt2=-0.019151
+  at=9501.31199999999 lat=0.011777806215168
+  ute=-1.2986
+  ua1=3.0044e-9
+  ub1=-3.9963632672e-18 lub1=4.41962178224179e-25
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.81e-6
+  sbref=2.81e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.5 nmos
* DC IV MOS Parameters
+  lmin=8.0e-07 lmax=1e-06 wmin=2.0e-05 wmax=1.0e-4
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.80172216336+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-7.46631287920889e-9
+  k1=0.88325
+  k2=-0.034783520344 lk2=9.35975191816358e-9
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=109622.5588 lvsat=-0.0125226133733568
+  ua=-1.611781619232e-10 lua=9.10094295140447e-18
+  ub=7.526737312e-19 lub=5.72433901491917e-25
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.044773155776 lu0=-1.57483987845275e-9
+  a0=-0.24955524808 la0=8.39975121588315e-7
+  keta=-0.07771021344 lketa=4.10572594969958e-08 wketa=4.2351647362715e-22
+  a1=0.0
+  a2=0.65972622
+  ags=-0.18364432224 lags=2.10578873703153e-7
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.7226301416+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=3.26557921732223e-8
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-1.7899905 lpclm=1.725434563608e-06 ppclm=3.23117426778526e-27
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=5.60955976e-06 lalpha0=7.19521757480064e-12
+  alpha1=0.0
+  beta0=23.37007024 lbeta0=7.41657062151935e-6
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.33823656 lkt1=-1.989690307584e-8
+  kt2=-0.019151
+  at=8691.60000000001 lat=0.0124355644224
+  ute=-1.45627652 lute=1.2808631355072e-7
+  ua1=6.043729736e-09 lua1=-2.4689569604233e-15
+  ub1=-9.591886904e-18 lub1=4.98740746724774e-24
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.41e-6
+  sbref=2.41e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.6 nmos
* DC IV MOS Parameters
+  lmin=6e-07 lmax=8.0e-07 wmin=2.0e-05 wmax=1.0e-4
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.79360287968+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-2.4945831877327e-9
+  k1=0.88325
+  k2=-0.00691865331199999 lk2=-7.70290930074318e-9
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=76135.378856 lvsat=0.00798279244483238
+  ua=-2.80615603048e-10 lua=8.22367879000002e-17
+  ub=1.025401468e-18 lub=4.05432890050752e-25
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0359226803448 lu0=3.84462484518654e-9
+  a0=1.1222
+  keta=-0.01066
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.7171196528+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=3.60300628430592e-8
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=1.031511024 lpclm=-2.27239359206404e-9
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.67621128e-05 lalpha0=3.66107856499198e-13
+  alpha1=0.0
+  beta0=32.43483696 lbeta0=1.86588762726145e-6
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.37073
+  kt2=-0.019151
+  at=9620.208 lat=0.011866944314112
+  ute=-1.13989264 lute=-6.56469259929603e-8
+  ua1=2.0117e-9
+  ub1=-1.653168e-18 lub1=1.26244088448e-25
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.02e-6
+  sbref=2.01e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.7 nmos
* DC IV MOS Parameters
+  lmin=5e-07 lmax=6e-07 wmin=2.0e-05 wmax=1.0e-4
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.99226738448+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-8.44111104389452e-8
+  k1=0.88325
+  k2=0.00623535913600001 lk2=-1.31267821775017e-8
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=102214.584368 lvsat=-0.00277060283916364
+  ua=1.4315937032e-10 lua=-9.25008895186676e-17
+  ub=5.3820762016e-18 lub=-1.39098094290294e-24
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0496818299664 lu0=-1.8287678731855e-9
+  a0=1.1222
+  keta=-0.01066
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.8546985664+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-4.33034676075111e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.217674432 lpclm=3.33301731406848e-7
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=2.759165488e-05 lalpha0=-4.09930220659968e-12
+  alpha1=0.0
+  beta0=36.96
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.4331972 lkt1=2.57574753792001e-8
+  kt2=-0.019151
+  at=3418.36799999999 lat=0.014424186212352
+  ute=-1.30066168 lute=6.43936884480031e-10
+  ua1=-1.088859472e-09 lua1=1.27847229044659e-15
+  ub1=5.07306648e-18 lub1=-2.64722453209728e-24
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=1.81e-6
+  sbref=1.81e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.8 nmos
* DC IV MOS Parameters
+  lmin=2.0e-05 lmax=1.0e-04 wmin=1.5e-05 wmax=2.0e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.793111+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+  k1=0.88325
+  k2=-0.0384371
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=105660.0
+  ua=-5.84299e-11
+  ub=1.6951e-18
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0418565
+  a0=0.94501626
+  keta=-0.02132
+  a1=0.0
+  a2=0.65972622
+  ags=0.1410462
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.92473+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.33405
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.4467e-5
+  alpha1=0.0
+  beta0=24.0
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.40273
+  kt2=-0.019151
+  at=160000.0
+  ute=-1.2986
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.9 nmos
* DC IV MOS Parameters
+  lmin=8e-06 lmax=2.0e-05 wmin=1.5e-05 wmax=2.0e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.793111+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+  k1=0.88325
+  k2=-0.0384371
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=105660.0
+  ua=-5.84299e-11
+  ub=1.6951e-18
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0418565
+  a0=0.94501626
+  keta=-0.02132
+  a1=0.0
+  a2=0.65972622
+  ags=0.1410462
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.92473+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.33405
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.4467e-5
+  alpha1=0.0
+  beta0=24.0
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.40273
+  kt2=-0.019151
+  at=160000.0
+  ute=-1.2986
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.10 nmos
* DC IV MOS Parameters
+  lmin=4e-06 lmax=8e-06 wmin=1.5e-05 wmax=2.0e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.788258849356+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=3.79066311535443e-8
+  k1=0.88325
+  k2=-0.0396087261612 lk2=9.15313723768443e-9
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=110425.42 lvsat=-0.0372290622211207
+  ua=-1.009810976472e-10 lua=3.32424253222336e-16 pua=3.00926553810506e-36
+  ub=1.84142698652e-18 lub=-1.14315558456171e-24 wub=-2.35098870164458e-38
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0419580987544 lu0=-7.93723606554419e-10
+  a0=1.03070800431664 la0=-6.69452699027682e-07 wa0=1.35525271560688e-20
+  keta=-0.017304657108 lketa=-3.13692078275156e-8
+  a1=0.0
+  a2=0.65972622
+  ags=0.1570791696648 lags=-1.25254946099225e-7
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.962338694640001+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-2.93811759049078e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.26057675444 lpclm=5.73997681325227e-7
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.4467e-5
+  alpha1=0.0
+  beta0=21.5219816 lbeta0=1.93591123549823e-5
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.414167008 lkt1=8.93497493306868e-8
+  kt2=-0.019151
+  at=236246.72 lat=-0.59566499553792
+  ute=-1.33672336 lute=2.97832497768957e-7
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.11 nmos
* DC IV MOS Parameters
+  lmin=2e-06 lmax=4e-06 wmin=1.5e-05 wmax=2.0e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.805263767223999+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-2.69218294116758e-8
+  k1=0.88325
+  k2=-0.0416511041712 lk2=1.6939368450816e-8
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=93909.0484000001 lvsat=0.0257368958189377
+  ua=1.047175735464e-10 lua=-4.51768196121189e-16 pua=-1.1284745767894e-36
+  ub=1.49940600296e-18 lub=1.60743323819487e-25
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0422586227152 lu0=-1.93942192117469e-9
+  a0=0.4891605022816 la0=1.39510833869058e-6
+  keta=-0.039010436664 lketa=5.13805169818872e-8
+  a1=0.0
+  a2=0.65972622
+  ags=0.112641360624 lags=4.41569130681423e-8
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.92460675288+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.49964919127526e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.59742095576 lpclm=-7.10165593758256e-7
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.4467e-5
+  alpha1=0.0
+  beta0=23.910493376 lbeta0=1.02533029249137e-5
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.407041024 lkt1=6.21831039920639e-8
+  kt2=-0.019151
+  at=137994.752 lat=-0.221095480860672
+  ute=-1.22235328 lute=-1.38184675537918e-7
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.12 nmos
* DC IV MOS Parameters
+  lmin=1e-06 lmax=2e-06 wmin=1.5e-05 wmax=2.0e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.788121461336924+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=4.1457886704852e-09 wvth0=1.12874433717955e-08 pvth0=-2.04566399706748e-14
+  k1=0.88325
+  k2=-0.0382218329283343 lk2=1.07243767236057e-08 wk2=-2.85997428810288e-08 pk2=5.18323436140331e-14
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=126725.487551853 lvsat=-0.0337375182477747 wvsat=-0.146590173659812 pvsat=2.6567064896993e-7
+  ua=-1.46865750096547e-10 lua=4.18531831657549e-18 wua=1.34362598640933e-16 pua=-2.43510174570518e-22
+  ub=1.74915156727746e-18 lub=-2.91879553233358e-25 wub=-1.09796040071201e-24 pub=1.98987316078477e-30
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0389863502500038 lu0=3.99103526930906e-09 wu0=1.73196290179069e-08 pu0=-3.13889871757966e-14
+  a0=1.77253117495417 la0=-9.30790532738142e-07 wa0=-2.56581667295891e-06 pa0=4.65012192580365e-12
+  keta=0.00275004268800001 lketa=-2.43035031249992e-8
+  a1=0.0
+  a2=0.65972622
+  ags=-0.0256962366997688 lags=2.94871120851512e-07 wags=4.25658773595117e-06 pags=-7.7143671910228e-12
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.91486921551977+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.32317229618238e-07 wnfactor=-1.76396842303965e-07 pnfactor=3.19690347593812e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.10120107072 lpclm=1.89151567815598e-7
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.4467e-5
+  alpha1=0.0
+  beta0=27.2472440158654 lbeta0=4.2059896172625e-06 wbeta0=-1.22158478049837e-06 pbeta0=2.21392207474912e-12
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.38085336 lkt1=1.472225776896e-8
+  kt2=-0.019151
+  at=9501.31200000001 lat=0.011777806215168
+  ute=-1.2986
+  ua1=3.0044e-9
+  ub1=-3.9963632672e-18 lub1=4.41962178224178e-25
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.81e-6
+  sbref=2.81e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.13 nmos
* DC IV MOS Parameters
+  lmin=8.0e-07 lmax=1e-06 wmin=1.5e-05 wmax=2.0e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.804540971715383+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-9.19237071231057e-09 wvth0=-5.64372168590044e-08 pvth0=3.45585396225751e-14
+  k1=0.88325
+  k2=-0.0419257217743284 lk2=1.37331789732052e-08 wk2=1.42998714405146e-07 pk2=-8.75632607839899e-14
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=73014.6580807362 lvsat=0.00989372212147444 wvsat=0.732950868299056 pvsat=-4.48812202890772e-7
+  ua=-1.27623848229266e-10 lua=-1.14455712786844e-17 wua=-6.71812993204677e-16 pua=4.11375281006977e-22
+  ub=4.78480554812709e-19 lub=7.40332254348204e-25 wub=5.48980200355994e-24 pub=-3.36160339965189e-30
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.049098379245981 lu0=-4.22332991716704e-09 wu0=-8.65981450895336e-08 pu0=5.30271617715445e-14
+  a0=-0.89031553700285 la0=1.23233571386618e-06 wa0=1.28290833647945e-05 pa0=-7.85570959126481e-12
+  keta=-0.07771021344 lketa=4.10572594969958e-8
+  a1=0.0
+  a2=0.65972622
+  ags=0.879351493578842 lags=-4.40331732172093e-07 wags=-2.12829386797558e-05 pags=1.3032309539407e-11
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.678578634401152+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=5.96301158853361e-08 wnfactor=8.81984211519867e-07 pnfactor=-5.4007068414522e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-1.7899905 lpclm=1.725434563608e-06 ppclm=-6.46234853557053e-27
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=5.60955976e-06 lalpha0=7.19521757480063e-12
+  alpha1=0.0
+  beta0=23.0650044006728 lbeta0=7.60337341730962e-06 wbeta0=6.10792390249096e-06 pbeta0=-3.74010169075579e-12
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.33823656 lkt1=-1.98969030758398e-8
+  kt2=-0.019151
+  at=8691.59999999998 lat=0.0124355644224
+  ute=-1.45627652 lute=1.28086313550721e-7
+  ua1=6.043729736e-09 lua1=-2.4689569604233e-15
+  ub1=-9.591886904e-18 lub1=4.98740746724774e-24
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.41e-6
+  sbref=2.41e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.14 nmos
* DC IV MOS Parameters
+  lmin=6e-07 lmax=8.0e-07 wmin=1.5e-05 wmax=2.0e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.79360287968+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-2.49458318773206e-9
+  k1=0.88325
+  k2=-0.00691865331200001 lk2=-7.70290930074316e-9
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=76135.378856 lvsat=0.00798279244483241
+  ua=-2.80615603048e-10 lua=8.22367879000002e-17
+  ub=1.025401468e-18 lub=4.05432890050752e-25
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0359226803448 lu0=3.84462484518655e-9
+  a0=1.1222
+  keta=-0.01066
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.717119652799999+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=3.60300628430588e-8
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=1.031511024 lpclm=-2.27239359206341e-9
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.67621128e-05 lalpha0=3.66107856499192e-13
+  alpha1=0.0
+  beta0=32.43483696 lbeta0=1.86588762726144e-6
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.37073
+  kt2=-0.019151
+  at=9620.20799999998 lat=0.011866944314112
+  ute=-1.13989264 lute=-6.56469259929595e-8
+  ua1=2.0117e-9
+  ub1=-1.653168e-18 lub1=1.26244088448001e-25
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.02e-6
+  sbref=2.01e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.15 nmos
* DC IV MOS Parameters
+  lmin=5e-07 lmax=6e-07 wmin=1.5e-05 wmax=2.0e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={1.03974844675965+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-1.03989261735087e-07 wvth0=-9.50649590439865e-07 pvth0=3.91987049523615e-13
+  k1=0.88325
+  k2=0.0444970254295326 lk2=-2.89034446103118e-08 wk2=-7.66061997039237e-07 pk2=3.15874939611171e-13
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=153123.479068748 lvsat=-0.0237621728444914 wvsat=-1.0192804788564 pvsat=4.20286035529732e-7
+  ua=1.15955349044321e-10 lua=-8.12836922019391e-17 wua=5.44669610206366e-16 pua=-2.24586888394052e-22
+  ub=1.46218346195651e-17 lub=-5.200865969933e-24 wub=-1.84995283047118e-22 pub=7.62802150305166e-29
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.069020510055754 lu0=-9.8028018665094e-09 wu0=-3.87192438920456e-07 pu0=1.59653381494705e-13
+  a0=1.1222
+  keta=-0.01066
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={2.66013127385287+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-7.65143576935397e-07 wnfactor=-1.61260982106354e-05 pnfactor=6.64937083178056e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-1.71159560845378 lpclm=1.1288092228074e-06 wpclm=3.86271849396118e-05 ppclm=-1.59273789292598e-11
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=2.759165488e-05 lalpha0=-4.09930220659968e-12
+  alpha1=0.0
+  beta0=36.96
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.4331972 lkt1=2.57574753792004e-8
+  kt2=-0.019151
+  at=-71049.9541840527 lat=0.0451301563084355 wat=1.49097927860291 pat=-6.14784431822011e-7
+  ute=-1.30066168 lute=6.43936884479184e-10
+  ua1=-1.088859472e-09 lua1=1.27847229044659e-15
+  ub1=1.78880327883842e-18 lub1=-1.29300458078312e-24 wub1=6.57563945956425e-23 pub1=-2.71137287219889e-29
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=1.81e-6
+  sbref=1.81e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.16 nmos
* DC IV MOS Parameters
+  lmin=2.0e-05 lmax=1.0e-04 wmin=1.0e-05 wmax=1.5e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.793111+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+  k1=0.88325
+  k2=-0.0384371
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=105660.0
+  ua=-5.84299e-11
+  ub=1.6951e-18
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0418565
+  a0=0.94501626
+  keta=-0.02132
+  a1=0.0
+  a2=0.65972622
+  ags=0.1410462
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.92473+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.33405
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.4467e-5
+  alpha1=0.0
+  beta0=24.0
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.40273
+  kt2=-0.019151
+  at=160000.0
+  ute=-1.2986
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.17 nmos
* DC IV MOS Parameters
+  lmin=8e-06 lmax=2.0e-05 wmin=1.0e-05 wmax=1.5e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.793111+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+  k1=0.88325
+  k2=-0.0384371
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=105660.0
+  ua=-5.84299e-11
+  ub=1.6951e-18
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0418565
+  a0=0.94501626
+  keta=-0.02132
+  a1=0.0
+  a2=0.65972622
+  ags=0.1410462
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.92473+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.33405
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.4467e-5
+  alpha1=0.0
+  beta0=24.0
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.40273
+  kt2=-0.019151
+  at=160000.0
+  ute=-1.2986
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.18 nmos
* DC IV MOS Parameters
+  lmin=4e-06 lmax=8e-06 wmin=1.0e-05 wmax=1.5e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.788258849356+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=3.79066311535443e-8
+  k1=0.88325
+  k2=-0.0396087261612 lk2=9.15313723768475e-9
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=110425.42 lvsat=-0.0372290622211202
+  ua=-1.009810976472e-10 lua=3.32424253222336e-16
+  ub=1.84142698652e-18 lub=-1.14315558456171e-24
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0419580987544 lu0=-7.93723606554313e-10
+  a0=1.03070800431664 la0=-6.69452699027682e-7
+  keta=-0.017304657108 lketa=-3.13692078275156e-8
+  a1=0.0
+  a2=0.65972622
+  ags=0.1570791696648 lags=-1.25254946099225e-7
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.96233869464+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-2.93811759049078e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.26057675444 lpclm=5.73997681325229e-7
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.4467e-5
+  alpha1=0.0
+  beta0=21.5219816 lbeta0=1.93591123549823e-5
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.414167008 lkt1=8.93497493306885e-8
+  kt2=-0.019151
+  at=236246.72 lat=-0.59566499553792
+  ute=-1.33672336 lute=2.97832497768957e-7
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.19 nmos
* DC IV MOS Parameters
+  lmin=2e-06 lmax=4e-06 wmin=1.0e-05 wmax=1.5e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.805263767224+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-2.69218294116741e-8
+  k1=0.88325
+  k2=-0.0416511041712 lk2=1.6939368450816e-8
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=93909.0484 lvsat=0.0257368958189377
+  ua=1.047175735464e-10 lua=-4.51768196121189e-16 wua=9.86076131526265e-32 pua=1.31655367292096e-36
+  ub=1.49940600296e-18 lub=1.60743323819484e-25
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0422586227152 lu0=-1.93942192117469e-9
+  a0=0.4891605022816 la0=1.39510833869057e-6
+  keta=-0.039010436664 lketa=5.13805169818871e-8
+  a1=0.0
+  a2=0.65972622
+  ags=0.112641360624 lags=4.41569130681423e-8
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.92460675288+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.49964919127526e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.59742095576 lpclm=-7.10165593758256e-7
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.4467e-5
+  alpha1=0.0
+  beta0=23.910493376 lbeta0=1.02533029249137e-5
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.407041024 lkt1=6.2183103992063e-8
+  kt2=-0.019151
+  at=137994.752 lat=-0.221095480860672
+  ute=-1.22235328 lute=-1.38184675537919e-7
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.20 nmos
* DC IV MOS Parameters
+  lmin=1e-06 lmax=2e-06 wmin=1.0e-05 wmax=1.5e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.783680572435085+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=1.21941714992884e-08 wvth0=7.79969576712294e-08 pvth0=-1.4135669427804e-13
+  k1=0.88325
+  k2=-0.0395307925880787 lk2=1.30966514375082e-08 wk2=-8.93699853655237e-09 pk2=1.61968441797412e-14
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=123842.74879583 lvsat=-0.0285130270216396 wvsat=-0.103286657963494 pvsat=1.87190128546926e-7
+  ua=-1.25745710973561e-10 lua=-3.40912889074203e-17 wua=-1.82895406011178e-16 pua=3.31467928548677e-22
+  ub=1.86750240630474e-18 lub=-5.06371039432703e-25 wub=-2.87578622859284e-24 pub=5.21189091038304e-30
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0392141080656185 lu0=3.57826158078913e-09 wu0=1.38983290049147e-08 pu0=-2.51884419954513e-14
+  a0=2.3309313600211 la0=-1.94279929054159e-06 wa0=-1.0953913280171e-05 pa0=1.9852171378532e-11
+  keta=0.0296282150049073 lketa=-7.30157824291338e-08 wketa=-4.0375471220965e-07 pketa=7.31739200107188e-13
+  a1=0.0
+  a2=0.65972622
+  ags=0.387363927850294 lags=-4.53732685528491e-07 wags=-1.9482607893436e-06 pags=3.53090316591581e-12
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.933361882690448+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.65832156067677e-07 wnfactor=-4.54187364049744e-07 pnfactor=8.23140110612459e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.728770899762208 lpclm=-9.4821582587144e-07 wpclm=-9.42713934299051e-06 ppclm=1.70851440083181e-11
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.25831833431874e-05 lalpha0=3.41410874454105e-12 walpha0=2.82980495533417e-11 palpha0=-5.12855739353052e-17
+  alpha1=0.0
+  beta0=27.6136748945198 lbeta0=3.54189374436552e-06 wbeta0=-6.72598412028414e-06 pbeta0=1.21897431566195e-11
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.397135267146176 lkt1=4.42305442386322e-08 wkt1=2.44581240737611e-07 pkt1=-4.43263387513441e-13
+  kt2=-0.019151
+  at=9501.31199999999 lat=0.011777806215168
+  ute=-1.2986
+  ua1=3.0044e-9
+  ub1=-4.48514611972821e-18 lub1=1.32780093804373e-24 wub1=7.34232884694311e-24 pub1=-1.33067668931535e-29
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.81e-6
+  sbref=2.81e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.21 nmos
* DC IV MOS Parameters
+  lmin=8.0e-07 lmax=1e-06 wmin=1.0e-05 wmax=1.5e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.826745416224577+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-2.27889514452931e-08 wvth0=-3.89984788356126e-07 pvth0=2.38801725362838e-13
+  k1=0.88325
+  k2=-0.0353809234756064 lk2=9.72556336215891e-09 wk2=4.46849926827619e-08 pk2=-2.73622296793917e-14
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=87428.3518608494 lvsat=0.00106769852693478 wvsat=0.516433289817467 pvsat=-3.16230694953669e-7
+  ua=-2.33224043844195e-10 lua=5.32172301033789e-17 wua=9.14477030055895e-16 pua=-5.59967206676306e-22
+  ub=-1.13273640323688e-19 lub=1.10268465118124e-24 wub=1.43789311429642e-23 pub=-8.80473718035812e-30
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0479595901679072 lu0=-3.52600836825568e-09 wu0=-6.94916450245733e-08 pu0=4.25522359477674e-14
+  a0=-3.68231646233748 la0=2.94197839248188e-06 wa0=5.47695664008549e-05 pa0=-3.35373772116339e-11
+  keta=-0.212101075024537 lketa=1.23349622116225e-07 wketa=2.01877356104825e-06 pketa=-1.23616772727804e-12
+  a1=0.0
+  a2=0.65972622
+  ags=-1.18594932917147 lags=8.24326312427541e-07 wags=9.74130394671797e-06 pags=-5.96495109351749e-12
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.586115298547755+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.16248745108461e-07 wnfactor=2.27093682024873e-06 pnfactor=-1.39057636876382e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-4.92783964521104 lpclm=3.64685255778994e-06 wpclm=4.71356967149525e-05 ppclm=-2.88628839836472e-11
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.50286430440628e-05 lalpha0=1.42757379297076e-12 walpha0=-1.41490247766708e-10 palpha0=8.66395723564753e-17
+  alpha1=0.0
+  beta0=21.2328500074008 lbeta0=8.72526750986819e-06 wbeta0=3.36299206014209e-05 pbeta0=-2.0592811061392e-11
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.25682702426912 lkt1=-6.97468925471441e-08 wkt1=-1.22290620368806e-06 pkt1=7.48829493141529e-13
+  kt2=-0.019151
+  at=8691.59999999992 lat=0.0124355644224
+  ute=-1.45627652 lute=1.28086313550721e-7
+  ua1=6.043729736e-09 lua1=-2.4689569604233e-15
+  ub1=-7.14797264135899e-18 lub1=3.4909107833192e-24 wub1=-3.67116442347155e-23 pub1=2.24798613841087e-29
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.41e-6
+  sbref=2.41e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.22 nmos
* DC IV MOS Parameters
+  lmin=6e-07 lmax=8.0e-07 wmin=1.0e-05 wmax=1.5e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.793602879679999+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-2.49458318773248e-9
+  k1=0.88325
+  k2=-0.00691865331200001 lk2=-7.70290930074316e-9
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=76135.3788559999 lvsat=0.00798279244483241
+  ua=-2.80615603048e-10 lua=8.22367879000002e-17
+  ub=1.025401468e-18 lub=4.05432890050751e-25
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0359226803448001 lu0=3.84462484518655e-9
+  a0=1.1222
+  keta=-0.01066
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.7171196528+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=3.60300628430597e-8
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=1.031511024 lpclm=-2.27239359206341e-9
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.67621128e-05 lalpha0=3.66107856499218e-13
+  alpha1=0.0
+  beta0=32.43483696 lbeta0=1.86588762726144e-6
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.37073
+  kt2=-0.019151
+  at=9620.20799999998 lat=0.011866944314112
+  ute=-1.13989264 lute=-6.56469259929595e-8
+  ua1=2.0117e-9
+  ub1=-1.653168e-18 lub1=1.26244088448e-25
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.02e-6
+  sbref=2.01e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.23 nmos
* DC IV MOS Parameters
+  lmin=5e-07 lmax=6e-07 wmin=1.0e-05 wmax=1.5e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.974146890695916+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-7.69393785139906e-08 wvth0=3.47945490173935e-08 pvth0=-1.43470451636387e-14
+  k1=0.88325
+  k2=-0.00154264996514331 lk2=-9.91962901677271e-09 wk2=-7.44697388294024e-08 pk2=3.07065542299603e-14
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=74524.9537504183 lvsat=0.00864682869116756 wvsat=0.1613996877799 pvsat=-6.65509016604134e-8
+  ua=1.85836285987859e-10 lua=-1.1009811821749e-16 wua=-5.05057925279025e-16 pua=2.08253564677853e-22
+  ub=3.06619090080042e-18 lub=-4.36058061512439e-25 wub=-1.14103551339871e-23 pub=4.70490019452769e-30
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.041941889085115 lu0=1.36268839004005e-09 wu0=1.95733444121125e-08 pu0=-8.07079454151293e-15
+  a0=1.1222
+  keta=-0.01066
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.61701411426298+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-3.35028819818739e-07 wnfactor=-4.56748985344622e-07 pnfactor=1.88334049621062e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=2.14694447245379 lpclm=-4.62205759993706e-07 wpclm=-1.9334484535074e-05 ppclm=7.97230401525429e-12
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=2.759165488e-05 lalpha0=-4.09930220659967e-12
+  alpha1=0.0
+  beta0=36.96
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.4331972 lkt1=2.57574753792002e-8
+  kt2=-0.019151
+  at=77886.6901840529 lat=-0.0162817838837316 wat=-0.74629605676239 pat=3.07724730861177e-7
+  ute=-1.30066168 lute=6.43936884480878e-10
+  ua1=-1.088859472e-09 lua1=1.27847229044659e-15
+  ub1=6.16624248e-18 lub1=-3.09798035123328e-24
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=1.81e-6
+  sbref=1.81e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.24 nmos
* DC IV MOS Parameters
+  lmin=2.0e-05 lmax=1.0e-04 wmin=7e-06 wmax=1.0e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.793111+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+  k1=0.88325
+  k2=-0.0384371
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=105660.0
+  ua=-5.84299e-11
+  ub=1.6951e-18
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0418565
+  a0=0.94501626
+  keta=-0.02132
+  a1=0.0
+  a2=0.65972622
+  ags=0.1410462
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.92473+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.33405
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.4467e-5
+  alpha1=0.0
+  beta0=24.0
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.40273
+  kt2=-0.019151
+  at=160000.0
+  ute=-1.2986
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.25 nmos
* DC IV MOS Parameters
+  lmin=8e-06 lmax=2.0e-05 wmin=7e-06 wmax=1.0e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.793111+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+  k1=0.88325
+  k2=-0.0384371
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=105660.0
+  ua=-5.84299e-11
+  ub=1.6951e-18
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0418565
+  a0=0.94501626
+  keta=-0.02132
+  a1=0.0
+  a2=0.65972622
+  ags=0.1410462
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.92473+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.33405
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.4467e-5
+  alpha1=0.0
+  beta0=24.0
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.40273
+  kt2=-0.019151
+  at=160000.0
+  ute=-1.2986
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.26 nmos
* DC IV MOS Parameters
+  lmin=4e-06 lmax=8e-06 wmin=7e-06 wmax=1.0e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.788258849356001+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=3.79066311535443e-8
+  k1=0.88325
+  k2=-0.0396087261612 lk2=9.15313723768475e-9
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=110425.42 lvsat=-0.0372290622211202
+  ua=-1.009810976472e-10 lua=3.32424253222336e-16
+  ub=1.84142698652e-18 lub=-1.14315558456171e-24
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0419580987544 lu0=-7.93723606554207e-10
+  a0=1.03070800431664 la0=-6.69452699027682e-7
+  keta=-0.017304657108 lketa=-3.13692078275156e-8
+  a1=0.0
+  a2=0.65972622
+  ags=0.1570791696648 lags=-1.25254946099225e-7
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.962338694640001+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-2.93811759049081e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.26057675444 lpclm=5.73997681325229e-7
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.4467e-5
+  alpha1=0.0
+  beta0=21.5219816 lbeta0=1.93591123549825e-5
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.414167008 lkt1=8.93497493306868e-8
+  kt2=-0.019151
+  at=236246.72 lat=-0.59566499553792
+  ute=-1.33672336 lute=2.97832497768964e-7
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.27 nmos
* DC IV MOS Parameters
+  lmin=2e-06 lmax=4e-06 wmin=7e-06 wmax=1.0e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.805263767223999+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-2.69218294116758e-8
+  k1=0.88325
+  k2=-0.0416511041712 lk2=1.6939368450816e-8
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=93909.0484000001 lvsat=0.0257368958189377
+  ua=1.047175735464e-10 lua=-4.51768196121188e-16 pua=-3.76158192263132e-37
+  ub=1.49940600296e-18 lub=1.60743323819487e-25
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0422586227152 lu0=-1.93942192117469e-9
+  a0=0.489160502281599 la0=1.39510833869057e-6
+  keta=-0.039010436664 lketa=5.13805169818872e-8
+  a1=0.0
+  a2=0.65972622
+  ags=0.112641360624 lags=4.41569130681423e-8
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.92460675288+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.49964919127526e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.59742095576 lpclm=-7.10165593758255e-7
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.4467e-5
+  alpha1=0.0
+  beta0=23.910493376 lbeta0=1.02533029249137e-5
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.407041024 lkt1=6.21831039920647e-8
+  kt2=-0.019151
+  at=137994.752 lat=-0.221095480860672
+  ute=-1.22235328 lute=-1.38184675537921e-7
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.28 nmos
* DC IV MOS Parameters
+  lmin=1e-06 lmax=2e-06 wmin=7e-06 wmax=1.0e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.791463412128+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-1.91094905841112e-9
+  k1=0.88325
+  k2=-0.0404225610496 lk2=1.47128355239879e-8
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=113536.40448 lvsat=-0.00983446818966538
+  ua=-1.439957256928e-10 lua=-1.01613023121362e-18
+  ub=1.5805452752e-18 lub=1.36916997251329e-26
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0406009373712 lu0=1.06486090442886e-9
+  a0=1.2379073035056 la0=3.81275559474756e-8
+  keta=-0.01066
+  a1=0.0
+  a2=0.65972622
+  ags=0.192958891344 lags=-1.0140543928682e-7
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.888041301599999+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-8.36960354165376e-8
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-0.21190571712 lpclm=7.56606271262393e-07 ppclm=-1.61558713389263e-27
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.5406872752e-05 lalpha0=-1.70336522386868e-12
+  alpha1=0.0
+  beta0=26.942530048 lbeta0=4.75823371092789e-6
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.37273
+  kt2=-0.019151
+  at=9501.31199999999 lat=0.011777806215168
+  ute=-1.2986
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.81e-6
+  sbref=2.81e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.29 nmos
* DC IV MOS Parameters
+  lmin=8.0e-07 lmax=1e-06 wmin=7e-06 wmax=1.0e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.787831217759999+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=1.03961318571207e-9
+  k1=0.88325
+  k2=-0.030922081168 lk2=6.9952536988884e-9
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=138960.07344 lvsat=-0.0304870297379557
+  ua=-1.41973970248e-10 lua=-2.65847496222067e-18
+  ub=1.3215120152e-18 lub=2.24113742020493e-25
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.04102544364 lu0=7.20019180056902e-10
+  a0=1.78280382024 la0=-4.04511500870481e-7
+  keta=-0.01066
+  a1=0.0
+  a2=0.65972622
+  ags=-0.21392414664 lags=2.29120300256951e-7
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.812718203999999+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-2.25083716045437e-8
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-0.2244565608 lpclm=7.66801773414029e-7
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=9.1019600000002e-07 lalpha0=1.0072807182144e-11
+  alpha1=0.0
+  beta0=24.58857424 lbeta0=6.67043675617535e-6
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.37885336 lkt1=4.97422576895975e-9
+  kt2=-0.019151
+  at=8691.59999999998 lat=0.0124355644224
+  ute=-1.45627652 lute=1.28086313550721e-7
+  ua1=6.043729736e-09 lua1=-2.4689569604233e-15
+  ub1=-1.081120324e-17 lub1=5.73403875516864e-24
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.41e-6
+  sbref=2.41e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.30 nmos
* DC IV MOS Parameters
+  lmin=6e-07 lmax=8.0e-07 wmin=7e-06 wmax=1.0e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.79360287968+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-2.49458318773248e-9
+  k1=0.88325
+  k2=-0.00691865331200001 lk2=-7.70290930074318e-9
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=76135.3788559999 lvsat=0.00798279244483246
+  ua=-2.80615603048e-10 lua=8.22367879000001e-17
+  ub=1.025401468e-18 lub=4.05432890050752e-25
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0359226803448 lu0=3.84462484518658e-9
+  a0=1.1222
+  keta=-0.01066
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.717119652799999+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=3.60300628430592e-8
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=1.031511024 lpclm=-2.27239359206426e-9
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.67621128e-05 lalpha0=3.66107856499205e-13
+  alpha1=0.0
+  beta0=32.43483696 lbeta0=1.86588762726144e-6
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.37073
+  kt2=-0.019151
+  at=9620.20799999998 lat=0.011866944314112
+  ute=-1.13989264 lute=-6.56469259929595e-8
+  ua1=2.0117e-9
+  ub1=-1.653168e-18 lub1=1.26244088447999e-25
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.02e-6
+  sbref=2.01e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.31 nmos
* DC IV MOS Parameters
+  lmin=5e-07 lmax=6e-07 wmin=7e-06 wmax=1.0e-5
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.961243555667611+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-7.1618868961759e-08 wvth0=1.64107359730501e-07 pvth0=-6.7667372281834e-14
+  k1=0.88325
+  k2=-0.0321357652152401 lk2=2.69501375299124e-09 wk2=2.32123999361653e-07 pk2=-9.57130814007865e-14
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=94464.3409366158 lvsat=0.000425101536359718 wvsat=-0.0384260313297524 pvsat=1.58444360543848e-8
+  ua=1.59282401750269e-10 lua=-9.91489958064991e-17 wua=-2.38943978878309e-16 pua=9.85252044747666e-23
+  ub=4.89230552649467e-18 lub=-1.1890308618127e-24 wub=-2.97110513814929e-23 pub=1.22509360824393e-29
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0445835589928638 lu0=2.73432786958509e-10 wu0=-6.9005679522386e-09 pu0=2.84535258715446e-15
+  a0=1.1222
+  keta=-0.01066
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={2.22614901520396+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-5.86197068333141e-07 wnfactor=-6.56129063843905e-06 pnfactor=2.70545633669141e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.217674432000001 lpclm=3.33301731406847e-7
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=2.759165488e-05 lalpha0=-4.09930220659968e-12
+  alpha1=0.0
+  beta0=36.96
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.4331972 lkt1=2.57574753792e-8
+  kt2=-0.019151
+  at=-66761.3623388162 lat=0.0433618155013381 wat=0.70331725598784 pat=-2.90003024065002e-7
+  ute=-1.30066168 lute=6.43936884480031e-10
+  ua1=-1.088859472e-09 lua1=1.27847229044659e-15
+  ub1=7.628320195392e-18 lub1=-3.70084762808716e-24 wub1=-1.465244283308e-23 pub1=6.04172966802085e-30
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=1.81e-6
+  sbref=1.81e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.32 nmos
* DC IV MOS Parameters
+  lmin=2.0e-05 lmax=1.0e-04 wmin=5.0e-06 wmax=7.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.776604810154+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} wvth0=1.15900819981683e-7
+  k1=0.88325
+  k2=-0.0369901092473 wk2=-1.01602741946219e-8
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=119394.23463 wvsat=-0.0964370984636167
+  ua=-3.8164891717e-10 wua=2.26953339766387e-15
+  ub=2.14742584435e-18 wub=-3.17607738358693e-24
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0412646976047 wu0=4.15543402337759e-9
+  a0=1.23137349532152 wa0=-2.01070257225324e-6
+  keta=-0.016973755001 wketa=-3.05178459671884e-8
+  a1=0.0
+  a2=0.65972622
+  ags=0.168954064335 wags=-1.95959478870767e-7
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.85259388283+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} wnfactor=5.06515144215664e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.65757031665 wpclm=-2.27164901956801e-6
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=2.3910227869e-05 walpha0=-6.63071165121868e-11
+  alpha1=0.0
+  beta0=26.724249465 wbeta0=-1.91287480499129e-5
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.40273
+  kt2=-0.019151
+  at=180086.632 wat=-0.141041460275856
+  ute=-1.2986
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.33 nmos
* DC IV MOS Parameters
+  lmin=8e-06 lmax=2.0e-05 wmin=5.0e-06 wmax=7.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.776604810154+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} wvth0=1.15900819981683e-7
+  k1=0.88325
+  k2=-0.0369901092473 wk2=-1.01602741946219e-8
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=119394.23463 wvsat=-0.0964370984636167
+  ua=-3.8164891717e-10 wua=2.26953339766387e-15
+  ub=2.14742584435e-18 wub=-3.17607738358694e-24
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0412646976047 wu0=4.15543402337749e-9
+  a0=1.23137349532152 wa0=-2.01070257225323e-6
+  keta=-0.016973755001 wketa=-3.05178459671884e-8
+  a1=0.0
+  a2=0.65972622
+  ags=0.168954064335 wags=-1.95959478870768e-7
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.852593882830001+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} wnfactor=5.06515144215661e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.65757031665 wpclm=-2.27164901956801e-6
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=2.3910227869e-05 walpha0=-6.63071165121868e-11
+  alpha1=0.0
+  beta0=26.724249465 wbeta0=-1.9128748049913e-5
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.40273
+  kt2=-0.019151
+  at=180086.632 wat=-0.141041460275856
+  ute=-1.2986
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.34 nmos
* DC IV MOS Parameters
+  lmin=4e-06 lmax=8e-06 wmin=5.0e-06 wmax=7.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.76736384075387+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=7.21935579195349e-08 wvth0=1.46717604311214e-07 pvth0=-2.40751073621845e-13
+  k1=0.88325
+  k2=-0.0336257452491515 lk2=-2.62835419798394e-08 wk2=-4.20104457849326e-08 pk2=2.48824242121163e-13
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=142418.480752833 lvsat=-0.179873146858266 wvsat=-0.224644330979614 pvsat=1.00159797804509e-6
+  ua=-5.30977394959193e-10 lua=1.16660424285771e-15 wua=3.01928694099113e-15 pua=-5.85732659766316e-21
+  ub=2.43477414455526e-18 lub=-2.24486147023235e-24 wub=-4.16628081899554e-24 pub=7.7358019457664e-30
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0409164065411324 lu0=2.72096681438726e-09 wu0=7.3144064628282e-09 pu0=-2.46789541117275e-14
+  a0=1.53508849805127 la0=-2.37272364956577e-06 wa0=-3.54158732887575e-06 pa0=1.19597860960133e-11
+  keta=-0.00287657273082251 lketa=-1.10131924547869e-07 wketa=-1.01309074091683e-07 pketa=5.53044859961204e-13
+  a1=0.0
+  a2=0.65972622
+  ags=0.218716805192635 lags=-3.88763251860769e-07 wags=-4.32798396605103e-07 pags=1.85026520321699e-12
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.886876264454175+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-2.67825484128287e-07 wnfactor=5.29871376613729e-07 pnfactor=-1.82466735187745e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.39961831541383 lpclm=2.01520770552937e-06 wpclm=-9.76302288944385e-07 ppclm=-1.01196838961332e-11
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=3.56791540645559e-05 lalpha0=-9.1942805798884e-11 walpha0=-1.48944491284621e-10 palpha0=6.4559093788018e-16
+  alpha1=0.0
+  beta0=26.868992982513 lbeta0=-1.13078499263384e-06 wbeta0=-3.75448852501139e-05 pbeta0=1.43873051630069e-10
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.414167008 lkt1=8.93497493306885e-8
+  kt2=-0.019151
+  at=275477.599573088 lat=-0.745226290046068 wat=-0.275465819401409 pat=1.0501682600735e-6
+  ute=-1.33672336 lute=2.97832497768957e-7
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.35 nmos
* DC IV MOS Parameters
+  lmin=2e-06 lmax=4e-06 wmin=5.0e-06 wmax=7.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.791175938953565+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-1.85861612826966e-08 wvth0=9.8919912077724e-08 pvth0=-5.8530210803175e-14
+  k1=0.88325
+  k2=-0.0478256327677362 lk2=2.78512004032114e-08 wk2=4.33554281160971e-08 pk2=-7.66191521231938e-14
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=73196.092717212 lvsat=0.084025855055899 wvsat=0.145439290973693 pvsat=-4.09285136937885e-7
+  ua=1.17508881255757e-10 lua=-1.30564333346248e-15 wua=-8.9816188107868e-17 pua=5.99561918911361e-21
+  ub=1.70950579557174e-18 lub=5.20105166258072e-25 wub=-1.47524888959057e-24 pub=-2.52331595585366e-30
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0435456326698101 lu0=-7.30252660811118e-09 wu0=-9.03694374386762e-09 pu0=3.76578869298654e-14
+  a0=0.288472353273105 la0=2.37979595735327e-06 wa0=1.40916354699069e-06 pa0=-6.91413969508383e-12
+  keta=-0.0508894422831011 lketa=7.29092665095863e-08 wketa=8.34103148374063e-08 pketa=-1.51167516351165e-13
+  a1=0.0
+  a2=0.65972622
+  ags=0.118576138575625 lags=-6.99338345274517e-09 wags=-4.16719810822501e-08 pags=3.59159888768263e-13
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.830819364549343+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-5.41177465727e-08 wnfactor=6.58542965571057e-07 pnfactor=-6.7300606594698e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=1.58222070588992 lpclm=-2.4932699613687e-06 wpclm=-6.91492704389779e-06 ppclm=1.25203490476668e-11
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=8.92952638948431e-06 lalpha0=1.00357627733876e-11 walpha0=3.88822458770665e-11 palpha0=-7.04676939638593e-17
+  alpha1=0.0
+  beta0=23.857846695174 lbeta0=1.03487163998552e-05 wbeta0=3.6966698759521e-07 pbeta0=-6.69960789630321e-13
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.407041024 lkt1=6.21831039920647e-8
+  kt2=-0.019151
+  at=147095.683573088 lat=-0.255791289930292 wat=-0.0639036289876258 pat=2.4362210532017e-7
+  ute=-1.22235328 lute=-1.38184675537921e-7
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.36 nmos
* DC IV MOS Parameters
+  lmin=1e-06 lmax=2e-06 wmin=5.0e-06 wmax=7.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.773891908751926+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=1.27383088768192e-08 wvth0=1.23381087252634e-07 pvth0=-1.02862079174971e-13
+  k1=0.88325
+  k2=-0.0385906373726994 lk2=1.11142857889521e-08 wk2=-1.28631415412985e-08 pk2=2.5267785535412e-14
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=125673.142317065 lvsat=-0.0110801911077003 wvsat=-0.0852200223275328 pvsat=8.74704029320424e-9
+  ua=-9.79902027211758e-10 lua=6.83233962745898e-16 wua=5.86944816931101e-15 pua=-4.80457013935348e-21
+  ub=2.29960908737638e-18 lub=-5.49360273197983e-25 wub=-5.0490201692788e-24 pub=3.95355839009138e-30
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0364205839007869 lu0=5.6104557777453e-09 wu0=2.93530123883543e-08 pu0=-3.19176126069811e-14
+  a0=1.59274671740178 la0=1.60125733657515e-08 wa0=-2.49156100929945e-06 pa0=1.55283844364818e-13
+  keta=-0.01066
+  a1=0.0
+  a2=0.65972622
+  ags=0.14972523214998 lags=-6.34460071049165e-08 wags=3.03571968948967e-07 pags=-2.66538150655517e-13
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.830006948183031+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-5.26453751450426e-08 wnfactor=4.07497381945087e-07 pnfactor=-2.18027117100623e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.156647424016692 lpclm=9.03478180083073e-08 wpclm=-2.58785411188758e-06 ppclm=4.67823899835917e-12
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=4.72741579049635e-05 lalpha0=-5.94575933288499e-11 walpha0=-2.23761177732588e-10 palpha0=4.05530437807166e-16
+  alpha1=0.0
+  beta0=32.6535130503232 lbeta0=-5.5919863795706e-06 wbeta0=-4.01005694861268e-05 pbeta0=7.26757057002091e-11
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.37273
+  kt2=-0.019151
+  at=3537.26957308804 lat=0.00438479186481198 wat=0.0418774662192659 pat=5.19112183572921e-8
+  ute=-1.2986
+  ua1=3.0044e-9
+  ub1=-3.1406089640368e-18 lub1=-1.1089521525534e-24 wub1=-4.2964895877993e-24 pub1=7.78668275359383e-30
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.81e-6
+  sbref=2.81e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.37 nmos
* DC IV MOS Parameters
+  lmin=8.0e-07 lmax=1e-06 wmin=5.0e-06 wmax=7.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.788938948110349+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=5.15057112556408e-10 wvth0=-7.77810367636855e-09 pvth0=3.68325334752087e-15
+  k1=0.88325
+  k2=-0.0343694886543655 lk2=7.68529472369559e-09 wk2=2.42065163558985e-08 pk2=-4.8452320821653e-15
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=203346.345622789 lvsat=-0.0741769303882586 wvsat=-0.452098383162458 pvsat=3.06775540420404e-7
+  ua=-1.18242830544528e-10 lua=-1.67228224379739e-17 wua=-1.66631946948003e-16 pua=9.8755037967903e-23
+  ub=1.10345223320547e-18 lub=4.22321001091803e-25 wub=1.53114121272017e-24 pub=-1.39174358631614e-30
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0437453420793826 lu0=-3.39708982022485e-10 wu0=-1.90981966360783e-08 pu0=7.44104872709063e-15
+  a0=3.11347305796524 la0=-1.2193281792222e-06 wa0=-9.3435042984273e-06 pa0=5.72136404808179e-12
+  keta=-0.01066
+  a1=0.0
+  a2=0.65972622
+  ags=-0.199728274605654 lags=2.20427656758928e-07 wags=-9.96785584369424e-08 pags=6.10367697590443e-14
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.824810286160789+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-4.84239395045419e-08 wnfactor=-8.49064654409584e-08 pnfactor=1.81970254669562e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-3.5992729597461 lpclm=3.14141715887264e-06 wpclm=2.36968065661911e-05 ppclm=-1.66737371182286e-11
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=-0.000136179024589526 lalpha0=8.95680311259934e-11 walpha0=9.62593622466207e-10 palpha0=-5.58188275167122e-16
+  alpha1=0.0
+  beta0=-3.96634077161605 lbeta0=2.41556391947283e-05 wbeta0=0.000200502847430634 pbeta0=-1.22775111584285e-10
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.378853359999999 lkt1=4.97422576896059e-9
+  kt2=-0.019151
+  at=-52497.50359632 lat=0.0499038553621562 wat=0.429648958779929 pat=-2.63089524823467e-7
+  ute=-1.45627652 lute=1.28086313550719e-7
+  ua1=6.043729736e-09 lua1=-2.4689569604233e-15
+  ub1=-1.24100609825992e-17 lub1=6.4209574223975e-24 wub1=1.12266322591836e-23 pub1=-4.82330795509689e-30
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.41e-6
+  sbref=2.41e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.38 nmos
* DC IV MOS Parameters
+  lmin=6e-07 lmax=8.0e-07 wmin=5.0e-06 wmax=7.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.794371615173271+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-2.81156050608631e-09 wvth0=-5.39779772621422e-09 pvth0=2.22570632323883e-15
+  k1=0.88325
+  k2=-0.0140233067408198 lk2=-4.77340492451729e-09 wk2=4.98864465857003e-08 pk2=-2.05699778393613e-14
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=54816.0374210876 lvsat=0.0167735244147384 wvsat=0.149697124341184 pvsat=-6.17255134623465e-8
+  ua=-2.7828018461944e-10 lua=8.12738108068413e-17 wua=-1.63985094922476e-17 pua=6.76169580999544e-24
+  ub=1.34880849001953e-18 lub=2.72080532219307e-25 wub=-2.27085350341961e-24 pub=9.36354650186033e-31
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0389514981882917 lu0=2.59573421087258e-09 wu0=-2.12673230412961e-08 pu0=8.7692829135559e-15
+  a0=1.1222
+  keta=-0.01066
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.62456389941005+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=7.41941319728576e-08 wnfactor=6.49894846236566e-07 pnfactor=-2.67975041317801e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=2.57198007896776 lpclm=-6.37463241841253e-07 wpclm=-1.08166468635668e-05 ppclm=4.4600929011357e-12
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=-5.48509237529169e-06 lalpha0=9.53943144965828e-12 walpha0=1.56212266196728e-10 palpha0=-6.44119409944943e-17
+  alpha1=0.0
+  beta0=32.43483696 lbeta0=1.86588762726144e-6
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.37073
+  kt2=-0.019151
+  at=9620.20799999998 lat=0.011866944314112
+  ute=-1.13989264 lute=-6.56469259929595e-8
+  ua1=2.0117e-9
+  ub1=-3.1137654372168e-18 lub1=7.28500993320229e-25 wub1=1.02558156798129e-23 pub1=-4.22884201415132e-30
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.02e-6
+  sbref=2.01e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.39 nmos
* DC IV MOS Parameters
+  lmin=5e-07 lmax=6e-07 wmin=5.0e-06 wmax=7.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={1.06091998096073+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-1.12719047461424e-07 wvth0=-5.35786409340352e-07 pvth0=2.20924024881761e-13
+  k1=0.88325
+  k2=-0.00404474018696965 lk2=-8.88792714306566e-09 wk2=3.48784287436979e-08 pk2=-1.43816317944614e-14
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=95442.0681148244 lvsat=2.19494226058048e-05 wvsat=-0.0452912971924393 pvsat=1.86752323191415e-8
+  ua=1.39044952457449e-10 lua=-9.0804366914895e-17 wua=-9.68435311517854e-17 pua=3.9932074261003e-23
+  ub=3.53389412817445e-19 lub=6.82527652836508e-25 wub=2.15966525943768e-24 pub=-8.90507734415496e-31
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0372932651526123 lu0=3.27948338787244e-09 wu0=4.42893821135138e-08 pu0=-1.82621066631579e-14
+  a0=1.1222
+  keta=-0.01066
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={2.5366658062886+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-7.14234319901815e-07 wnfactor=-8.7416333486928e-06 pnfactor=3.6044901284666e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.217674431999997 lpclm=3.33301731406847e-7
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=2.759165488e-05 lalpha0=-4.09930220659968e-12
+  alpha1=0.0
+  beta0=36.96
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.4331972 lkt1=2.57574753792e-8
+  kt2=-0.019151
+  at=108687.963508224 lat=-0.028982257721127 wat=-0.528627906440636 pat=2.17972316430106e-7
+  ute=-1.30066168 lute=6.43936884480031e-10
+  ua1=-1.088859472e-09 lua1=1.27847229044659e-15
+  ub1=5.54157048e-18 lub1=-2.84040559744128e-24
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=1.81e-6
+  sbref=1.81e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.40 nmos
* DC IV MOS Parameters
+  lmin=2.0e-05 lmax=1.0e-04 wmin=3.0e-06 wmax=5.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.800603584032+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} wvth0=-4.61281485296475e-9
+  k1=0.88325
+  k2=-0.0415250021296 wk2=1.26124069269229e-8
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=133679.035614 wvsat=-0.168170483603328
+  ua=3.988788169096e-10 wua=-1.65000994239883e-15
+  ub=1.21900881548e-18 wub=1.48611541677434e-24
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0454752482968 wu0=-1.69885115440121e-8
+  a0=0.62809289928104 wa0=1.01876625909821e-6
+  keta=-0.012053675709 wketa=-5.52248015044945e-8
+  a1=0.0
+  a2=0.65972622
+  ags=0.0982374824866999 wags=1.59155010100403e-7
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.92922630284+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} wnfactor=1.21693339213092e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-0.84355705864 wpclm=5.26649927357602e-6
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=5.023772131e-06 walpha0=2.85342050361868e-11
+  alpha1=0.0
+  beta0=21.577916335 wbeta0=6.71437688301655e-6
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.40273
+  kt2=-0.019151
+  at=210015.8336 wat=-0.291335674924109
+  ute=-1.2986
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.41 nmos
* DC IV MOS Parameters
+  lmin=8e-06 lmax=2.0e-05 wmin=3.0e-06 wmax=5.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.800603584032+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} wvth0=-4.6128148529639e-9
+  k1=0.88325
+  k2=-0.0415250021296 wk2=1.26124069269229e-8
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=133679.035614 wvsat=-0.168170483603328
+  ua=3.988788169096e-10 wua=-1.65000994239883e-15
+  ub=1.21900881548e-18 wub=1.48611541677433e-24
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0454752482968 wu0=-1.69885115440121e-8
+  a0=0.62809289928104 wa0=1.01876625909821e-6
+  keta=-0.012053675709 wketa=-5.52248015044945e-8
+  a1=0.0
+  a2=0.65972622
+  ags=0.0982374824866999 wags=1.59155010100403e-7
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.92922630284+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} wnfactor=1.2169333921309e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-0.843557058639999 wpclm=5.26649927357602e-6
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=5.023772131e-06 walpha0=2.85342050361868e-11
+  alpha1=0.0
+  beta0=21.577916335 wbeta0=6.71437688301655e-6
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.40273
+  kt2=-0.019151
+  at=210015.8336 wat=-0.291335674924109
+  ute=-1.2986
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.42 nmos
* DC IV MOS Parameters
+  lmin=4e-06 lmax=8e-06 wmin=3.0e-06 wmax=5.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.795107637565637+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=4.29361804332383e-08 wvth0=7.3977451010289e-09 pvth0=-9.38305299087451e-14
+  k1=0.88325
+  k2=-0.0457326257158378 lk2=3.28713692172148e-08 wk2=1.87861673656463e-08 pk2=-4.82314909308149e-14
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=138951.018099728 lvsat=-0.0411864985646198 wvsat=-0.207231919407947 pvsat=3.05161061148118e-7
+  ua=3.98819907918775e-10 lua=4.60216829742726e-19 wua=-1.64983712338444e-15 pua=-1.35012020759785e-24
+  ub=1.29805417145197e-18 lub=-6.1752888009264e-25 wub=1.54193812769837e-24 pub=-4.36105774169468e-31
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0456091522546432 lu0=-1.04610271040052e-09 wu0=-1.62509575913888e-08 pu0=-5.76201929602071e-15
+  a0=0.627032334241484 la0=8.28549043887326e-09 wa0=1.018360170569e-06 pa0=3.17250003592349e-15
+  keta=-0.012053675709 wketa=-5.52248015044944e-8
+  a1=0.0
+  a2=0.65972622
+  ags=0.0961443780564972 lags=1.63520350918329e-08 wags=1.82718412702498e-07 pags=-1.84085218430837e-13
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.97377557733188+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-3.48033900886795e-07 wnfactor=9.34927469069086e-08 pnfactor=2.20312502494935e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-0.843557058639999 wpclm=5.26649927357602e-6
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=-7.57888334665808e-06 lalpha0=9.84561790837055e-11 walpha0=6.82825783457007e-11 palpha0=-3.10527647747355e-16
+  alpha1=0.0
+  beta0=16.9091201014777 lbeta0=3.64742048918104e-05 wbeta0=1.24701900819202e-05 pbeta0=-4.496634666307e-11
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.414167008 lkt1=8.93497493306877e-8
+  kt2=-0.019151
+  at=305132.905418102 lat=-0.743086524379147 wat=-0.424384623240473 pat=1.03942308869407e-6
+  ute=-1.33672336 lute=2.97832497768961e-7
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.43 nmos
* DC IV MOS Parameters
+  lmin=2e-06 lmax=4e-06 wmin=3.0e-06 wmax=5.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.810651369602644+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-1.63217487857957e-08 wvth0=1.12095995533308e-09 pvth0=-6.99013159335446e-14
+  k1=0.88325
+  k2=-0.0390149644616333 lk2=7.2613873820058e-09 wk2=-8.88734868590747e-10 pk2=2.67758471532477e-14
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=145713.764705023 lvsat=-0.0669683609068664 wvsat=-0.218719656705276 pvsat=3.48956175605265e-7
+  ua=4.7360752173533e-10 lua=-2.84655295677206e-16 wua=-1.87802177486124e-15 pua=8.68566441264867e-22
+  ub=1.10824530861904e-18 lub=1.06086280804407e-25 wub=1.54407564479936e-24 pub=-4.44254707564163e-31
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0457703051846262 lu0=-1.66047182688017e-09 wu0=-2.02084882752738e-08 pu0=9.32541740125808e-15
+  a0=0.192076707329375 la0=1.66648248531847e-06 wa0=1.89322951360919e-06 pa0=-3.33212339173253e-12
+  keta=-0.0402460864895334 lketa=1.07478942545415e-07 wketa=2.99630220697904e-08 pketa=-3.24764606573895e-13
+  a1=0.0
+  a2=0.65972622
+  ags=0.0141066713072558 lags=3.29107337889409e-07 wags=4.82937954981692e-07 pags=-1.32862298736533e-12
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.888626290988336+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-2.34162111849963e-08 wnfactor=3.68256350963281e-07 pnfactor=-8.2717867673893e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-0.84355705864 wpclm=5.26649927357602e-6
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=2.16719321747202e-05 lalpha0=-1.30577579578037e-11 walpha0=-2.51057580736096e-11 palpha0=4.55000691640934e-17
+  alpha1=0.0
+  beta0=24.1296802120651 lbeta0=8.9470036420542e-06 wbeta0=-9.95387967169024e-07 pbeta0=6.36896129428254e-12
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.407041024 lkt1=6.21831039920643e-8
+  kt2=-0.019151
+  at=178277.30893272 lat=-0.25947036709645 wat=-0.220487087427825 pat=2.62097172604225e-7
+  ute=-1.22235328 lute=-1.38184675537921e-7
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.44 nmos
* DC IV MOS Parameters
+  lmin=1e-06 lmax=2e-06 wmin=3.0e-06 wmax=5.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.812865674091839+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-2.03348125265255e-08 wvth0=-7.23318332566585e-08 pvth0=6.32198255051045e-14
+  k1=0.88325
+  k2=-0.0458932436477358 lk2=1.97271403690301e-08 wk2=2.38080496805884e-08 pk2=-1.79830245694738e-14
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=122927.076973593 lvsat=-0.0256712264104361 wvsat=-0.07143022132696 pvsat=8.20182294494695e-8
+  ua=6.97672542114505e-10 lua=-6.90736398451119e-16 wua=-2.55475758734278e-15 pua=2.09503911671441e-21
+  ub=8.02770447445528e-19 lub=6.59709368804165e-25 wub=2.46759156163911e-24 pub=-2.11797585022585e-30
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0466223705966031 lu0=-3.20470064736071e-09 wu0=-2.18768713869848e-08 pu0=1.23490881764039e-14
+  a0=1.08398346090606 la0=5.00477671683128e-08 wa0=6.32740677883437e-08 pa0=-1.56292588753612e-14
+  keta=0.0431990129013204 lketa=-4.3751615104207e-08 wketa=-2.70461543008019e-07 pketa=2.19705648000962e-13
+  a1=0.0
+  a2=0.65972622
+  ags=0.2829424044518 lags=-1.58113339374842e-07 wags=-3.65399110077846e-07 pags=2.0884881577641e-13
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.02440339930684+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-2.69489952566511e-07 wnfactor=-5.68695112012374e-07 pnfactor=8.70892189864513e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-2.25939133038738 lpclm=2.56596742072156e-06 wpclm=9.54466622747567e-06 ppclm=-7.75347598456268e-12
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=-9.71393997733106e-06 lalpha0=4.38239880347563e-11 walpha0=6.24135599028203e-11 palpha0=-1.13114341500038e-16
+  alpha1=0.0
+  beta0=21.7989308027566 lbeta0=1.31711047035227e-05 wbeta0=1.44074302940239e-05 pbeta0=-2.15461207419347e-11
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.37273
+  kt2=-0.019151
+  at=31894.133146176 lat=0.00582513217583197 wat=-0.10052100459744 pat=4.4678321911736e-8
+  ute=-1.2986
+  ua1=3.0044e-9
+  ub1=-3.9962008e-18 lub1=4.41667733068801e-25
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.81e-6
+  sbref=2.81e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.45 nmos
* DC IV MOS Parameters
+  lmin=8.0e-07 lmax=1e-06 wmin=3.0e-06 wmax=5.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.78294720779271+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=3.96903471304207e-09 wvth0=2.23103670236201e-08 pvth0=-1.36614409017764e-14
+  k1=0.88325
+  k2=-0.0309003236939849 lk2=7.54785174547997e-09 wk2=6.78555637928356e-09 pk2=-4.155040451065e-15
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=89427.231845921 lvsat=0.00154190378119601 wvsat=0.119964445888062 pvsat=-7.34585489373118e-8
+  ua=-1.71058002975951e-10 lua=1.4964697625482e-17 wua=9.85877862136336e-17 pua=-6.03688506589116e-23
+  ub=1.52133277580138e-18 lub=7.59953212368886e-26 wub=-5.67311957050918e-25 pub=3.47385534532729e-31
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0453410727040071 lu0=-2.16385624248089e-09 wu0=-2.71114100930686e-08 pu0=1.66012924107492e-14
+  a0=1.21721548333449 la0=-5.81814010031106e-08 wa0=1.78852721277755e-07 pa0=-1.09517959936334e-13
+  keta=-0.01066
+  a1=0.0
+  a2=0.65972622
+  ags=-0.131979411560422 lags=1.78942588957263e-07 wags=-4.39890178538935e-07 pags=2.69360592365818e-13
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.40074519606403+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=2.37130057622938e-07 wnfactor=2.04460338676415e-06 pnfactor=-1.25198425943762e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=1.119647876 lpclm=-1.78947772038337e-7
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=0.000117653757726655 lalpha0=-5.96413780473092e-11 walpha0=-3.12067799514101e-10 palpha0=1.91090348083267e-16
+  alpha1=0.0
+  beta0=45.7612750205539 lbeta0=-6.29437014898585e-06 wbeta0=-4.92122322330426e-05 pbeta0=3.01344214366523e-11
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.37885336 lkt1=4.97422576896017e-9
+  kt2=-0.019151
+  at=69880.70359632 lat=-0.0250327265173562 wat=-0.184892544394649 pat=1.13216361064442e-7
+  ute=-1.45627652 lute=1.28086313550719e-7
+  ua1=6.043729736e-09 lua1=-2.4689569604233e-15
+  ub1=-1.017441844e-17 lub1=5.46045633787584e-24
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.41e-6
+  sbref=2.41e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.46 nmos
* DC IV MOS Parameters
+  lmin=6e-07 lmax=8.0e-07 wmin=3.0e-06 wmax=5.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.78036698621328+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=5.54899727410532e-09 wvth0=6.49286593277593e-08 pvth0=-3.97581555381244e-14
+  k1=0.88325
+  k2=-0.00116296238680283 lk2=-1.06614051279147e-08 wk2=-1.46938045224041e-08 pk2=8.99754548603088e-15
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=80211.664859556 lvsat=0.00718492720735892 wvsat=0.0221689686497801 pvsat=-1.35748575871317e-8
+  ua=-4.79846489531346e-10 lua=2.04047004328867e-16 wua=9.95798538099068e-16 pua=-6.09763293625431e-22
+  ub=1.49215513273606e-18 lub=9.38618424809303e-26 wub=-2.99069131859024e-24 pub=1.83130795926027e-30
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0303872409536685 lu0=6.99291327619449e-09 wu0=2.17394478150077e-08 pu0=-1.33118465172505e-14
+  a0=1.1222
+  keta=-0.01066
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.890879758743044+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-6.29969799496804e-08 wnfactor=-6.87452319309837e-07 pnfactor=4.20951803396908e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=1.22410309618793 lpclm=-2.42909463747335e-07 wpclm=-4.04806962997465e-06 ppclm=2.47877876494015e-12
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=2.74229956691121e-05 lalpha0=-4.38983413204146e-12 walpha0=-9.0408973961567e-12 palpha0=5.53606694797299e-18
+  alpha1=0.0
+  beta0=32.43483696 lbeta0=1.86588762726144e-6
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.37073
+  kt2=-0.019151
+  at=9620.20800000001 lat=0.011866944314112
+  ute=-1.13989264 lute=-6.56469259929586e-8
+  ua1=2.0117e-9
+  ub1=-1.58851322483152e-18 lub1=2.02997482040433e-25 wub1=2.5965207054706e-24 pub1=-1.58994310270505e-30
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.02e-6
+  sbref=2.01e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.47 nmos
* DC IV MOS Parameters
+  lmin=5e-07 lmax=6e-07 wmin=3.0e-06 wmax=5.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.953941810338902+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-6.60221514065579e-08 wvth0=1.42137698811066e-09 pvth0=-1.35718167673215e-14
+  k1=0.88325
+  k2=0.0294436810328514 lk2=-2.32816260490012e-08 wk2=-1.33288969582186e-07 pk2=5.78986014661211e-14
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=95903.4215643189 lvsat=0.000714651014743828 wvsat=-0.0476080564329213 pvsat=1.51967218273691e-8
+  ua=5.27703064967779e-10 lua=-2.11401948775085e-16 wua=-2.04855165110418e-15 pua=6.45531885989881e-22
+  ub=-3.34987023744358e-19 lub=8.47258330715442e-25 wub=5.61645629910973e-24 pub=-1.71772886083166e-30
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0509364529081776 lu0=-1.48026658428001e-09 wu0=-2.42220408247226e-08 pu0=5.63972986250127e-15
+  a0=1.1222
+  keta=-0.01066
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.22717705826796+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-2.01664463246586e-07 wnfactor=-2.16582870128498e-06 pnfactor=1.03053960723501e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-1.39456982277588 lpclm=8.36863652966527e-07 wpclm=8.09613925994931e-06 ppclm=-2.52871575189553e-12
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=2.39908929817757e-05 lalpha0=-2.97465463835588e-12 walpha0=1.80817947923133e-11 palpha0=-5.647595458252e-18
+  alpha1=0.0
+  beta0=36.96
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.4331972 lkt1=2.57574753792002e-8
+  kt2=-0.019151
+  at=3418.36799999996 lat=0.014424186212352
+  ute=-1.30066168 lute=6.43936884480031e-10
+  ua1=-1.088859472e-09 lua1=1.27847229044659e-15
+  ub1=6.57569932966304e-18 lub1=-3.16340126582964e-24 wub1=-5.19304141094121e-24 pub1=1.62197378212773e-30
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=1.81e-6
+  sbref=1.81e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.48 nmos
* DC IV MOS Parameters
+  lmin=2.0e-05 lmax=1.0e-04 wmin=1.5e-06 wmax=3.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.797280429121333+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} wvth0=5.42862276809016e-9
+  k1=0.88325
+  k2=-0.0397531907626667 wk2=7.25859893553785e-9
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=39317.0782346666 wvsat=0.116959079807594
+  ua=-1.46640386864267e-10 wua=-1.63747616189373e-18
+  ub=1.83044246318667e-18 wub=-3.61427956287696e-25
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0415518804350667 wu0=-5.13343565766268e-9
+  a0=0.803755902738373 wa0=4.87972739397332e-7
+  keta=-0.0352530708493333 wketa=1.48758364164549e-8
+  a1=0.0
+  a2=0.65972622
+  ags=0.1600428043108 wags=-2.75995350319634e-8
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.90327744384+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} wnfactor=2.00101916601312e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=1.36597135350667 wpclm=-1.40993992921425e-6
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.4467e-5
+  alpha1=0.0
+  beta0=20.8581278666667 wbeta0=8.88933146666373e-6
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.414903264 wkt1=3.67834405517118e-8
+  kt2=-0.019151
+  at=157829.525866667 wat=-0.13364650067122
+  ute=-1.415767666 wute=3.54040615310227e-7
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.49 nmos
* DC IV MOS Parameters
+  lmin=8e-06 lmax=2.0e-05 wmin=1.5e-06 wmax=3.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.797280429121333+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} wvth0=5.42862276809016e-9
+  k1=0.88325
+  k2=-0.0397531907626667 wk2=7.25859893553785e-9
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=39317.0782346666 wvsat=0.116959079807594
+  ua=-1.46640386864267e-10 wua=-1.63747616189373e-18
+  ub=1.83044246318667e-18 wub=-3.61427956287697e-25
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0415518804350667 wu0=-5.13343565766268e-9
+  a0=0.803755902738373 wa0=4.87972739397332e-7
+  keta=-0.0352530708493333 wketa=1.48758364164548e-8
+  a1=0.0
+  a2=0.65972622
+  ags=0.1600428043108 wags=-2.75995350319634e-8
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.90327744384+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} wnfactor=2.00101916601314e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=1.36597135350667 wpclm=-1.40993992921425e-6
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.4467e-5
+  alpha1=0.0
+  beta0=20.8581278666667 wbeta0=8.88933146666374e-6
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.414903264 wkt1=3.67834405517118e-8
+  kt2=-0.019151
+  at=157829.525866667 wat=-0.13364650067122
+  ute=-1.415767666 wute=3.54040615310228e-7
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.50 nmos
* DC IV MOS Parameters
+  lmin=4e-06 lmax=8e-06 wmin=1.5e-06 wmax=3.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.794216222018893+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=2.39386154578585e-08 wvth0=1.00912980191765e-08 pvth0=-3.64263857203738e-14
+  k1=0.88325
+  k2=-0.0441133501170805 lk2=3.40630298902239e-08 wk2=1.38932702984565e-08 pk2=-5.18322819366981e-14
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=23896.2064008263 lvsat=0.120473032178898 wvsat=0.140424372800532 pvsat=-1.83318753199278e-7
+  ua=-1.46643842736939e-10 lua=2.69984384863922e-20 wua=-1.63221750559547e-18 pua=-4.10823899102831e-26
+  ub=2.02688962529306e-18 lub=-1.53471123662162e-24 wub=-6.60353352084187e-25 pub=2.33530563089518e-30
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0423133243804478 lu0=-5.94865594648289e-09 wu0=-6.29209292870342e-09 pu0=9.05181991021329e-15
+  a0=0.801348733828036 la0=1.88056123363121e-08 wa0=4.91635627227098e-07 pa0=-2.86157104564461e-14
+  keta=-0.0352530708493333 wketa=1.48758364164549e-8
+  a1=0.0
+  a2=0.65972622
+  ags=0.171535308881291 lags=-8.97833071862135e-08 wags=-4.50871965516879e-08 pags=1.36619487646359e-13
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.9742188300776+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-5.5421794559391e-07 wnfactor=9.21533887017791e-08 pnfactor=8.43330170656537e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=1.36597135350667 wpclm=-1.40993992921425e-6
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.5578639042803e-05 lalpha0=-8.68449771309537e-12 walpha0=-1.69153444259351e-12 palpha0=1.32148354211133e-17
+  alpha1=0.0
+  beta0=15.2903330063408 lbeta0=4.34974842279387e-05 wbeta0=1.73616110582375e-05 pbeta0=-6.61882948553167e-11
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.437942415146176 lkt1=1.79989589908712e-07 wkt1=7.18411492064998e-08 pkt1=-2.7388259940131e-13
+  kt2=-0.019151
+  at=260737.734319586 lat=-0.803953501592247 wat=-0.290237599329273 pat=1.22334227732586e-6
+  ute=-1.49256483648725 lute=5.99965299695709e-07 wute=4.70899644159522e-07 pute=-9.12941998004367e-13
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.51 nmos
* DC IV MOS Parameters
+  lmin=2e-06 lmax=4e-06 wmin=1.5e-06 wmax=3.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.81704241398592+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-6.30824979209516e-08 wvth0=-1.8190590433747e-08 pvth0=7.13936757766938e-14
+  k1=0.88325
+  k2=-0.0406034332735292 lk2=2.06820475505467e-08 wk2=3.91107462462475e-09 pk2=-1.37767980103052e-14
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=25218.6312424859 lvsat=0.115431504347744 wvsat=0.145375427282869 pvsat=-2.02193836440252e-7
+  ua=-1.47558768818895e-10 lua=3.51500407806814e-18 wua=-1.06968367774112e-18 pua=-2.18565035305715e-24
+  ub=1.63111040662524e-18 lub=-2.58678732424156e-26 wub=-3.58438615118643e-26 pub=-4.55343823553526e-32
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0406682670858836 lu0=3.22855199646697e-10 wu0=-4.79187403790361e-09 pu0=3.33248142493715e-15
+  a0=0.507267793715319 la0=1.13994096724187e-06 wa0=9.4082984590241e-07 pa0=-1.74109500130421e-12
+  keta=-0.0273162503099861 lketa=-3.0257826667693e-08 wketa=-9.10652086082813e-09 pketa=9.1428804013048e-14
+  a1=0.0
+  a2=0.65972622
+  ags=0.205055733539886 lags=-2.17574428847461e-07 wags=-9.40448065060311e-08 pags=3.2326234654926e-13
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.919468989584295+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-3.45493157687022e-07 wnfactor=2.75060264009216e-07 pnfactor=1.46027705274488e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=1.36597135350667 wpclm=-1.40993992921425e-6
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.11801475150397e-05 lalpha0=8.08402988389149e-12 walpha0=6.59682697759108e-12 palpha0=-1.83831832020676e-17
+  alpha1=0.0
+  beta0=22.8157436604076 lbeta0=1.48080902766564e-05 wbeta0=2.97487892563934e-06 pbeta0=-1.13412380238561e-11
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.407041024 lkt1=6.21831039920643e-8
+  kt2=-0.019151
+  at=95164.0133333333 lat=-0.1727308444224 wat=0.0306528671264267
+  ute=-1.27283664657477 lute=-2.37712388922502e-07 wute=1.52543468477576e-07 pute=3.00738711370229e-13
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.52 nmos
* DC IV MOS Parameters
+  lmin=1e-06 lmax=2e-06 wmin=1.5e-06 wmax=3.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.777582191977712+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=8.43268299251421e-09 wvth0=3.42827827413472e-08 pvth0=-2.37057074699652e-14
+  k1=0.88325
+  k2=-0.0363564649941381 lk2=1.29851140469483e-08 wk2=-5.00883383228424e-09 pk2=2.38907320285538e-15
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=80698.3013691131 lvsat=0.0148837009091332 wvsat=0.0561706963085202 pvsat=-4.05248911251254e-8
+  ua=-1.47823012066296e-10 lua=3.99390162808943e-18 wua=4.08179120694292e-20 pua=-4.19825236232797e-24
+  ub=1.63469588734106e-18 lub=-3.23659690209981e-26 wub=-4.62025992247443e-26 pub=-2.67608690837427e-32
+  uc=6.6204e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0408239367287185 lu0=4.07295018298211e-11 wu0=-4.35598730262046e-09 pu0=2.54250820266098e-15
+  a0=1.11954721766702 la0=3.02849251549391e-08 wa0=-4.41874423384527e-08 pa0=4.40872907970831e-14
+  keta=-0.0711045487294919 lketa=4.91012829367205e-08 wketa=7.49247284222181e-08 pketa=-6.0864054187591e-14
+  a1=0.0
+  a2=0.65972622
+  ags=0.104996123812249 lags=-3.62327959921153e-08 wags=1.72293692386896e-07 pags=-1.59432503180352e-13
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.732923050326026+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-7.40923631544965e-09 wnfactor=3.12058816328279e-07 pnfactor=7.89738969587641e-14
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=1.95675182758835 lpclm=-1.07069272127529e-06 wpclm=-3.19507647496695e-06 ppclm=3.23526722678326e-12
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=2.04604740457748e-05 lalpha0=-8.73503997951475e-12 walpha0=-2.87631996254097e-11 palpha0=4.57010659715084e-17
+  alpha1=0.0
+  beta0=29.7548150782496 lbeta0=2.23216133953027e-06 wbeta0=-9.63253107409359e-06 pbeta0=1.15076249854198e-11
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.37273
+  kt2=-0.019151
+  at=-19757.74115392 lat=0.0355459884180108 wat=0.0555532945964396 pat=-4.51279411192934e-8
+  ute=-1.48962053602923 lute=1.55172858155839e-07 wute=5.77198730857006e-07 pute=-4.68879308229458e-13
+  ua1=3.0044e-9
+  ub1=-4.2434203146176e-18 lub1=8.89712559312803e-25 wub1=7.47012824100389e-25 pub1=-1.3538382335788e-30
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.81e-6
+  sbref=2.81e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.53 nmos
* DC IV MOS Parameters
+  lmin=8.0e-07 lmax=1e-06 wmin=1.5e-06 wmax=3.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.771743538153427+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=1.31756316855194e-08 wvth0=5.61640250185202e-08 pvth0=-4.14806282964334e-14
+  k1=0.88325
+  k2=-0.0265649295913923 lk2=5.03109734402334e-09 wk2=-6.31452189396836e-09 pk2=3.44973062013162e-15
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=135887.584061388 lvsat=-0.0299485402359789 wvsat=-0.020422849066623 pvsat=2.1694803150737e-8
+  ua=-1.24453426036967e-10 lua=-1.49900544086318e-17 wua=-4.2235306530664e-17 pua=3.01441654629845e-23
+  ub=1.37782221698547e-18 lub=1.76301760860978e-25 wub=-1.33672128920369e-25 pub=4.42937787910834e-32
+  uc=6.49709630289469e-11 luc=1.00164032091741e-18 wuc=3.72581602787839e-18 puc=-3.0266144888226e-24
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0356684797366112 lu0=4.22869281297034e-09 wu0=2.11585782760664e-09 pu0=-2.71480458304729e-15
+  a0=1.26284987282847 la0=-8.61249805282931e-08 wa0=4.0961203188171e-08 pa0=-2.50820193154316e-14
+  keta=-0.01066
+  a1=0.0
+  a2=0.65972622
+  ags=-0.245337543794839 lags=2.48355854217157e-07 wags=-9.73606714077506e-08 pags=5.96174440871364e-14
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.38080862255111+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-5.33710010514488e-07 wnfactor=-9.16813106387955e-07 pnfactor=1.07723079917038e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.683360119059578 lpclm=-3.62707943358703e-08 wpclm=1.31831239106108e-06 ppclm=-4.3112103109048e-13
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.51850123805024e-05 lalpha0=-4.44959255219404e-12 walpha0=-2.44229538893578e-12 palpha0=2.43196479076682e-17
+  alpha1=0.0
+  beta0=27.9713146054231 lbeta0=3.68096297962428e-06 wbeta0=4.54294397502088e-06 pbeta0=-7.62371407763502e-15
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.37885336 lkt1=4.97422576895996e-9
+  kt2=-0.019151
+  at=8691.59999999998 lat=0.0124355644224
+  ute=-1.45627652 lute=1.2808631355072e-7
+  ua1=6.043729736e-09 lua1=-2.46895696042329e-15
+  ub1=-1.06285443420936e-17 lub1=6.07657867129658e-24 wub1=1.37221316506844e-24 pub1=-1.86171097775943e-30
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.41e-6
+  sbref=2.41e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.54 nmos
* DC IV MOS Parameters
+  lmin=6e-07 lmax=8.0e-07 wmin=1.5e-06 wmax=3.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.791257381070887+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=1.22660316881338e-09 wvth0=3.20216105831145e-08 pvth0=-2.66973588107159e-14
+  k1=0.88325
+  k2=0.0065665611906177 lk2=-1.52565071954695e-08 wk2=-3.80497812763055e-08 pk2=2.28823724092744e-14
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=69009.0981801694 lvsat=0.0110035642945832 wvsat=0.056019293877082 pvsat=-2.51134728908396e-8
+  ua=-1.55742748206169e-10 lua=4.1695239711692e-18 wua=1.64678752939168e-17 pua=-5.801906082752e-24
+  ub=-3.870775488576e-19 lub=1.25701342387826e-24 wub=2.68770714760872e-24 pub=-1.68333832188163e-30
+  uc=5.30374181086835e-11 luc=8.30897948321181e-18 wuc=3.97849075045517e-17 puc=-2.51068943272829e-23
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0368950144749426 lu0=3.4776414374394e-09 wu0=2.07518189226119e-09 pu0=-2.68989724350152e-15
+  a0=1.1222
+  keta=-0.01066
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.500303222503197+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=5.45514412925311e-09 wnfactor=4.92736396031588e-07 pnfactor=2.14112895056806e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.229324232153652 lpclm=2.41751724508558e-07 wpclm=-1.04218811723455e-06 ppclm=1.01429840815723e-12
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=-1.03102919696392e-05 lalpha0=1.11621001323542e-11 walpha0=1.04976193063777e-10 palpha0=-4.14565596375124e-17
+  alpha1=0.0
+  beta0=27.8443365992531 lbeta0=3.75871618401037e-06 wbeta0=1.38709221390537e-05 pbeta0=-5.71948055112885e-12
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.37073
+  kt2=-0.019151
+  at=9620.20799999998 lat=0.011866944314112
+  ute=-1.13989264 lute=-6.56469259929595e-8
+  ua1=2.0117e-9
+  ub1=3.58258267435095e-19 lub1=-6.5103609141181e-25 wub1=-3.28595694830875e-24 pub1=9.90654276785512e-31
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.02e-6
+  sbref=2.01e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.55 nmos
* DC IV MOS Parameters
+  lmin=5e-07 lmax=6e-07 wmin=1.5e-06 wmax=3.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.961142370368162+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-6.88230937780674e-08 wvth0=-2.03362528287746e-08 pvth0=-5.10832684291116e-15
+  k1=0.88325
+  k2=-0.015317189549187 lk2=-6.23304895042141e-09 wk2=1.96307309899473e-09 pk2=6.3836320875806e-15
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=89362.7898897667 lvsat=0.00261100446981466 wvsat=-0.0278445044084579 pvsat=9.46659023902673e-9
+  ua=-1.44294085900614e-10 lua=-5.51171649254253e-19 wua=-1.80060842054948e-17 pua=8.41294848139722e-24
+  ub=3.1918427981612e-18 lub=-2.18704276330081e-25 wub=-5.04041724688976e-24 pub=1.50324557844829e-30
+  uc=9.50032377247392e-11 luc=-8.99503871399415e-18 wuc=-8.702144706486e-17 puc=2.71799306904501e-23
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0460179242459859 lu0=-2.84062685913455e-10 wu0=-9.35992934438145e-09 pu0=2.0252107833708e-15
+  a0=1.1222
+  keta=-0.01066
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={-0.190813510164692+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=2.90427453210599e-07 wnfactor=2.11885384374408e-06 pnfactor=-4.56393868863172e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-0.649789317021334 lpclm=6.04241888921176e-07 wpclm=5.84566728649205e-06 ppclm=-1.82581233759378e-12
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=2.39223067076111e-05 lalpha0=-2.95323267582841e-12 walpha0=1.8289039056333e-11 palpha0=-5.71232530269882e-18
+  alpha1=0.0
+  beta0=36.96
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.4331972 lkt1=2.57574753792e-8
+  kt2=-0.019151
+  at=3418.36800000002 lat=0.014424186212352
+  ute=-1.30066168 lute=6.43936884480031e-10
+  ua1=-1.088859472e-09 lua1=1.27847229044659e-15
+  ub1=5.42891186470908e-18 lub1=-2.74184911309738e-24 wub1=-1.72784189316335e-24 pub1=3.48187347407076e-31
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=1.81e-6
+  sbref=1.81e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.56 nmos
* DC IV MOS Parameters
+  lmin=2.0e-05 lmax=1.0e-04 wmin=1e-06 wmax=1.5e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.795429125968+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} wvth0=8.24567302178501e-9
+  k1=0.88325
+  k2=-0.027755791308 wk2=-1.09973399238513e-8
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=124925.39248 wvsat=-0.0133074964303319
+  ua=-1.45640490944e-10 wua=-3.15897578813488e-18
+  ub=1.34704778572e-18 wub=3.74133421836875e-25
+  uc=9.3907278328e-11 wuc=-4.21549150940279e-17
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.03808569691888 wu0=1.40910219210928e-10
+  a0=1.1221892700996 wa0=3.42605848518229e-9
+  keta=-0.032912626924 wketa=1.131448119392e-8
+  a1=0.0
+  a2=0.65972622
+  ags=0.146725182444 wags=-7.33466917737219e-9
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.76777989828+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} wnfactor=4.06282840783052e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-0.76291756756 wpclm=1.82950092863822e-6
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=-1.8937129968e-05 walpha0=5.0829661598847e-11
+  alpha1=0.0
+  beta0=26.156477944 wbeta0=8.27054684688863e-7
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.386643368 wkt1=-6.21845627585605e-9
+  kt2=-0.019151
+  at=-93465.28 wat=0.24873825103424
+  ute=-1.2125237504 wute=4.47728851861624e-8
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.57 nmos
* DC IV MOS Parameters
+  lmin=8e-06 lmax=2.0e-05 wmin=1e-06 wmax=1.5e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.795429125968+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} wvth0=8.24567302178501e-9
+  k1=0.88325
+  k2=-0.027755791308 wk2=-1.09973399238513e-8
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=124925.39248 wvsat=-0.0133074964303319
+  ua=-1.45640490944e-10 wua=-3.15897578813478e-18
+  ub=1.34704778572e-18 wub=3.74133421836874e-25
+  uc=9.3907278328e-11 wuc=-4.21549150940278e-17
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.03808569691888 wu0=1.40910219210901e-10
+  a0=1.1221892700996 wa0=3.42605848518314e-9
+  keta=-0.032912626924 wketa=1.131448119392e-8
+  a1=0.0
+  a2=0.65972622
+  ags=0.146725182444 wags=-7.33466917737219e-9
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.76777989828+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} wnfactor=4.06282840783053e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-0.762917567560001 wpclm=1.82950092863821e-6
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=-1.8937129968e-05 walpha0=5.0829661598847e-11
+  alpha1=0.0
+  beta0=26.156477944 wbeta0=8.27054684688836e-7
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.386643368 wkt1=-6.21845627585541e-9
+  kt2=-0.019151
+  at=-93465.2800000001 wat=0.24873825103424
+  ute=-1.2125237504 wute=4.47728851861632e-8
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.58 nmos
* DC IV MOS Parameters
+  lmin=4e-06 lmax=8e-06 wmin=1e-06 wmax=1.5e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.78929854774396+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=4.78941369604878e-08 wvth0=1.75743164210212e-08 pvth0=-7.28784966590243e-14
+  k1=0.88325
+  k2=-0.0242114290564899 lk2=-2.76897488145132e-08 wk2=-1.63906470987596e-08 pk2=4.21343278015945e-14
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=124925.39248 wvsat=-0.0133074964303318
+  ua=-1.44900654010292e-10 lua=-5.77985471133715e-18 wua=-4.28475457700714e-18 pua=8.79496216034383e-24
+  ub=8.53407706866828e-19 lub=3.85648215906748e-24 wub=1.12528479694444e-24 pub=-5.86824692920231e-30
+  uc=9.3907278328e-11 wuc=-4.21549150940278e-17
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0368221512507345 lu0=9.87124331089696e-09 wu0=2.06359459350981e-09 pu0=-1.50206563539729e-14
+  a0=1.12897146569142 la0=-5.29847907810019e-08 wa0=-6.89412369467189e-09 pa0=8.06247307702334e-14
+  keta=-0.032912626924 wketa=1.131448119392e-8
+  a1=0.0
+  a2=0.65972622
+  ags=0.087764132154594 lags=4.60623535773739e-07 wags=8.2383884683905e-08 pags=-7.00911488198395e-13
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.5312229297685+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.84806252115326e-06 wnfactor=7.66241644374325e-07 pnfactor=-2.81211911981302e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-0.76291756756 wpclm=1.82950092863822e-6
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=-3.66862055505621e-05 lalpha0=1.3866174214037e-10 walpha0=7.78376844516571e-11 palpha0=-2.10995749221832e-16
+  alpha1=0.0
+  beta0=28.3454137520754 lbeta0=-1.7100702015117e-05 wbeta0=-2.50375699915563e-06 pbeta0=2.60214200269188e-11
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.382748464426912 lkt1=-3.0428295400564e-08 wkt1=-1.21451674570737e-08 pkt1=4.63014591226308e-14
+  kt2=-0.019151
+  at=-307684.97651984 lat=1.67355624703102 wat=0.574707366001227 pat=-2.54658025174473e-6
+  ute=-1.2125237504 wute=4.47728851861641e-8
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.59 nmos
* DC IV MOS Parameters
+  lmin=2e-06 lmax=4e-06 wmin=1e-06 wmax=1.5e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.80634770595522+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-1.71029826579983e-08 wvth0=-1.91690240116967e-09 pvth0=1.42857854069805e-15
+  k1=0.88325
+  k2=-0.0345414522041578 lk2=1.16917703121742e-08 wk2=-5.31318736543281e-09 pk2=-9.66707283178637e-17
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=135334.041735227 lvsat=-0.039681268267076 wvsat=-0.0221825680166952 pvsat=3.38347549112699e-8
+  ua=-1.45555522057482e-10 lua=-3.2832776797835e-18 wua=-4.11794013821911e-18 pua=8.15900947003216e-24
+  ub=2.21601301411591e-18 lub=-1.33822710754926e-24 wub=-9.258655934209e-25 pub=1.95142754540153e-30
+  uc=1.18276022377411e-10 luc=-9.29018402143561e-17 wuc=-7.92358094267668e-17 puc=1.41364828376897e-22
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0412851738234057 lu0=-7.14329831171008e-09 wu0=-5.73059511030802e-09 pu0=1.46934136447212e-14
+  a0=1.11805048617408 la0=-1.13503474117893e-08 wa0=1.14274756609977e-08 pa0=1.07766379690386e-14
+  keta=-0.0567230885420418 lketa=9.0773480003079e-08 wketa=3.56406297896853e-08 pketa=-9.27394520329857e-14
+  a1=0.0
+  a2=0.65972622
+  ags=0.223599899597389 lags=-5.72280505360598e-08 wags=-1.2226268514076e-07 pags=7.92699972206898e-14
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.23082009283674+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-8.19036929109666e-07 wnfactor=-1.98709633063696e-07 pnfactor=8.66599373409925e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-0.76291756756 wpclm=1.82950092863821e-6
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=-9.44594004483783e-06 lalpha0=3.48126973033397e-11 walpha0=3.79826781217793e-11 palpha0=-5.90550738102103e-17
+  alpha1=0.0
+  beta0=20.7251755779197 lbeta0=1.19502063047913e-05 wbeta0=6.15600857290169e-06 pbeta0=-6.99251601499577e-12
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.407041024 lkt1=6.21831039920647e-8
+  kt2=-0.019151
+  at=232155.50719264 lat=-0.384497063283481 wat=-0.177801335436538 pat=3.22235761059714e-7
+  ute=-1.18053378575218 lute=-1.21956493865615e-07 wute=1.20900818839993e-08 pute=1.24597827609757e-13
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.60 nmos
* DC IV MOS Parameters
+  lmin=1e-06 lmax=2e-06 wmin=1e-06 wmax=1.5e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.814288702581149+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-3.14947367190467e-08 wvth0=-2.15719727704564e-08 pvth0=3.70501701534892e-14
+  k1=0.88325
+  k2=-0.0360973284903804 lk2=1.45115409172419e-08 wk2=-5.40315096631917e-09 pk2=6.63735442581699e-17
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=129183.402395662 lvsat=-0.0285342431689657 wvsat=-0.0176070455493361 pvsat=2.55423708248665e-8
+  ua=-3.69141694944644e-12 lua=-2.60388702474861e-16 wua=-2.19278176850246e-16 pua=3.98101652231759e-22
+  ub=1.23259449596298e-18 lub=4.4405767596596e-25 wub=5.65658199776845e-25 pub=-7.51714719867304e-31
+  uc=3.47076980308303e-11 luc=5.8552042458629e-17 wuc=4.79265998618029e-17 puc=-8.90961838235125e-23
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.036324604785805 lu0=1.84691953561906e-09 wu0=2.49045714296943e-09 pu0=-2.05895311774636e-16
+  a0=0.00555375737445463 la0=2.00486752407401e-06 wa0=1.65092961846341e-06 pa0=-2.96055211750891e-12
+  keta=-0.00336831363285089 lketa=-5.92329933674445e-09 wketa=-2.81466556024665e-08 pketa=2.28645416254852e-14
+  a1=0.0
+  a2=0.65972622
+  ags=-0.389758852887688 lags=1.05438409750774e-06 wags=9.2514156072217e-07 pags=-1.81897842410955e-12
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.708469457199696+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.27637932478234e-07 wnfactor=3.49268821937707e-07 pnfactor=-1.26521707813495e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-2.53525898980504 lpclm=3.21207816382588e-06 wpclm=3.64022772140623e-06 ppclm=-3.28164535269802e-12
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=-2.9503199336359e-06 lalpha0=2.30404511334844e-11 walpha0=6.86002231971246e-12 palpha0=-2.65036428451569e-18
+  alpha1=0.0
+  beta0=20.6878821589759 lbeta0=1.20177945105061e-05 wbeta0=4.16423993798254e-06 pbeta0=-3.382762014261e-12
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.37273
+  kt2=-0.019151
+  at=16750.656 lat=0.005888903107584
+  ute=-0.861662112825202 lute=-6.99859106091399e-07 wute=-3.78339227478783e-07 pute=8.32186920423067e-13
+  ua1=3.0044e-9
+  ub1=-3.00506542647695e-18 lub1=-1.35460258524047e-24 wub1=-1.13733979827794e-24 pub1=2.06124186065185e-30
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.81e-6
+  sbref=2.81e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.61 nmos
* DC IV MOS Parameters
+  lmin=8.0e-07 lmax=1e-06 wmin=1e-06 wmax=1.5e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.744491438544566+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=2.52040935593752e-08 wvth0=9.76324004051387e-08 pvth0=-5.9783833534481e-14
+  k1=0.88325
+  k2=-0.0165104491485989 lk2=-1.39958629974358e-09 wk2=-2.16140024955885e-08 pk2=1.32350318321387e-14
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=85534.2731175842 lvsat=0.00692351591227114 wvsat=0.0561976693575044 pvsat=-3.44118560636968e-8
+  ua=-8.75020098929532e-10 lua=4.47422953730114e-16 wua=1.09987047580969e-15 pua=-6.73490287675403e-22
+  ub=2.2501462697927e-18 lub=-3.82536261779784e-25 wub=-1.46105100246691e-24 pub=8.94654126646577e-31
+  uc=2.32251799471008e-10 luc=-1.01920142728879e-16 wuc=-2.50818406990875e-16 puc=1.53585140063164e-22
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0310878804285038 lu0=6.10089925313163e-09 wu0=9.08596340958284e-09 pu0=-5.56366249037032e-15
+  a0=6.61107790962271 la0=-3.36103754366674e-06 wa0=-8.09721277482409e-06 pa0=4.95821488168469e-12
+  keta=-0.01066
+  a1=0.0
+  a2=0.65972622
+  ags=3.19821052994181 lags=-1.86025259906245e-06 wags=-5.33726314619372e-06 pags=3.26819836588768e-12
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.261751149710028+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=4.9052329551116e-07 wnfactor=7.86009649620466e-07 pnfactor=-4.81302004809997e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=2.61618538141808 lpclm=-9.72625550916022e-07 wpclm=-1.62278663200883e-06 ppclm=9.93690675097761e-13
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=3.97770467937183e-06 lalpha0=1.74125673314521e-11 walpha0=1.46113940329511e-11 palpha0=-8.9470825765612e-18
+  alpha1=0.0
+  beta0=30.95683696 lbeta0=3.6759528432614e-6
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.378853360000001 lkt1=4.97422576896017e-9
+  kt2=-0.019151
+  at=8691.59999999998 lat=0.0124355644224
+  ute=-3.18087017287686 lute=1.18411709257873e-06 wute=2.6242417286493e-06 pute=-1.6069176831542e-12
+  ua1=6.043729736e-09 lua1=-2.4689569604233e-15
+  ub1=-1.34639290516153e-17 lub1=7.14150885654988e-24 wub1=5.68669899138971e-24 pub1=-3.48217051359161e-30
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.41e-6
+  sbref=2.41e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.62 nmos
* DC IV MOS Parameters
+  lmin=6e-07 lmax=8.0e-07 wmin=1e-06 wmax=1.5e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.81230127568+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-1.63183108727881e-8
+  k1=0.88325
+  k2=-0.01843891394 lk2=-2.18717883236157e-10
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=105823.73976 lvsat=-0.00550045493367934
+  ua=-1.449204246e-10 lua=3.56639549865696e-19
+  ub=1.3792241744e-18 lub=1.50760690424602e-25
+  uc=7.91831798399999e-11 luc=-8.19071645850625e-18
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0382587781408 lu0=1.70990043157511e-9
+  a0=1.1222
+  keta=-0.01066
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.824118689599999+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.46165405605094e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-0.45557876 lpclm=9.08326216383361e-7
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=5.867774152e-05 lalpha0=-1.60822344273907e-11
+  alpha1=0.0
+  beta0=36.96
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.37073
+  kt2=-0.019151
+  at=9620.20800000001 lat=0.011866944314112
+  ute=-1.13989264 lute=-6.56469259929595e-8
+  ua1=2.0117e-9
+  ub1=-1.8012e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.02e-6
+  sbref=2.01e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.63 nmos
* DC IV MOS Parameters
+  lmin=5e-07 lmax=6e-07 wmin=1e-06 wmax=1.5e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.950202998915469+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-7.31801558248086e-08 wvth0=-3.6902707428133e-09 pvth0=1.52163147700909e-15
+  k1=0.88325
+  k2=0.00770173311985431 lk2=-1.09974477293082e-08 wk2=-3.30638547317334e-08 pk2=1.3633417604664e-14
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=89527.1562788717 lvsat=0.00121921311259515 wvsat=-0.0280946138393705 pvsat=1.15844206920706e-8
+  ua=-1.13147630210777e-10 lua=-1.27444273974089e-17 wua=-6.54003376775803e-17 pua=2.69669136366229e-23
+  ub=-1.40530690085229e-18 lub=1.29892309586983e-24 wub=1.95487236981171e-24 pub=-8.0606425347868e-31
+  uc=-8.89384632420158e-11 luc=6.11318893633597e-17 wuc=1.9287491374481e-16 puc=-7.952927043388e-23
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0415012187257568 lu0=3.72925450536367e-10 wu0=-2.48704825588061e-09 pu0=1.02549952963682e-15
+  a0=1.1222
+  keta=-0.01066
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.82274775225848+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-2.65605307575255e-07 wnfactor=-9.45097759712248e-07 pnfactor=3.8969782984871e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=3.191854 lpclm=-5.95641618144e-7
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=3.594145888e-05 lalpha0=-6.70724658874369e-12
+  alpha1=0.0
+  beta0=36.96
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.4331972 lkt1=2.57574753792e-8
+  kt2=-0.019151
+  at=-52130.6597631592 lat=0.037329050124102 wat=0.0845266224880332 pat=-3.48533694102257e-8
+  ute=-0.306344294257789 lute=-4.0934891668292e-07 wute=-1.51301100455372e-06 pute=6.23868905573663e-13
+  ua1=-1.088859472e-09 lua1=1.27847229044659e-15
+  ub1=1.70133994124339e-17 lub1=-7.75793666332534e-24 wub1=-1.93554700460592e-23 pub1=7.98095709691185e-30
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=1.81e-6
+  sbref=1.81e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.64 nmos
* DC IV MOS Parameters
+  lmin=2.0e-05 lmax=1.0e-04 wmin=7.5e-07 wmax=1.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.820109166792+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} wvth0=-1.69688881263809e-8
+  k1=0.88325
+  k2=-0.029358876224 wk2=-9.3595353947406e-9
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=145544.2888 wvsat=-0.0343729568068303
+  ua=-1.53513692968e-10 wua=4.88474404530103e-18
+  ub=2.41014977296e-18 wub=-7.11993228242768e-25
+  uc=3.9200631008e-11 wuc=1.37365687936287e-17
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.03963334656704 wu0=-1.44025842502898e-9
+  a0=2.1057418918264 wa0=-1.00142834592298e-6
+  keta=-0.026727225088 wketa=4.9951159249559e-9
+  a1=0.0
+  a2=0.65972622
+  ags=0.0756403710719999 wags=6.52896970393226e-8
+  b0=-4.600021304e-07 wb0=5.03611119454203e-13
+  b1=4.957130992e-10 wb1=-5.06449253502473e-16
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.21532997312+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} wnfactor=-5.09602735778334e-8
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=3.56572142936 wpclm=-2.59288773167708e-6
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=3.9300151368e-05 walpha0=-8.66892277632815e-12
+  alpha1=0.0
+  beta0=21.53352768 wbeta0=5.55012880550654e-6
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.398903264 wkt1=6.30696455171185e-9
+  kt2=-0.019151
+  at=427796.88 wat=-0.28381340482704
+  ute=-1.279818752 wute=1.13525361930816e-7
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.65 nmos
* DC IV MOS Parameters
+  lmin=8e-06 lmax=2.0e-05 wmin=7.5e-07 wmax=1.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.830922199430262+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-2.14231435808209e-07 wvth0=-2.80161094255225e-08 pvth0=2.18871260244948e-13
+  k1=0.88325
+  k2=-0.0233947281343583 lk2=-1.1816370590574e-07 wk2=-1.54528550037078e-08 pk2=1.20722895448247e-13
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=167447.662848886 lvsat=-0.433957006190218 wvsat=-0.0567507141308676 pvsat=4.43355647030286e-7
+  ua=-1.56626383463571e-10 lua=6.16696699622618e-17 wua=8.06484919162513e-18 pua=-6.30053116743039e-23
+  ub=2.8638510383506e-18 lub=-8.98888191354379e-24 wub=-1.1755207556392e-24 pub=9.18356311802733e-30
+  uc=3.04473193238762e-11 luc=1.73423552198586e-16 wuc=2.26794597022073e-17 puc=-1.77179559492103e-22
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0405511180345269 lu0=-1.81831966850639e-08 wu0=-2.37790698695869e-09 pu0=1.85770083588691e-14
+  a0=2.74387901128276 la0=-1.26429870247415e-05 wa0=-1.65338623911252e-06 pa0=1.29168088377234e-11
+  keta=-0.0299102475185905 lketa=6.30631098903949e-08 wketa=8.24707625534809e-09 pketa=-6.44289307244011e-14
+  a1=0.0
+  a2=0.65972622
+  ags=0.0340360172822619 lags=8.24279436345164e-07 wags=1.07795117923439e-07 pags=-8.42131680377527e-13
+  b0=-7.80916702474051e-07 lb0=6.35806732922732e-12 wb0=8.31476059330234e-13 pb0=-6.49577035144373e-18
+  b1=8.18436206745978e-10 lb1=-6.39389864166505e-15 wb1=-8.36161898111682e-16 pb1=6.53237769844623e-21
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.24780323226037+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-6.43371121104036e-07 wnfactor=-8.41368385646633e-08 pnfactor=6.57305252844908e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=5.21797934167338 lpclm=-3.27350889174113e-05 wpclm=-4.28093024585535e-06 ppclm=3.34440654731846e-11
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=4.48242224928063e-05 lalpha0=-1.09444753212561e-10 walpha0=-1.43126342335555e-11 palpha0=1.11815107677638e-16
+  alpha1=0.0
+  beta0=17.996836090455 lbeta0=7.00701221004387e-05 wbeta0=9.16341806149788e-06 pbeta0=-7.158770080489e-11
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.402922231715392 lkt1=7.96251387504987e-08 wkt1=1.04129750698837e-08 pkt1=-8.13496600055541e-14
+  kt2=-0.019151
+  at=608650.42719264 lat=-3.58313124377244 wat=-0.468583878144778 pat=3.66073470025007e-6
+  ute=-1.35216017087706 lute=1.43325249750898e-06 wute=1.87433551257912e-07 pute=-1.46429388010003e-12
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.66 nmos
* DC IV MOS Parameters
+  lmin=4e-06 lmax=8e-06 wmin=7.5e-07 wmax=1.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.799931225325294+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=2.78804668670901e-08 wvth0=6.71135630863041e-09 pvth0=-5.24313704987396e-14
+  k1=0.88325
+  k2=-0.0543400449959453 lk2=1.23591507043443e-07 wk2=1.43904944047125e-08 pk2=-1.12423377495734e-13
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=79834.1666533409 lvsat=0.250509064224106 wvsat=0.0327603151652811 pvsat=-2.55934589537072e-7
+  ua=-1.45655295348703e-10 lua=-2.40401566766957e-17 wua=-3.51376921648919e-18 pua=2.74507457456691e-23
+  ub=2.03632613449454e-18 lub=-2.52397931625252e-24 wub=-8.32532779888331e-26 pub=6.50402580750174e-31
+  uc=6.54605660603713e-11 luc=-1.00111695757817e-16 wuc=-1.30921039321069e-17 puc=1.0227991486454e-22
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0394071235008702 lu0=-9.24592700597444e-09 wu0=-5.77362985619325e-10 pu0=4.51055363762122e-15
+  a0=0.177766142273692 la0=7.4043489218813e-06 wa0=9.64912404617634e-07 pa0=-7.53821991544092e-12
+  keta=-0.0171781577962286 lketa=-3.64042530028426e-08 wketa=-4.76076506622066e-09 pketa=3.7192696314378e-14
+  a1=0.0
+  a2=0.65972622
+  ags=0.318375533020026 lags=-1.39707639867554e-06 wags=-1.53222097901471e-07 pags=1.19702251143118e-12
+  b0=5.02741585822153e-07 lb0=-3.6703025281275e-12 wb0=-4.79983700173889e-13 pb0=3.74979394028168e-18
+  b1=-4.72456223437932e-10 lb1=3.6909867627882e-15 wb1=4.82688680325151e-16 pb1=-3.77092615409667e-21
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.5910241327219+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-3.32472811773205e-06 wnfactor=-3.16512733032638e-07 pnfactor=2.47270381872926e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-1.39105230758014 lpclm=1.88968869611914e-05 wpclm=2.47123981085771e-06 ppclm=-1.93061557389969e-11
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=5.82260891587051e-05 lalpha0=-2.14144638633761e-10 walpha0=-1.91302207364233e-11 palpha0=1.49451712147107e-16
+  alpha1=0.0
+  beta0=27.765730832484 lbeta0=-6.24776597292433e-06 wbeta0=-1.91151930689163e-06 pbeta0=1.49334310959245e-11
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.394636168 lkt1=1.48916248884492e-8
+  kt2=-0.019151
+  at=313675.63146176 lat=-1.27868902799144 wat=-0.0601106700280387 pat=4.69604751444168e-7
+  ute=-1.06279449536883 lute=-8.27369386428235e-07 wute=-1.0819920605047e-07 pute=8.45288552599504e-13
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.67 nmos
* DC IV MOS Parameters
+  lmin=2e-06 lmax=4e-06 wmin=7.5e-07 wmax=1.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.816591495340202+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-3.56340802804629e-08 wvth0=-1.23825517766513e-08 pvth0=2.03610226754717e-14
+  k1=0.88325
+  k2=-0.0205886927833808 lk2=-5.07998804519598e-09 wk2=-1.95681356497449e-08 pk2=1.70383303715562e-14
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=180550.393039494 lvsat=-0.133455031411977 wvsat=-0.0683782150575103 pvsat=1.29639470218364e-7
+  ua=-1.53929242046186e-10 lua=7.50290818019935e-18 wua=4.43713787799991e-18 pua=-2.86078360330635e-24
+  ub=1.26006832351362e-18 lub=4.35376281831252e-25 wub=5.07829472904586e-26 pub=1.39411453813813e-31
+  uc=-9.53685709082235e-12 luc=1.85803680428712e-16 wuc=5.13452413849898e-17 puc=-1.43376896432259e-22
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0367298568313111 lu0=9.60713099985856e-10 wu0=-1.0766190627986e-09 pu0=6.4138855538707e-15
+  a0=1.74418889139448 la0=1.43261908418917e-06 wa0=-6.28271835139666e-07 pa0=-1.46446628358153e-12
+  keta=-0.026727225088 wketa=4.9951159249559e-9
+  a1=0.0
+  a2=0.65972622
+  ags=-0.0699130136715613 lags=8.32100062644805e-08 wags=1.7760713080377e-07 pags=-6.42096670140367e-14
+  b0=-5.69952481316178e-07 lb0=4.19167681010381e-13 wb0=6.15942775070524e-13 pb0=-4.28246014645704e-19
+  b1=3.66966860261518e-10 lb1=4.90823921569774e-16 wb1=-3.74914628521062e-16 pb1=-5.01454186063132e-22
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.417667824345905+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.14850037751684e-06 wnfactor=6.32053887258115e-07 pnfactor=-1.1435508562035e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=3.56572142936 wpclm=-2.59288773167708e-6
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=2.66992179178013e-05 lalpha0=-9.39536124346994e-11 walpha0=1.05468832798526e-12 palpha0=7.25000566641353e-17
+  alpha1=0.0
+  beta0=27.6405330330995 lbeta0=-5.77046989521036e-06 wbeta0=-9.09121694042404e-07 pbeta0=1.11119545901454e-11
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.407041024 lkt1=6.21831039920647e-8
+  kt2=-0.019151
+  at=-59549.42292352 lat=0.144170282943521 wat=0.120221340056078 pat=-2.17881462551872e-7
+  ute=-1.38051100926234 lute=3.83872717282467e-07 wute=2.1639841210094e-07 pute=-3.92186632593369e-13
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.68 nmos
* DC IV MOS Parameters
+  lmin=1e-06 lmax=2e-06 wmin=7.5e-07 wmax=1.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.745009951687237+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=9.4095728217376e-08 wvth0=4.92072173103161e-08 pvth0=-9.1260333072527e-14
+  k1=0.88325
+  k2=-0.0233759104803806 lk2=-2.86130730860051e-11 wk2=-1.84000894475796e-08 pk2=1.49214381897086e-14
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=103597.471586061 lvsat=0.00600951844325293 wvsat=0.00853302534973943 pvsat=-9.74953957634982e-9
+  ua=-4.36389729591993e-10 lua=5.19416218337017e-16 wua=2.22791515847513e-16 pua=-3.98592283555063e-22
+  ub=2.04685732074306e-18 lub=-9.90549742251571e-25 wub=-2.66239929262326e-25 pub=7.13963425813982e-31
+  uc=1.57599791602339e-10 luc=-1.17104084917258e-16 wuc=-7.76270906722779e-17 puc=9.03643039590813e-23
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0366910183807602 lu0=1.0311014221036e-09 wu0=2.11610776237477e-09 pu0=6.27591790443301e-16
+  a0=5.67363734161128 la0=-5.68886180228295e-06 wa0=-4.13991332004082e-06 pa0=4.89980799859829e-12
+  keta=-0.0397792104470855 lketa=2.36545829377437e-08 wketa=9.05282841497086e-09 pketa=-7.35393842330377e-15
+  a1=0.0
+  a2=0.65972622
+  ags=1.61313246439456 lags=-2.96703390327196e-06 wags=-1.12112837670977e-06 pags=2.28953544773103e-12
+  b0=-1.16036802656051e-08 lb0=-5.92747951690411e-13 wb0=4.55012556867978e-14 pb0=6.05585686828122e-19
+  b1=5.81836854585723e-09 lb1=-9.38894760369602e-15 wb1=-5.94438277182341e-15 pb1=9.59229343089687e-21
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.0250884791188+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=4.7650057728345e-08 wnfactor=2.57924652418744e-08 pnfactor=-4.48014556722731e-14
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=6.27176362073505 lpclm=-4.90425768094789e-06 wpclm=-5.35753738483293e-06 ppclm=5.01047409380186e-12
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=-7.12461962841845e-05 lalpha0=8.35563877584709e-11 walpha0=7.66350507602612e-11 palpha0=-6.44769550649261e-17
+  alpha1=0.0
+  beta0=15.5001572278651 lbeta0=1.6231970230145e-05 wbeta0=9.46432061565137e-06 pbeta0=-7.68820835163577e-12
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.37273
+  kt2=-0.019151
+  at=16750.656 lat=0.005888903107584
+  ute=-1.75301501475075 lute=1.05897513657331e-06 wute=5.32318595596662e-07 pute=-9.64740154269272e-13
+  ua1=3.0044e-9
+  ub1=-4.4951544593405e-18 lub1=1.34593941222333e-24 wub1=3.85021582859374e-25 pub1=-6.97788475393028e-31
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.81e-6
+  sbref=2.81e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.69 nmos
* DC IV MOS Parameters
+  lmin=8.0e-07 lmax=1e-06 wmin=7.5e-07 wmax=1.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.960726842238767+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-8.11388677856887e-08 wvth0=-1.2328622966227e-07 pvth0=4.88623036673949e-14
+  k1=0.88325
+  k2=-0.0555437668748299 lk2=2.61024947189553e-08 wk2=1.82646988259573e-08 pk2=-1.48626892572632e-14
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=176898.485082619 lvsat=-0.0535355336564873 wvsat=-0.0371453087102691 pvsat=2.73566156006216e-8
+  ua=1.26170089005449e-09 lua=-8.60003923264129e-16 wua=-1.08312761635375e-15 pua=6.62252840620782e-22
+  ub=-1.12853893740362e-18 lub=1.58893895250627e-24 wub=1.99080976894687e-24 pub=-1.11951929783048e-30
+  uc=-2.01361339887947e-10 luc=1.74492964793035e-16 wuc=1.92185925740316e-16 puc=-1.28814522541459e-22
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0379236983943896 lu0=2.9751070551946e-11 wu0=2.10209529819184e-09 pu0=6.38974619547758e-16
+  a0=-8.83562698973907 la0=6.09753594758886e-06 wa0=7.68403685924808e-06 pa0=-4.70521239424453e-12
+  keta=0.0477691878561698 lketa=-4.74641327463296e-08 wketa=-5.96946472067588e-08 pketa=4.84921109333496e-14
+  a1=0.0
+  a2=0.65972622
+  ags=-8.77377586837771 lags=5.47062566413893e-06 wags=6.89401253354061e-06 pags=-4.22145205873813e-12
+  b0=-3.11170050195326e-06 lb0=1.92557230005205e-12 wb0=3.21273997433857e-12 pb0=-1.96727634492658e-18
+  b1=-2.33123868631427e-08 lb1=1.42750137222294e-14 wb1=2.38172865378247e-14 pb1=-1.45841819694254e-20
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.93918332703677+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-6.94902094649943e-07 wnfactor=-9.27752353802816e-07 pnfactor=7.29797328451216e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-1.46556969917063 lpclm=1.38105671881101e-06 wpclm=2.54737110011526e-06 ppclm=-1.41096764522702e-12
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=2.804625977232e-05 lalpha0=2.89755117535417e-12 walpha0=-9.97843782620009e-12 palpha0=5.88229979944561e-18
+  alpha1=0.0
+  beta0=30.9568369599999 lbeta0=3.6759528432614e-6
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.378853360000001 lkt1=4.97422576896017e-9
+  kt2=-0.019151
+  at=8691.59999999998 lat=0.0124355644224
+  ute=1.99291078575373 lute=-1.9839752445053e-06 wute=-2.66159297798332e-06 pute=1.62978919776639e-12
+  ua1=6.043729736e-09 lua1=-2.4689569604233e-15
+  ub1=-6.01348388729746e-18 lub1=2.57933306641218e-24 wub1=-1.92510791429688e-24 pub1=1.17881287980889e-30
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.41e-6
+  sbref=2.41e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.70 nmos
* DC IV MOS Parameters
+  lmin=6e-07 lmax=8.0e-07 wmin=7.5e-07 wmax=1.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.861219937758836+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-2.02072079240679e-08 wvth0=-4.99781424621387e-08 pvth0=3.97312278361622e-15
+  k1=0.88325
+  k2=-0.00564469523729805 lk2=-4.45250321128438e-09 wk2=-1.30713158913651e-08 pk2=4.32548065068307e-15
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=152849.321047124 lvsat=-0.0388093647476486 wvsat=-0.0480440613266411 pvsat=3.40303141827202e-8
+  ua=-1.20069947997467e-10 lua=-1.38958953747454e-17 wua=-2.5388688224791e-17 pua=1.45612163260081e-23
+  ub=2.19014049343661e-18 lub=-4.43207935456718e-25 wub=-8.28479144674308e-25 pub=6.06832798380657e-31
+  uc=1.68829556810732e-10 luc=-5.21882481278472e-17 wuc=-9.15879382031643e-17 puc=4.49504302102356e-23
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0334461506063181 lu0=2.77151477290846e-09 wu0=4.91685942162368e-09 pu0=-1.08460678473797e-15
+  a0=1.1222
+  keta=-0.0297440283296 wketa=1.94973502151625e-8
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.466116679618073+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=2.07109643963832e-07 wnfactor=3.65755617514116e-07 pnfactor=-6.22641686731105e-14
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-5.27220243593632 lpclm=3.71199498231117e-06 wpclm=4.92094211150975e-06 ppclm=-2.86439062406027e-12
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=5.79028712003449e-05 lalpha0=-1.53847268400369e-11 walpha0=7.91652461038112e-13 palpha0=-7.12614206680737e-19
+  alpha1=0.0
+  beta0=34.6690869137664 lbeta0=1.40280855557193e-06 wbeta0=2.34052968185527e-06 pbeta0=-1.4331905832685e-12
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.37073
+  kt2=-0.019151
+  at=9620.20799999993 lat=0.011866944314112
+  ute=-1.13989264 lute=-6.56469259929603e-8
+  ua1=2.0117e-9
+  ub1=-1.8012e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.02e-6
+  sbref=2.01e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.71 nmos
* DC IV MOS Parameters
+  lmin=5e-07 lmax=6e-07 wmin=7.5e-07 wmax=1.0e-6
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={1.05889416799735+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-1.01715409323695e-07 wvth0=-1.14735473164668e-07 pvth0=3.06749014961742e-14
+  k1=0.88325
+  k2=-0.00577842263336609 lk2=-4.39736259169926e-09 wk2=-1.92917457652097e-08 pk2=6.89038782314464e-15
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=-61867.4892469116 lvsat=0.0497261059417532 wvsat=0.126578936919211 pvsat=-3.79730344219814e-8
+  ua=-2.50132665583184e-10 lua=3.97336453436791e-17 wua=7.45515195909221e-17 pua=-2.66477292038918e-23
+  ub=-1.86313811840312e-18 lub=1.22810475423483e-24 wub=2.42261929587225e-24 pub=-7.3371212820055e-31
+  uc=-5.09057224953751e-11 luc=3.84165180001159e-17 wuc=1.54018459899079e-16 puc=-5.6321929557651e-23
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0334483048357185 lu0=2.77062650657445e-09 wu0=5.740275643188e-09 pu0=-1.42413093587296e-15
+  a0=1.1222
+  keta=-0.0893503190531394 lketa=2.45778194917813e-08 wketa=8.03945939831923e-08 pketa=-2.51101259063344e-14
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={-0.39921016233917+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=5.63915052669114e-07 wnfactor=1.32498331939977e-06 pnfactor=-4.57788282357833e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=11.3678682588692 lpclm=-3.14930520770219e-06 wpclm=-8.35309037568783e-06 ppclm=2.60897083558084e-12
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=3.97214654722855e-05 lalpha0=-7.88787872775175e-12 walpha0=-3.86187397506119e-12 palpha0=1.20620226987471e-18
+  alpha1=0.0
+  beta0=41.5418261724672 lbeta0=-1.43106925940372e-06 wbeta0=-4.68105936371049e-06 pbeta0=1.46206335742389e-12
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.4331972 lkt1=2.57574753792e-8
+  kt2=-0.019151
+  at=30604.09344 lat=0.00321453292732415
+  ute=-1.787281168 lute=2.01294670088448e-7
+  ua1=-1.088859472e-09 lua1=1.27847229044659e-15
+  ub1=-4.24455148335244e-18 lub1=1.00748177723961e-24 wub1=2.36288555022811e-24 pub1=-9.74302776238857e-31
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=1.81e-6
+  sbref=1.81e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.72 nmos
* DC IV MOS Parameters
+  lmin=2.0e-05 lmax=1.0e-04 wmin=7e-07 wmax=7.5e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.798119+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+  k1=0.88325
+  k2=-0.041488
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=101000.0
+  ua=-1.471835e-10
+  ub=1.48747e-18
+  uc=5.7002e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0377669
+  a0=0.80798
+  keta=-0.020254
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=1.92633e-7
+  b1=-1.606e-10
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.14929+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.20557
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=2.8066e-5
+  alpha1=0.0
+  beta0=28.726
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.39073
+  kt2=-0.019151
+  at=60000.0
+  ute=-1.1327
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.73 nmos
* DC IV MOS Parameters
+  lmin=8e-06 lmax=2.0e-05 wmin=7e-07 wmax=7.5e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.794615818332005+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=6.94062122754346e-08 wvth0=-1.6940658945086e-21
+  k1=0.88325
+  k2=-0.0434202511039998 lk2=3.8282408108819e-08 wk2=-1.05879118406788e-22
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=93903.7948000003 lvsat=0.140592401747352
+  ua=-1.46175057628e-10 lua=-1.99795991107014e-17
+  ub=1.34048089816001e-18 lub=2.91219747399231e-24
+  uc=5.98378779679999e-11 luc=-5.61853671570138e-17
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.03746956249184 lu0=5.89095061706839e-9
+  a0=0.601237790544403 la0=4.09604611911673e-6
+  keta=-0.019222771648 lketa=-2.04310426025509e-8
+  a1=0.0
+  a2=0.65972622
+  ags=0.173728883712001 lags=-2.6704817300707e-7
+  b0=2.966021716e-07 lb0=-2.05987216138086e-12 pb0=-3.08148791101958e-33
+  b1=-2.651550968e-10 lb1=2.07148070831413e-15
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.13876938752+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=2.0843790937957e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-0.329724752439998 lpclm=1.06054394943781e-05 ppclm=6.46234853557053e-27
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=2.62763240280001e-05 lalpha0=3.54576616883907e-11
+  alpha1=0.0
+  beta0=29.87180928 lbeta0=-2.27011584472778e-5
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.389427944000001 lkt1=-2.57967709628204e-8
+  kt2=-0.019151
+  at=1407.48000000021 lat=1.16085469332672
+  ute=-1.109262992 lute=-4.64341877330686e-7
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.74 nmos
* DC IV MOS Parameters
+  lmin=4e-06 lmax=8e-06 wmin=7e-07 wmax=7.5e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.808628545004005+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-4.00659167623841e-8
+  k1=0.88325
+  k2=-0.0356912466880002 lk2=-2.20991713344567e-8
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=122288.615600001 lvsat=-0.0811593556420398
+  ua=-1.50208827116e-10 lua=1.15335634761027e-17
+  ub=1.92843730552001e-18 lub=-1.6811155336569e-24
+  uc=4.84943660960001e-11 luc=3.243395900704e-17
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0386589125244801 lu0=-3.40065145952614e-9
+  a0=1.4282066283668 la0=-2.36451230348138e-6
+  keta=-0.023347685056 lketa=1.17941669116508e-8
+  a1=0.0
+  a2=0.65972622
+  ags=0.119813348864001 lags=1.54158100845209e-7
+  b0=-1.192745148e-07 lb0=1.18909624734257e-12 wb0=-1.0097419586829e-28 pb0=3.85185988877447e-34
+  b1=1.530652904e-10 lb1=-1.19579747854238e-15
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.18085183744+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.20324329098672e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=1.81145425732 lpclm=-6.12217036601431e-6
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=3.3435027916e-05 lalpha0=-2.04685384091718e-11
+  alpha1=0.0
+  beta0=25.2885721600001 lbeta0=1.31046299018346e-5
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.394636168000002 lkt1=1.48916248884475e-8
+  kt2=-0.019151
+  at=235777.560000001 lat=-0.670123119980158
+  ute=-1.203011024 lute=2.68049247992069e-7
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.75 nmos
* DC IV MOS Parameters
+  lmin=2e-06 lmax=4e-06 wmin=7e-07 wmax=7.5e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.800544811736003+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-9.24800941037119e-9
+  k1=0.88325
+  k2=-0.045947252728 lk2=1.70001697080527e-08 wk2=-1.05879118406788e-22
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=91938.3200000003 lvsat=0.0345461688844795
+  ua=-1.481791067816e-10 lua=3.7955875753364e-18
+  ub=1.325878497568e-18 lub=6.16041102015601e-25
+  uc=5.7002e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0353346544711999 lu0=9.27253719028327e-9
+  a0=0.930004582880002 la0=-4.65198710198412e-7
+  keta=-0.020254
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=2.2825446408e-07 lb0=-1.35800989884891e-13
+  b1=-1.18889086960001e-10 lb1=-1.59016015375262e-16
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.23675333536+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-3.3343962207301e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.20557
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=2.8066e-5
+  alpha1=0.0
+  beta0=26.4623923360001 lbeta0=8.62963298734311e-6
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.407041024 lkt1=6.21831039920622e-8
+  kt2=-0.019151
+  at=96246.7200000002 lat=-0.13818467553792
+  ute=-1.100077952 lute=-1.24366207984124e-7
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.76 nmos
* DC IV MOS Parameters
+  lmin=1e-06 lmax=2e-06 wmin=7e-07 wmax=7.5e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.808778120111999+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-2.41695305792976e-8
+  k1=0.88325
+  k2=-0.0472207866399998 lk2=1.9308241063991e-8
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=114655.512 lvsat=-0.00662501599603216
+  ua=-1.476717796096e-10 lua=2.87614027774418e-18
+  ub=1.701834098976e-18 lub=-6.53167688177685e-26
+  uc=5.7002e-11
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0394333054592 lu0=1.84440445329525e-9
+  a0=0.308678616320002 la0=6.60852706733074e-7
+  keta=-0.028047551584 lketa=1.41245341035403e-8
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=4.73618921599994e-08 lb0=1.92037130338314e-13
+  b1=-1.88502177968e-09 lb1=3.04180984441814e-15 wb1=1.57772181044202e-30 pb1=2.63310734584192e-36
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.05851321552+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-1.04086362426566e-8
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-0.671127381280001 lpclm=1.58887022519947e-06 ppclm=1.21169035041947e-27
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=2.8066e-5
+  alpha1=0.0
+  beta0=27.7650733119999 lbeta0=6.26873735802319e-6
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.37273
+  kt2=-0.019151
+  at=16750.6560000001 lat=0.00588890310758405
+  ute=-1.0631775536 lute=-1.91242128418788e-7
+  ua1=3.0044e-9
+  ub1=-3.9962008e-18 lub1=4.4166773306881e-25
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.81e-6
+  sbref=2.81e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.77 nmos
* DC IV MOS Parameters
+  lmin=8.0e-07 lmax=1e-06 wmin=7e-07 wmax=7.5e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.800958875520003+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-1.78176767044149e-8
+  k1=0.88325
+  k2=-0.0318743448952004 lk2=6.8417739627872e-9
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=128761.475280001 lvsat=-0.0180837977830546
+  ua=-1.41935975440002e-10 lua=-1.78325993817145e-18
+  ub=1.45137310776002e-18 lub=1.38141710942682e-25
+  uc=4.76944928000004e-11 luc=7.56082316881947e-18
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0406478265680001 lu0=8.57805233857115e-10
+  a0=1.1222
+  keta=-0.0295897551040001 lketa=1.5377321542163e-8
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=1.0517241944e-06 lb0=-6.23842524814118e-13
+  b1=7.55269396e-09 lb1=-4.62478640869056e-15
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.736898955200019+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=2.50850205528653e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=1.83559623200001 lpclm=-4.47431607917948e-7
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.51150936000002e-05 lalpha0=1.05204875013504e-11
+  alpha1=0.0
+  beta0=30.9568369600001 lbeta0=3.6759528432614e-6
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.378853360000001 lkt1=4.97422576895763e-9
+  kt2=-0.019151
+  at=8691.60000000033 lat=0.0124355644223999
+  ute=-1.45627652 lute=1.28086313550724e-7
+  ua1=6.043729736e-09 lua1=-2.46895696042331e-15
+  ub1=-8.50825218400005e-18 lub1=4.10696950614182e-24
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.41e-6
+  sbref=2.41e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.78 nmos
* DC IV MOS Parameters
+  lmin=6e-07 lmax=8.0e-07 wmin=7e-07 wmax=7.5e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.796452719039998+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-1.50583948700779e-8
+  k1=0.88325
+  k2=-0.0225839557534401 lk2=1.15293423727837e-9
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=90588.4991200007 lvsat=0.00529088974685599
+  ua=-1.52971425368e-10 lua=4.97414332893958e-18
+  ub=1.11650535368001e-18 lub=3.43193292005005e-25
+  uc=5.01397509600001e-11 luc=6.06350356815741e-18
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0398179622400001 lu0=1.36596103700738e-9
+  a0=1.1222
+  keta=-0.0044772
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.940103364800002+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.26420830171825e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=1.1049
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=5.892878224e-05 lalpha0=-1.63082113457126e-11
+  alpha1=0.0
+  beta0=37.7022047999999 lbeta0=-4.54478718412885e-7
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.37073
+  kt2=-0.019151
+  at=9620.20799999987 lat=0.0118669443141121
+  ute=-1.13989264000001 lute=-6.56469259929595e-8
+  ua1=2.0117e-9
+  ub1=-1.8012e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.02e-6
+  sbref=2.01e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.79 nmos
* DC IV MOS Parameters
+  lmin=5e-07 lmax=6e-07 wmin=7e-07 wmax=7.5e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.910207219680011+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-6.19634706459721e-8
+  k1=0.88325
+  k2=-0.0307788059187202 lk2=4.53196597502935e-9
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=102167.532640001 lvsat=0.000516437381353096
+  ua=-1.53520540016001e-10 lua=5.20056306643769e-18
+  ub=1.27636059200001e-18 lub=2.77279222457084e-25
+  uc=1.4868847584e-10 luc=-3.45716834539624e-17
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0408871905120005 lu0=9.25079728243973e-10
+  a0=1.1222
+  keta=0.0148339102079999 lketa=-7.96266593872588e-9
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.3178501408+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-2.93377644569125e-8
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=0.543007536000005 lpclm=2.31688491035903e-7
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=3.471682096e-05 lalpha0=-6.32474807936256e-12
+  alpha1=0.0
+  beta0=35.4755904000003 lbeta0=4.63634556825622e-7
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.433197200000006 lkt1=2.57574753792004e-8
+  kt2=-0.019151
+  at=30604.0934400004 lat=0.00321453292732421
+  ute=-1.78728116800001 lute=2.0129467008845e-7
+  ua1=-1.08885947199999e-09 lua1=1.27847229044659e-15
+  ub1=-1.18246238400003e-18 lub1=-2.55127793630978e-25
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=1.81e-6
+  sbref=1.81e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.80 nmos
* DC IV MOS Parameters
+  lmin=2.0e-05 lmax=1.0e-04 wmin=4.2e-07 wmax=7.0e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.83241216635+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} wvth0=-2.47479378418083e-8
+  k1=0.88325
+  k2=-0.02922094905 wk2=-8.85261545447511e-9
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=57307.405 wvsat=0.03153111072251
+  ua=-3.8958307672e-10 wua=1.74929593736602e-16
+  ub=1.0350702465e-18 wub=3.26477901311303e-25
+  uc=2.369310005e-11 wuc=2.40376341201171e-17
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.032634045365 wu0=3.70416561018483e-9
+  a0=0.341052853 wa0=3.36961711049726e-7
+  keta=-0.0287149054 wketa=6.1058800691532e-9
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=3.505194256e-07 wb0=-1.13940002125645e-13
+  b1=-1.0851006085e-09 wb1=6.67173260128893e-16
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.604489083500001+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} wnfactor=3.93159939799557e-7
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-0.25880184 wpclm=3.3511765331072e-7
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=1.33083134e-05 walpha0=1.06500025963828e-11
+  alpha1=0.0
+  beta0=35.7578263 wbeta0=-5.0745737040054e-6
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.39546205 wkt1=3.41492173889994e-9
+  kt2=-0.019151
+  at=-255470 wat=0.22766144926
+  ute=-1.28065543 wute=1.0677321970294e-7
+  ua1=3.0044e-9
+  ub1=-4.22602047e-18 wub1=3.4171983533926e-25
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.81 nmos
* DC IV MOS Parameters
+  lmin=8e-06 lmax=2.0e-05 wmin=4.2e-07 wmax=7.0e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.825888874676532+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=1.29241646460744e-07 wvth0=-2.25684512954826e-08 pvth0=-4.31807197632866e-14
+  k1=0.88325
+  k2=-0.0365731731593924 lk2=1.45664734402583e-07 wk2=-4.94124857534963e-09 pk2=-7.74933148285051e-14
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=39018.00052778 lvsat=0.362355826643525 wvsat=0.0396087725229018 pvsat=-1.60037349683726e-7
+  ua=-3.85299750696712e-10 lua=-8.4862694370922e-17 wua=1.72566247750581e-16 pua=4.68234047592998e-23
+  ub=4.69660871682132e-19 lub=1.12020805114415e-23 wub=6.28434238667965e-25 pub=-5.98246041303954e-30
+  uc=3.10021501308248e-11 luc=-1.44809356042128e-16 wuc=2.08095336795202e-17 puc=6.39562105708542e-23
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0314506788480275 lu0=2.34452550454101e-08 wu0=4.34357553262649e-09 pu0=-1.26682042251481e-14
+  a0=-0.396208698625538 la0=1.46068735806865e-05 wa0=7.19815238481399e-07 pa0=-7.58522272426153e-12
+  keta=-0.0260570690069728 lketa=-5.2657947651683e-08 wketa=4.93202536348159e-09 pketa=2.32568038439469e-14
+  a1=0.0
+  a2=0.65972622
+  ags=0.194989800935123 lags=-6.88276608699775e-07 wags=-1.53431110014046e-08 pags=3.03982870445125e-13
+  b0=6.16224165289484e-07 lb0=-5.2642315795206e-12 wb0=-2.30657768721966e-13 pb0=2.31245160897589e-18
+  b1=3.28344764263096e-08 lb1=-6.72026057191533e-13 wb1=-2.38866138857043e-14 pb1=4.86467881005728e-19
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.34720463752326+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=5.09740589126502e-06 wnfactor=5.71239034353148e-07 pnfactor=-3.5281628558715e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-1.63844377020123 lpclm=2.73339294808354e-05 wpclm=9.44447548919536e-07 ppclm=-1.20722486266468e-11
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=-8.38369239721979e-06 lalpha0=4.29769307368467e-10 walpha0=2.50126781333913e-11 palpha0=-2.84558153598192e-16
+  alpha1=0.0
+  beta0=39.7491727527818 lbeta0=-7.9077897014921e-05 wbeta0=-7.12807836904077e-06 pbeta0=4.06847244012481e-11
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.4075096812054 lkt1=2.3869171744547e-07 wkt1=1.30488303081745e-08 pkt1=-1.90870233567746e-13
+  kt2=-0.019151
+  at=-476312.5644964 lat=4.37540709090435 wat=0.344750491871183 pat=-2.31980745413108e-6
+  ute=-1.30024549076202 lute=3.88124866077558e-07 wute=1.37824048091602e-07 pute=-6.15189445114507e-13
+  ua1=3.0044e-9
+  ub1=-4.53429555454316e-18 lub1=6.1076495553975e-24 wub1=5.64189016300507e-25 pub1=-4.40763416284904e-30
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.82 nmos
* DC IV MOS Parameters
+  lmin=4e-06 lmax=8e-06 wmin=4.2e-07 wmax=7.0e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.841860005700259+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=4.46980460336768e-09 wvth0=-2.39817494631408e-08 pvth0=-3.2139559609356e-14
+  k1=0.88325
+  k2=-0.00460257335305317 lk2=-1.04100333406074e-07 wk2=-2.2435389821551e-08 pk2=5.91767946182789e-14
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=103155.53613226 lvsat=-0.138708151710635 wvsat=0.0138075398625303 pvsat=4.15305490732694e-8
+  ua=-3.96058412304773e-10 lua=-8.12414978449174e-19 wua=1.7741931994816e-16 pua=8.90957411955519e-24
+  ub=2.54264334997538e-18 lub=-4.992755131098e-24 wub=-4.43246705629579e-25 pub=2.38987120861015e-30
+  uc=-3.52359310701306e-11 luc=3.72664790295019e-16 wuc=6.04246387923154e-17 puc=-2.4553030124562e-22
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0355401110408115 lu0=-8.50276329383591e-09 wu0=2.25070804110125e-09 pu0=3.68197982212442e-15
+  a0=2.25358124462117 la0=-6.09417578537771e-06 wa0=-5.95638194816897e-07 pa0=2.69154148901835e-12
+  keta=-0.0453927939835276 lketa=9.83992326687552e-08 wketa=1.59090292184217e-08 pketa=-6.24992385441404e-14
+  a1=0.0
+  a2=0.65972622
+  ags=0.0560305971946303 lags=3.97319381213411e-07 wags=4.60293330042139e-08 pags=-1.75479283267953e-13
+  b0=-4.62761787616192e-07 lb0=3.16516922385872e-12 wb0=2.47880338325987e-13 pb0=-1.42604887208669e-18
+  b1=-1.08591894182133e-07 lb1=4.32844269262148e-13 wb1=7.84766699630294e-14 pb1=-3.13228486483953e-19
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.755820894145397+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=1.90515839947067e-06 wnfactor=3.06726980476097e-07 pnfactor=-1.46170581493388e-12
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=3.8801239506037 lpclm=-1.57789757928469e-05 wpclm=-1.49287203351573e-06 ppclm=6.96891089071719e-12
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=4.413658170484e-05 lalpha0=1.9463279271077e-11 walpha0=-7.72286190414671e-12 palpha0=-2.8817115683493e-17
+  alpha1=0.0
+  beta0=26.8866952474882 lbeta0=2.14080990488741e-05 wbeta0=-1.15329831107056e-06 pbeta0=-5.99226493771452e-12
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.363829197526 lkt1=-1.02554897700519e-07 wkt1=-2.22320966983258e-08 pkt1=8.47562225985085e-14
+  kt2=-0.019151
+  at=136455.2249572 lat=-0.411740770284432 wat=0.0716767576623169 pat=-1.86463689716719e-7
+  ute=-1.36289920076006 lute=8.77596700228801e-07 wute=1.15384581864311e-07 pute=-4.39884795286261e-13
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.83 nmos
* DC IV MOS Parameters
+  lmin=2e-06 lmax=4e-06 wmin=4.2e-07 wmax=7.0e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.841256003997288+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=6.77246203966564e-09 wvth0=-2.93795575848967e-08 pvth0=-1.15613013856931e-14
+  k1=0.88325
+  k2=-0.0402958437505104 lk2=3.19744062878866e-08 wk2=-4.0783844998772e-09 pk2=-1.08062776217298e-14
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=40557.6958624 lvsat=0.0999358482724015 wvsat=0.0370792384538921 pvsat=-4.71889852477287e-8
+  ua=-5.10985593954478e-10 lua=4.37328617003262e-16 wua=2.61822203920205e-16 pua=-3.12862578950897e-22
+  ub=8.8810129803352e-19 lub=1.31491509703381e-24 wub=3.15925418261654e-25 pub=-5.04348009496849e-31
+  uc=7.29449101156608e-11 luc=-3.97569250678563e-17 wuc=-1.15053286282475e-17 puc=2.8690903030619e-23
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0318976594566588 lu0=5.38348600868665e-09 wu0=2.48033494820381e-09 pu0=2.80656489760863e-15
+  a0=0.83095099925396 la0=-6.70631286275461e-07 wa0=7.14828110524003e-08 pa0=1.48252061986615e-13
+  keta=-0.0195820489 wketa=-4.84918886923806e-10
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=5.25508451826388e-07 lb0=-6.02448987696843e-13 wb0=-2.14515718289083e-13 pb0=3.36760260804978e-19
+  b1=7.648676584652e-09 lb1=-1.03038433326148e-14 wb1=-5.60552590744418e-15 pb1=7.32109579210448e-21
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.39696285099775+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-5.39090163748014e-07 wnfactor=-1.15616478636109e-07 pnfactor=1.48409358604106e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-0.25880184 wpclm=3.3511765331072e-7
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=5.10614787826804e-05 lalpha0=-6.93675515506865e-12 walpha0=-1.65948712273516e-11 palpha0=5.00596485169655e-18
+  alpha1=0.0
+  beta0=31.8008413316164 lbeta0=2.67372302309329e-06 wbeta0=-3.85253442527854e-06 pbeta0=4.2981300729806e-12
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.407041024 lkt1=6.21831039920643e-8
+  kt2=-0.019151
+  at=36112.8381040001 lat=-0.029201876558051 wat=0.0433960969413036 pat=-7.86483087462144e-8
+  ute=-1.100077952 lute=-1.24366207984129e-7
+  ua1=3.0044e-9
+  ub1=-3.7525e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=3.0e-6
+  sbref=3.0e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.84 nmos
* DC IV MOS Parameters
+  lmin=1e-06 lmax=2e-06 wmin=4.2e-07 wmax=7.0e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.82578172165797+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=3.48170609973746e-08 wvth0=-1.2270785084462e-08 pvth0=-4.25681457040414e-14
+  k1=0.88325
+  k2=-0.0299447508804896 lk2=1.32147480402046e-08 wk2=-1.24673894141367e-08 pk2=4.39741798855967e-15
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=109029.32033148 lvsat=-0.0241577417313932 wvsat=0.00406018622712084 pvsat=1.26526317887293e-8
+  ua=-2.67421201897886e-10 lua=-4.09189903901417e-18 wua=8.64181285897201e-17 pua=5.02854131725312e-24
+  ub=1.62833675632821e-18 lub=-2.66402725101606e-26 wub=5.30399453005169e-26 pub=-2.79112029723554e-32
+  uc=5.100807e-11 wuc=4.32556753594001e-18
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0337297308117397 lu0=2.0631571373047e-09 wu0=4.11603027293691e-09 pu0=-1.57864624436862e-16
+  a0=-0.0762723352915353 la0=9.73562222961385e-07 wa0=2.77802933838078e-07 pa0=-2.25669324062289e-13
+  keta=-0.0268297504152304 lketa=1.31352703733066e-08 wketa=-8.78835955851926e-10 pketa=7.13910085032933e-16
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=1.43040246936817e-07 lb0=9.0711908879902e-14 wb0=-6.9047050151528e-14 pb0=7.31221566672348e-20
+  b1=-3.43781898757057e-09 lb1=9.78861170676472e-15 wb1=1.12058852745189e-15 pb1=-4.86888353837732e-21
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={0.912293378048136+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=3.39293770179602e-07 wnfactor=1.05520715470271e-07 pnfactor=-2.52365539213873e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-1.70300390545384 lpclm=2.61737939449635e-06 wpclm=7.44661948682245e-07 ppclm=-7.42231870096448e-13
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=4.53798608396488e-05 lalpha0=3.36024558133346e-12 walpha0=-1.24946861858193e-11 palpha0=-2.42494810573393e-18
+  alpha1=0.0
+  beta0=27.6953096200224 lbeta0=1.01143259431567e-05 wbeta0=5.03455264251677e-08 pbeta0=-2.77519976717028e-12
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.37273
+  kt2=-0.019151
+  at=16750.656 lat=0.005888903107584
+  ute=-1.0631775536 lute=-1.9124212841879e-7
+  ua1=3.0044e-9
+  ub1=-4.38060225688e-18 lub1=1.13833233182487e-24 wub1=2.77406386569107e-25 pub1=-5.02753581009109e-31
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.81e-6
+  sbref=2.81e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.85 nmos
* DC IV MOS Parameters
+  lmin=8.0e-07 lmax=1e-06 wmin=4.2e-07 wmax=7.0e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.995633498752792+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-1.03159652200724e-07 wvth0=-1.4048849925293e-07 pvth0=6.15877193527158e-14
+  k1=0.88325
+  k2=-0.0378831936721389 lk2=1.96634309038018e-08 wk2=4.33633379066816e-09 pk2=-9.25285130473873e-15
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=50631.6168242882 lvsat=0.0232808151448251 wvsat=0.0563830373934321 pvsat=-2.98511038363074e-8
+  ua=-4.34840355940512e-10 lua=1.31908706879357e-16 wua=2.11376789423239e-16 pua=-9.64798773896042e-23
+  ub=2.28090763580987e-19 lub=1.11082995625415e-24 wub=8.82791489935539e-25 pub=-7.01948253734991e-31
+  uc=-1.40879838312959e-11 luc=5.28798679850996e-17 wuc=4.45858185207878e-17 puc=-3.27048512440273e-23
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0398236292169608 lu0=-2.88713591759892e-09 wu0=5.94788611956302e-10 pu0=2.70256674147754e-15
+  a0=1.1222
+  keta=-0.0594486043172943 lketa=3.96327396766936e-08 wketa=2.15478774055676e-08 pketa=-1.75041165401291e-14
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=9.3371294713784e-07 lb0=-5.51579989710597e-13 wb0=8.51637606767158e-14 pb0=-5.21488365577374e-20
+  b1=3.49797379083879e-08 lb1=-2.14193527918706e-14 wb1=-1.97929456817058e-14 pb1=1.2119933186953e-20
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.06815845962404+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=2.12678953272557e-07 wnfactor=-2.39056071443644e-07 pnfactor=2.75465895606292e-14
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=2.9386311435452 lpclm=-1.15318785466733e-06 wpclm=-7.96013968195884e-07 ppclm=5.09314641516664e-13
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=-6.21958694471117e-06 lalpha0=4.52763345966892e-11 walpha0=1.53963428925352e-11 palpha0=-2.50818351031281e-17
+  alpha1=0.0
+  beta0=28.483294988856 lbeta0=9.47421706057986e-06 wbeta0=1.78505135181182e-06 pbeta0=-4.18436375854159e-12
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.37885336 lkt1=4.97422576896017e-9
+  kt2=-0.019151
+  at=8691.60000000001 lat=0.0124355644224
+  ute=-1.45627652 lute=1.28086313550717e-7
+  ua1=6.04372973599999e-09 lua1=-2.4689569604233e-15
+  ub1=-6.5862448996e-18 lub1=2.93005525364147e-24 wub1=-1.38703193284554e-24 pub1=8.49329585630902e-31
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.41e-6
+  sbref=2.41e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.86 nmos
* DC IV MOS Parameters
+  lmin=6e-07 lmax=8.0e-07 wmin=4.2e-07 wmax=7.0e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.820888289311585+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=3.84313036766718e-09 wvth0=-1.76341247710513e-08 pvth0=-1.36404369000206e-14
+  k1=0.88325
+  k2=0.0120230776407434 lk2=-1.08959756468433e-08 wk2=-2.49744425051796e-08 pk2=8.69519220915552e-15
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=59172.032025216 lvsat=0.0180512114623498 wvsat=0.0226719448106876 pvsat=-9.20858824856005e-9
+  ua=-2.31855261729574e-10 lua=7.61362623060751e-18 wua=5.69271515810207e-17 pua=-1.9048039518518e-24
+  ub=1.87214806173783e-18 lub=1.04114486529982e-25 wub=-5.45315605411597e-25 pub=1.72533132601493e-31
+  uc=4.67480556367561e-11 luc=1.56277709213906e-17 wuc=2.44764406358163e-18 puc=-6.90213004959953e-24
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0321985968009628 lu0=1.78194593188357e-09 wu0=5.49857602400466e-09 pu0=-3.00198827266553e-16
+  a0=1.1222
+  keta=0.00527523957999999 wketa=-7.03792604242364e-9
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={1.00623161078272+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=2.50598992184657e-07 wnfactor=-4.77219777393979e-08 pnfactor=-8.96141640418544e-14
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=2.4595809013464 lpclm=-8.5984814556029e-07 wpclm=-9.77616309903841e-07 ppclm=6.20516293028748e-13
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=0.000136362758546264 lalpha0=-4.20319685118725e-11 walpha0=-5.58808484732259e-11 palpha0=1.85637551490166e-17
+  alpha1=0.0
+  beta0=50.0993090146281 lbeta0=-3.76204650390524e-06 wbeta0=-8.94646943332003e-06 pbeta0=2.38693275294292e-12
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.37073
+  kt2=-0.019151
+  at=9620.20799999998 lat=0.011866944314112
+  ute=-1.13989264 lute=-6.56469259929603e-8
+  ua1=2.0117e-9
+  ub1=-1.8012e-18
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=2.02e-6
+  sbref=2.01e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.87 nmos
* DC IV MOS Parameters
+  lmin=5e-07 lmax=6e-07 wmin=4.2e-07 wmax=7.0e-7
+  level=54.0
+  tnom=30.0
+  version=4.5
+  toxm=1.16e-8
+  xj=1.5e-7
+  lln=1.0
+  lwn=1.0
+  wln=1.0
+  wwn=1.0
+  lint=9.3832e-8
+  ll=0.0
+  lw=0.0
+  lwl=0.0
+  wint=-1.0829e-8
+  wl=0.0
+  ww=0.0
+  wwl=0.0
+  xl=0.0
+  xw=0.0
+  mobmod=0.0
+  binunit=2.0
+  dwg=-4.1292e-9
+  dwb=-1.6944e-9
* BSIM4 - Model Selectors
+  igcmod=0.0
+  igbmod=0.0
+  rgatemod=0.0
+  rbodymod=1.0
+  trnqsmod=0.0
+  acnqsmod=0.0
+  fnoimod=1.0
+  tnoimod=1.0
+  permod=1.0
+  geomod=0.0
+  rdsmod=0.0
+  tempmod=0.0
+  lintnoi=0.0
+  vfbsdoff=0.0
+  lambda=0.0
+  vtl=0.0
+  lc=5.0e-9
+  xn=3.0
+  rnoia=0.794
+  rnoib=0.38
+  tnoia=7.50e+6
+  tnoib=7.2e+6
* BSIM4 - Process Parameters
+  epsrox=3.9
+  toxe={1.0904e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.0904e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}
+  dtox=0.0
+  ndep=1.7000000000000000e+17
+  nsd=1.0e+20
+  rshg=0.1
+  rsh=1.0
* Threshold Voltage Parameters
+  vth0={0.924284804192327+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))} lvth0=-3.87909749921988e-08 wvth0=-1.01592014839976e-08 pvth0=-1.67226168685111e-14
+  k1=0.88325
+  k2=0.0128316267389061 lk2=-1.12293695477833e-08 wk2=-3.14718176108372e-08 pk2=1.13742938707219e-14
+  k3=-0.884
+  dvt0=0.0
+  dvt1=0.53
+  dvt2=-0.19251
+  dvt0w=0.16
+  dvt1w=6909100.0
+  dvt2w=-0.036016
+  w0=0.0
+  k3b=0.43
* NEW BSIM4 Parameters for Level 54
+  phin=0.0
+  lpe0=2.5e-8
+  lpeb=-2.182e-7
+  vbm=-3.0
+  dvtp0=0.0
+  dvtp1=0.0
* Mobility Parameters
+  vsat=121177.384856784 lvsat=-0.00751582770280768 wvsat=-0.0137186119310599 pvsat=5.79654835610521e-9
+  ua=-4.97692054119712e-10 lua=1.17227705857587e-16 wua=2.48374126525056e-16 pua=-8.08452838123757e-23
+  ub=2.59647279754237e-19 lub=7.69006608969969e-25 wub=7.33719295488652e-25 pub=-3.54859002296113e-31
+  uc=2.3034596854428e-10 luc=-6.00762580952462e-17 wuc=-5.89287828699853e-17 puc=1.84055803264797e-23
+  rdsw=724.62
+  prwb=0.05626
+  prwg=0.048
+  wr=1.0
+  u0=0.0236484514077593 lu0=5.30747868273555e-09 wu0=1.24404739844882e-08 pu0=-3.1625932647005e-15
+  a0=1.1222
+  keta=0.0550467294745888 lketa=-2.05225770571752e-08 wketa=-2.90199027262879e-08 pketa=9.06396033791787e-15
+  a1=0.0
+  a2=0.65972622
+  ags=0.16025
+  b0=3.2933e-8
+  b1=0.0
* BSIM4 - Mobility Parameters
+  eu=1.67
+  rdswmin=0.0
+  rdw=0.0
+  rdwmin=0.0
+  rsw=0.0
+  rswmin=0.0
* Subthreshold Current Parameters
+  voff={-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+  nfactor={2.55769186340056+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))} lnfactor=-3.89123922538774e-07 wnfactor=-8.94741697848475e-07 pnfactor=2.59642559269042e-13
+  up=0.0
+  ud=0.0
+  lp=1.0
+  tvfbsdoff=0.0
+  tvoff=0.0
+  cit=-8.0e-4
+  cdsc=0.0
+  cdscb=0.0
+  cdscd=0.0
+  eta0=0.032
+  etab=-0.01932
+  dsub=0.504
* BSIM4 - Sub-threshold parameters
+  voffl=-4.2579486e-7
+  minv=0.0
* Rout Parameters
+  pclm=-0.317684066054399 lpclm=2.85318182037887e-07 wpclm=6.21124980155373e-07 ppclm=-3.87022955491089e-14
+  pdiblc1=0.21098
+  pdiblc2=2.0e-4
+  pdiblcb=-0.26831
+  drout=0.36075
+  pscbe1=937310000.0
+  pscbe2=1.68e-6
+  pvag=1.99
+  delta=0.0246
+  alpha0=9.67674098405984e-05 lalpha0=-2.57053808079731e-11 walpha0=-4.47793038703949e-11 palpha0=1.39861886536637e-17
+  alpha1=0.0
+  beta0=53.517636179504 lbeta0=-5.17154585376156e-06 wbeta0=-1.30201866731453e-05 pbeta0=4.06667302474351e-12
* BSIM4 - Rout Parameters
+  fprout=10.125
+  pdits=0.0
+  pditsl=0.0
+  pditsd=0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+  agidl=5.06e-11
+  bgidl=1058000000.0
+  cgidl=4000.0
+  egidl=0.8
* BSIM4 - Gate Leakage Current Parameters
+  aigbacc=1.0
+  bigbacc=0.0
+  cigbacc=0.0
+  nigbacc=1.0
+  aigbinv=0.35
+  bigbinv=0.03
+  cigbinv=0.006
+  eigbinv=1.1
+  nigbinv=3.0
+  aigc=0.43
+  bigc=0.054
+  cigc=0.075
+  nigc=1.0
+  aigsd=0.43
+  bigsd=0.054
+  cigsd=0.075
+  dlcig=0.0
+  poxedge=1.0
+  pigcd=1.0
+  ntox=1.0
+  toxref=1.16e-8
* Temperature Effects Parameters
+  kt1=-0.35929772156 lkt1=-4.71393996283589e-09 wkt1=-5.33301498120534e-08 pkt1=2.19899406529029e-14
+  kt2=-0.019151
+  at=73485.497462784 lat=-0.0144670136818145 wat=-0.0309457082642743 pat=1.27600295628578e-8
+  ute=-2.5548504173968 lute=5.17791104107726e-07 wute=5.53922489381196e-07 pute=-2.28402183581485e-13
+  ua1=-1.088859472e-09 lua1=1.27847229044659e-15
+  ub1=-9.81983342406719e-18 lub1=3.30637123154617e-24 wub1=6.23322791003282e-24 pub1=-2.57018426351129e-30
+  uc1=-5.9821e-11
+  kt1l=0.0
+  prt=0.0
* BSIM4 - High Speed RF Model Parameters
+  xrcrg1=12.0
+  xrcrg2=1.0
+  rbpb=50.0
+  rbpd=50.0
+  rbps=50.0
+  rbdb=50.0
+  rbsb=50.0
+  gbmin=1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+  noia=2.6e+41
+  noib=0.0
+  noic=0.0
+  em=4.1000000e+7
+  af=1.0
+  ef=0.89
+  kf=0.0
+  ntnoi=1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+  dmcg=0.0
+  dmcgt=0.0
+  dmdg=0.0
+  xgw=0.0
+  xgl=0.0
+  ngcon=1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+  diomod=1.0
+  njs=1.0773
+  jss=0.000375
+  jsws=5.84e-11
+  xtis=0.76
+  bvs=12.636
+  xjbvs=1.0
+  ijthsrev=0.1
+  ijthsfwd=0.1
* Diode and FET Capacitance Parameters
+  tpb=0.001344
+  tpbsw=0.00099005
+  tpbswg=0.0
+  tcj=0.00067434
+  tcjsw=0.0002493
+  tcjswg=0.0
+  cgdo=2.338769804e-10
+  cgso=2.338769804e-10
+  cgbo=0.0
+  capmod=2.0
+  xpart=0.0
+  cgsl=3.8123e-11
+  cgdl=3.8123e-11
+  cf=0.0
+  clc=1.0e-7
+  cle=0.6
+  dlc=8.332e-8
+  dwc=-3.2175e-8
+  vfbcv=-1.0
+  acde=0.4176
+  moin=15.0
+  noff=4.0
+  voffcv=-0.4104
+  ngate=1.0e+23
+  lwc=0.0
+  llc=0.0
+  lwlc=0.0
+  wlc=0.0
+  wwc=0.0
+  wwlc=0.0
* BSIM4 - FET and Diode capacitance parameters
+  ckappas=0.6
+  cjs=0.000695881536
+  mjs=0.295
+  pbs=0.72468
+  cjsws=6.627678344e-11
+  mjsws=0.037586
+  pbsws=0.29067
+  cjswgs=4.200444e-11
+  mjswgs=0.78692
+  pbswgs=0.54958
* Stress Parameters
+  saref=1.81e-6
+  sbref=1.81e-6
+  wlod={0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+  kvth0={0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+  lkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+  wkvth0={0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+  pkvth0=0.0
+  llodvth=0.0
+  wlodvth=1.0
+  stk2=0.0
+  lodk2=1.0
+  lodeta0=1.0
+  ku0={0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+  lku0={0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+  wku0={0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+  pku0=0.0
+  llodku0=0.0
+  wlodku0=1.0
+  kvsat={0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+  steta0=0.0
+  tku0=0.0
.ends sky130_fd_pr__nfet_g5v0d10v5
