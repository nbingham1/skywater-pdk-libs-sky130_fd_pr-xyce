* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.subckt sky130_fd_pr__ind_05_125 a b ct sub
R31 net27 b r='1e-2'
R26 a net23 r='1e-2'
C24 net35 net27 c='103.1e-15'
C25 net23 net37 c='357e-15'
C1 net27 net31 c='357e-15'
R3 sub net31 r='3.67e3'
R2 net41 net27 r='1.7645'
R13 net23 net35 r='9.312'
R10 sub net37 r='3.67e3'
R9 net23 net39 r='1.7645'
L1 net39 ct l=2.895e-9
L2 ct net41 l=2.895e-9
.ends sky130_fd_pr__ind_05_125
