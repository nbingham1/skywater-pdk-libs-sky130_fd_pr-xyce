* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.subckt sky130_fd_pr__model__parasitic__rf_diode_ps2nw c0 c1
.param area=-1 perim=-1.0
+  ra1=7.6e+5
+  ra2=2000.0
+  rp1_diode=3750.0
+  wl={sqrt(0.0625*perim*perim-area)}
+  wi={perim/4+wl}
+  le={perim/4-wl}
rnwdiode_rf c0 a1 r={(ra1/area+ra2/(le/wi+wi/le))*(9.8286e-01*2-sky130_fd_pr__model__parasitic__diode_ps2nw__ajunction_mult)}
rp c0 p1 r={(rp1_diode/perim)*(9.8954e-01*2-sky130_fd_pr__model__parasitic__diode_ps2nw__pjunction_mult)}
da a1 c1 sky130_fd_pr__model__parasitic__diode_ps2nw_noresistor area={area}
dp p1 c1 sky130_fd_pr__model__parasitic__diode_ps2nw_noresistor area=1.0e-18
.ends sky130_fd_pr__model__parasitic__rf_diode_ps2nw
