* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 11
.param
+  sky130_fd_pr__nfet_05v0_nvt__toxe_mult=0.948
+  sky130_fd_pr__nfet_05v0_nvt__rshn_mult=1.0
+  sky130_fd_pr__nfet_05v0_nvt__overlap_mult=4.0927e-1
+  sky130_fd_pr__nfet_05v0_nvt__ajunction_mult=5.6418e-1
+  sky130_fd_pr__nfet_05v0_nvt__pjunction_mult=8.4099e-1
+  sky130_fd_pr__nfet_05v0_nvt__lint_diff=1.7325e-8
+  sky130_fd_pr__nfet_05v0_nvt__wint_diff=-3.2175e-8
+  sky130_fd_pr__nfet_05v0_nvt__dlc_diff=3.0000e-8
+  sky130_fd_pr__nfet_05v0_nvt__dwc_diff=-3.2175e-8
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 000, W = 10.0, L = 2.0
* -------------------------------------
+  sky130_fd_pr__nfet_05v0_nvt__eta0_diff_0=0.0
+  sky130_fd_pr__nfet_05v0_nvt__pdits_diff_0=0.0
+  sky130_fd_pr__nfet_05v0_nvt__keta_diff_0=0.0
+  sky130_fd_pr__nfet_05v0_nvt__kt1_diff_0=0.0
+  sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_0=0.0
+  sky130_fd_pr__nfet_05v0_nvt__pclm_diff_0=0.0
+  sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_0=0.084235
+  sky130_fd_pr__nfet_05v0_nvt__a0_diff_0=-0.088752
+  sky130_fd_pr__nfet_05v0_nvt__voff_diff_0=0.0
+  sky130_fd_pr__nfet_05v0_nvt__b0_diff_0=0.0
+  sky130_fd_pr__nfet_05v0_nvt__k2_diff_0=-0.00071772
+  sky130_fd_pr__nfet_05v0_nvt__u0_diff_0=-0.010239
+  sky130_fd_pr__nfet_05v0_nvt__ua_diff_0=-3.0465e-11
+  sky130_fd_pr__nfet_05v0_nvt__vsat_diff_0=0.0
+  sky130_fd_pr__nfet_05v0_nvt__vth0_diff_0=-0.042356
+  sky130_fd_pr__nfet_05v0_nvt__b1_diff_0=0.0
+  sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_0=0.0
+  sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_0=0.0
+  sky130_fd_pr__nfet_05v0_nvt__ags_diff_0=-0.0089574
+  sky130_fd_pr__nfet_05v0_nvt__ub_diff_0=-1.6353e-18
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 001, W = 10.0, L = 4.0
* -------------------------------------
+  sky130_fd_pr__nfet_05v0_nvt__ub_diff_1=-1.3876e-18
+  sky130_fd_pr__nfet_05v0_nvt__eta0_diff_1=0.0
+  sky130_fd_pr__nfet_05v0_nvt__pdits_diff_1=0.0
+  sky130_fd_pr__nfet_05v0_nvt__keta_diff_1=0.0
+  sky130_fd_pr__nfet_05v0_nvt__kt1_diff_1=0.0
+  sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_1=0.0
+  sky130_fd_pr__nfet_05v0_nvt__pclm_diff_1=0.0
+  sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_1=-0.036725
+  sky130_fd_pr__nfet_05v0_nvt__a0_diff_1=-0.051834
+  sky130_fd_pr__nfet_05v0_nvt__voff_diff_1=0.0
+  sky130_fd_pr__nfet_05v0_nvt__b0_diff_1=0.0
+  sky130_fd_pr__nfet_05v0_nvt__k2_diff_1=-0.0056229
+  sky130_fd_pr__nfet_05v0_nvt__u0_diff_1=-0.0086911
+  sky130_fd_pr__nfet_05v0_nvt__ua_diff_1=-2.5597e-11
+  sky130_fd_pr__nfet_05v0_nvt__vsat_diff_1=0.0
+  sky130_fd_pr__nfet_05v0_nvt__vth0_diff_1=-0.025235
+  sky130_fd_pr__nfet_05v0_nvt__b1_diff_1=0.0
+  sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_1=0.0
+  sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_1=0.0
+  sky130_fd_pr__nfet_05v0_nvt__ags_diff_1=-0.0075728
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 002, W = 10.0, L = 0.9
* -------------------------------------
+  sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_2=0.0
+  sky130_fd_pr__nfet_05v0_nvt__ags_diff_2=0.0
+  sky130_fd_pr__nfet_05v0_nvt__ub_diff_2=-1.9312e-18
+  sky130_fd_pr__nfet_05v0_nvt__eta0_diff_2=0.0
+  sky130_fd_pr__nfet_05v0_nvt__pdits_diff_2=0.0
+  sky130_fd_pr__nfet_05v0_nvt__keta_diff_2=0.0
+  sky130_fd_pr__nfet_05v0_nvt__kt1_diff_2=0.0
+  sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_2=0.0
+  sky130_fd_pr__nfet_05v0_nvt__pclm_diff_2=0.0
+  sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_2=0.12544
+  sky130_fd_pr__nfet_05v0_nvt__a0_diff_2=0.0
+  sky130_fd_pr__nfet_05v0_nvt__voff_diff_2=0.0
+  sky130_fd_pr__nfet_05v0_nvt__b0_diff_2=0.0
+  sky130_fd_pr__nfet_05v0_nvt__k2_diff_2=0.00061719
+  sky130_fd_pr__nfet_05v0_nvt__u0_diff_2=-0.011151
+  sky130_fd_pr__nfet_05v0_nvt__ua_diff_2=-4.1518e-11
+  sky130_fd_pr__nfet_05v0_nvt__vsat_diff_2=-7949.5
+  sky130_fd_pr__nfet_05v0_nvt__vth0_diff_2=0.024064
+  sky130_fd_pr__nfet_05v0_nvt__b1_diff_2=0.0
+  sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_2=0.0
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 003, W = 1.0, L = 25.0
* -------------------------------------
+  sky130_fd_pr__nfet_05v0_nvt__b1_diff_3=0.0
+  sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_3=0.0
+  sky130_fd_pr__nfet_05v0_nvt__ua_diff_3=-1.9154e-11
+  sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_3=0.0
+  sky130_fd_pr__nfet_05v0_nvt__ags_diff_3=-0.0071658
+  sky130_fd_pr__nfet_05v0_nvt__ub_diff_3=-1.1337e-18
+  sky130_fd_pr__nfet_05v0_nvt__eta0_diff_3=0.0
+  sky130_fd_pr__nfet_05v0_nvt__pdits_diff_3=0.0
+  sky130_fd_pr__nfet_05v0_nvt__keta_diff_3=0.0
+  sky130_fd_pr__nfet_05v0_nvt__kt1_diff_3=0.0
+  sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_3=0.0
+  sky130_fd_pr__nfet_05v0_nvt__pclm_diff_3=0.0
+  sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_3=0.010177
+  sky130_fd_pr__nfet_05v0_nvt__a0_diff_3=0.0013249
+  sky130_fd_pr__nfet_05v0_nvt__voff_diff_3=0.0
+  sky130_fd_pr__nfet_05v0_nvt__b0_diff_3=0.0
+  sky130_fd_pr__nfet_05v0_nvt__k2_diff_3=-0.0054271
+  sky130_fd_pr__nfet_05v0_nvt__u0_diff_3=-0.0080273
+  sky130_fd_pr__nfet_05v0_nvt__vsat_diff_3=0.0
+  sky130_fd_pr__nfet_05v0_nvt__vth0_diff_3=-0.029234
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 004, W = 1.0, L = 2.0
* ------------------------------------
+  sky130_fd_pr__nfet_05v0_nvt__u0_diff_4=-0.010027
+  sky130_fd_pr__nfet_05v0_nvt__vsat_diff_4=0.0
+  sky130_fd_pr__nfet_05v0_nvt__vth0_diff_4=-0.026425
+  sky130_fd_pr__nfet_05v0_nvt__b1_diff_4=0.0
+  sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_4=0.0
+  sky130_fd_pr__nfet_05v0_nvt__ua_diff_4=-2.2287e-11
+  sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_4=0.0
+  sky130_fd_pr__nfet_05v0_nvt__ags_diff_4=-0.068222
+  sky130_fd_pr__nfet_05v0_nvt__eta0_diff_4=0.0
+  sky130_fd_pr__nfet_05v0_nvt__ub_diff_4=-1.4787e-18
+  sky130_fd_pr__nfet_05v0_nvt__pdits_diff_4=0.0
+  sky130_fd_pr__nfet_05v0_nvt__keta_diff_4=0.0
+  sky130_fd_pr__nfet_05v0_nvt__kt1_diff_4=0.0
+  sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_4=0.0
+  sky130_fd_pr__nfet_05v0_nvt__pclm_diff_4=0.0
+  sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_4=-0.079945
+  sky130_fd_pr__nfet_05v0_nvt__a0_diff_4=-0.33061
+  sky130_fd_pr__nfet_05v0_nvt__voff_diff_4=0.0
+  sky130_fd_pr__nfet_05v0_nvt__b0_diff_4=0.0
+  sky130_fd_pr__nfet_05v0_nvt__k2_diff_4=-0.0024831
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 005, W = 1.0, L = 4.0
* ------------------------------------
+  sky130_fd_pr__nfet_05v0_nvt__b0_diff_5=0.0
+  sky130_fd_pr__nfet_05v0_nvt__k2_diff_5=-0.0012384
+  sky130_fd_pr__nfet_05v0_nvt__u0_diff_5=-0.009243
+  sky130_fd_pr__nfet_05v0_nvt__vsat_diff_5=0.0
+  sky130_fd_pr__nfet_05v0_nvt__vth0_diff_5=-0.023314
+  sky130_fd_pr__nfet_05v0_nvt__b1_diff_5=0.0
+  sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_5=0.0
+  sky130_fd_pr__nfet_05v0_nvt__ua_diff_5=-2.3342e-11
+  sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_5=0.0
+  sky130_fd_pr__nfet_05v0_nvt__ags_diff_5=-0.017982
+  sky130_fd_pr__nfet_05v0_nvt__eta0_diff_5=0.0
+  sky130_fd_pr__nfet_05v0_nvt__ub_diff_5=-1.3625e-18
+  sky130_fd_pr__nfet_05v0_nvt__pdits_diff_5=0.0
+  sky130_fd_pr__nfet_05v0_nvt__keta_diff_5=0.0
+  sky130_fd_pr__nfet_05v0_nvt__kt1_diff_5=0.0
+  sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_5=0.0
+  sky130_fd_pr__nfet_05v0_nvt__pclm_diff_5=0.0
+  sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_5=-0.012283
+  sky130_fd_pr__nfet_05v0_nvt__a0_diff_5=-0.089312
+  sky130_fd_pr__nfet_05v0_nvt__voff_diff_5=0.0
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 006, W = 1.0, L = 8.0
* ------------------------------------
+  sky130_fd_pr__nfet_05v0_nvt__voff_diff_6=0.0
+  sky130_fd_pr__nfet_05v0_nvt__a0_diff_6=-0.072963
+  sky130_fd_pr__nfet_05v0_nvt__b0_diff_6=0.0
+  sky130_fd_pr__nfet_05v0_nvt__k2_diff_6=-0.0029725
+  sky130_fd_pr__nfet_05v0_nvt__u0_diff_6=-0.0083572
+  sky130_fd_pr__nfet_05v0_nvt__vsat_diff_6=0.0
+  sky130_fd_pr__nfet_05v0_nvt__vth0_diff_6=-0.029505
+  sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_6=0.0
+  sky130_fd_pr__nfet_05v0_nvt__ua_diff_6=-2.0886e-11
+  sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_6=0.0
+  sky130_fd_pr__nfet_05v0_nvt__b1_diff_6=0.0
+  sky130_fd_pr__nfet_05v0_nvt__ags_diff_6=-0.013959
+  sky130_fd_pr__nfet_05v0_nvt__eta0_diff_6=0.0
+  sky130_fd_pr__nfet_05v0_nvt__ub_diff_6=-1.2199e-18
+  sky130_fd_pr__nfet_05v0_nvt__pdits_diff_6=0.0
+  sky130_fd_pr__nfet_05v0_nvt__keta_diff_6=0.0
+  sky130_fd_pr__nfet_05v0_nvt__kt1_diff_6=0.0
+  sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_6=0.0
+  sky130_fd_pr__nfet_05v0_nvt__pclm_diff_6=0.0
+  sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_6=-0.042692
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 007, W = 1.0, L = 0.9
* ------------------------------------
+  sky130_fd_pr__nfet_05v0_nvt__kt1_diff_7=0.0
+  sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_7=0.0
+  sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_7=0.079414
+  sky130_fd_pr__nfet_05v0_nvt__voff_diff_7=0.0
+  sky130_fd_pr__nfet_05v0_nvt__a0_diff_7=0.0
+  sky130_fd_pr__nfet_05v0_nvt__b0_diff_7=0.0
+  sky130_fd_pr__nfet_05v0_nvt__k2_diff_7=-8.6129e-5
+  sky130_fd_pr__nfet_05v0_nvt__u0_diff_7=-0.012564
+  sky130_fd_pr__nfet_05v0_nvt__vth0_diff_7=-0.049862
+  sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_7=0.0
+  sky130_fd_pr__nfet_05v0_nvt__ua_diff_7=-3.2654e-11
+  sky130_fd_pr__nfet_05v0_nvt__vsat_diff_7=-9440.5
+  sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_7=0.0
+  sky130_fd_pr__nfet_05v0_nvt__b1_diff_7=0.0
+  sky130_fd_pr__nfet_05v0_nvt__ags_diff_7=0.0
+  sky130_fd_pr__nfet_05v0_nvt__eta0_diff_7=0.0
+  sky130_fd_pr__nfet_05v0_nvt__ub_diff_7=-1.7558e-18
+  sky130_fd_pr__nfet_05v0_nvt__pdits_diff_7=0.0
+  sky130_fd_pr__nfet_05v0_nvt__keta_diff_7=0.0
+  sky130_fd_pr__nfet_05v0_nvt__pclm_diff_7=0.0
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 008, W = 0.42, L = 1.0
* -------------------------------------
+  sky130_fd_pr__nfet_05v0_nvt__pclm_diff_8=0.0
+  sky130_fd_pr__nfet_05v0_nvt__kt1_diff_8=0.0
+  sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_8=0.0
+  sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_8=0.050854
+  sky130_fd_pr__nfet_05v0_nvt__voff_diff_8=0.0
+  sky130_fd_pr__nfet_05v0_nvt__a0_diff_8=0.0
+  sky130_fd_pr__nfet_05v0_nvt__b0_diff_8=2.7274e-7
+  sky130_fd_pr__nfet_05v0_nvt__k2_diff_8=-0.011083
+  sky130_fd_pr__nfet_05v0_nvt__u0_diff_8=-0.012082
+  sky130_fd_pr__nfet_05v0_nvt__vth0_diff_8=-0.068342
+  sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_8=0.0
+  sky130_fd_pr__nfet_05v0_nvt__ua_diff_8=-2.1309e-11
+  sky130_fd_pr__nfet_05v0_nvt__vsat_diff_8=0.0
+  sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_8=0.0
+  sky130_fd_pr__nfet_05v0_nvt__b1_diff_8=-2.2962e-8
+  sky130_fd_pr__nfet_05v0_nvt__ags_diff_8=0.0
+  sky130_fd_pr__nfet_05v0_nvt__eta0_diff_8=0.0
+  sky130_fd_pr__nfet_05v0_nvt__ub_diff_8=-1.6897e-18
+  sky130_fd_pr__nfet_05v0_nvt__pdits_diff_8=0.0
+  sky130_fd_pr__nfet_05v0_nvt__keta_diff_8=0.0
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 009, W = 0.42, L = 0.9
* -------------------------------------
+  sky130_fd_pr__nfet_05v0_nvt__pdits_diff_9=0.0
+  sky130_fd_pr__nfet_05v0_nvt__keta_diff_9=0.0
+  sky130_fd_pr__nfet_05v0_nvt__pclm_diff_9=0.0
+  sky130_fd_pr__nfet_05v0_nvt__kt1_diff_9=0.0
+  sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_9=0.0
+  sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_9=-0.15711
+  sky130_fd_pr__nfet_05v0_nvt__voff_diff_9=0.0
+  sky130_fd_pr__nfet_05v0_nvt__a0_diff_9=0.0
+  sky130_fd_pr__nfet_05v0_nvt__b0_diff_9=0.0
+  sky130_fd_pr__nfet_05v0_nvt__k2_diff_9=-0.0083374
+  sky130_fd_pr__nfet_05v0_nvt__u0_diff_9=-0.012537
+  sky130_fd_pr__nfet_05v0_nvt__vth0_diff_9=-0.057364
+  sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_9=0.0
+  sky130_fd_pr__nfet_05v0_nvt__ua_diff_9=-1.3616e-10
+  sky130_fd_pr__nfet_05v0_nvt__vsat_diff_9=-13432.0
+  sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_9=0.0
+  sky130_fd_pr__nfet_05v0_nvt__b1_diff_9=0.0
+  sky130_fd_pr__nfet_05v0_nvt__ags_diff_9=0.0
+  sky130_fd_pr__nfet_05v0_nvt__eta0_diff_9=0.0
+  sky130_fd_pr__nfet_05v0_nvt__ub_diff_9=-1.1456e-18
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 010, W = 0.7, L = 0.9
* ------------------------------------
+  sky130_fd_pr__nfet_05v0_nvt__vsat_diff_10=-11514.0
+  sky130_fd_pr__nfet_05v0_nvt__vth0_diff_10=-0.047797
+  sky130_fd_pr__nfet_05v0_nvt__b0_diff_10=0.0
+  sky130_fd_pr__nfet_05v0_nvt__keta_diff_10=0.0
+  sky130_fd_pr__nfet_05v0_nvt__b1_diff_10=0.0
+  sky130_fd_pr__nfet_05v0_nvt__kt1_diff_10=0.0
+  sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_10=0.0
+  sky130_fd_pr__nfet_05v0_nvt__pclm_diff_10=0.0
+  sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_10=0.058
+  sky130_fd_pr__nfet_05v0_nvt__ags_diff_10=0.0
+  sky130_fd_pr__nfet_05v0_nvt__u0_diff_10=-0.012559
+  sky130_fd_pr__nfet_05v0_nvt__pdits_diff_10=0.0
+  sky130_fd_pr__nfet_05v0_nvt__k2_diff_10=0.0004686
+  sky130_fd_pr__nfet_05v0_nvt__ua_diff_10=-2.9266e-11
+  sky130_fd_pr__nfet_05v0_nvt__eta0_diff_10=0.0
+  sky130_fd_pr__nfet_05v0_nvt__ub_diff_10=-1.7087e-18
+  sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_10=0.0
+  sky130_fd_pr__nfet_05v0_nvt__voff_diff_10=0.0
+  sky130_fd_pr__nfet_05v0_nvt__a0_diff_10=0.0
+  sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_10=0.0
.include "sky130_fd_pr__nfet_05v0_nvt.pm3.spice"
