* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 49
.param
+  sky130_fd_pr__nfet_g5v0d10v5__toxe_mult=0.958
+  sky130_fd_pr__nfet_g5v0d10v5__rshn_mult=1.0
+  sky130_fd_pr__nfet_g5v0d10v5__overlap_mult=0.80232
+  sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult=8.7078e-1
+  sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult=8.4883e-1
+  sky130_fd_pr__nfet_g5v0d10v5__lint_diff=1.21275e-8
+  sky130_fd_pr__nfet_g5v0d10v5__wint_diff=-2.252e-8
+  sky130_fd_pr__nfet_g5v0d10v5__dlc_diff=1.21275e-8
+  sky130_fd_pr__nfet_g5v0d10v5__dwc_diff=-2.252e-8
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 000, W = 10.0, L = 0.5
* -------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_0=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_0=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_0=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_0=-0.0027974
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_0=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_0=0.0028713
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_0=-0.088847
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_0=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_0=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_0=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_0=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_0=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_0=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_0=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_0=-3.182e-12
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_0=-7539.2
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_0=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_0=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_0=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_0=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_0=0.067831
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_0=-1.431e-20
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_0=0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 001, W = 15.0, L = 1.0
* -------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_1=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_1=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_1=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_1=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_1=0.0057654
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_1=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_1=0.00045135
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_1=-0.034563
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_1=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_1=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_1=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_1=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_1=-0.12355
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_1=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_1=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_1=-5.9724e-12
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_1=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_1=0.065625
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_1=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_1=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_1=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_1=0.23772
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_1=-5.0923e-19
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 002, W = 15.0, L = 0.5
* -------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_2=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_2=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_2=0.061219
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_2=-1.2189e-19
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_2=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_2=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_2=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_2=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_2=-0.0035133
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_2=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_2=0.0040354
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_2=-0.077042
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_2=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_2=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_2=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_2=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_2=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_2=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_2=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_2=-1.0836e-11
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_2=-3684.4
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_2=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_2=0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 003, W = 1.5, L = 1.0
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_3=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_3=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_3=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_3=0.42574
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_3=-2.6147e-19
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_3=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_3=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_3=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_3=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_3=-0.0027391
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_3=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_3=-0.0016864
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_3=-0.061437
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_3=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_3=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_3=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_3=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_3=-0.065837
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_3=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_3=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_3=1.7763e-12
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_3=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_3=0.019369
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 004, W = 1.5, L = 2.0
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_4=-0.0028111
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_4=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_4=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_4=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_4=0.40835
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_4=-2.1584e-19
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_4=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_4=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_4=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_4=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_4=-0.012463
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_4=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_4=-0.0013555
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_4=-0.040788
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_4=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_4=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_4=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_4=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_4=-0.0049408
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_4=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_4=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_4=1.3358e-12
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_4=0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 005, W = 1.5, L = 4.0
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_5=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_5=3.462e-13
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_5=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_5=0.056417
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_5=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_5=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_5=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_5=-1.1837e-19
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_5=0.46504
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_5=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_5=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_5=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_5=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_5=-0.015753
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_5=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_5=-0.00055717
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_5=-0.024671
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_5=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_5=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_5=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_5=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_5=-0.0048985
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_5=0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 006, W = 1.5, L = 0.5
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_6=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_6=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_6=2.2098e-12
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_6=-12771.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_6=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_6=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_6=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_6=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_6=2.0562e-19
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_6=0.5662
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_6=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_6=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_6=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_6=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_6=0.0064292
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_6=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_6=0.00046466
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_6=-0.11792
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_6=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_6=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_6=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_6=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_6=0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 007, W = 1.0, L = 1.0
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_7=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_7=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_7=-0.070162
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_7=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_7=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_7=1.8609e-13
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_7=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_7=0.018372
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_7=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_7=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_7=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_7=1.1345e-19
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_7=0.47052
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_7=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_7=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_7=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_7=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_7=0.0070682
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_7=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_7=0.00067424
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_7=-0.053375
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_7=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_7=0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 008, W = 1.0, L = 2.0
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_8=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_8=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_8=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_8=-0.02736
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_8=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_8=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_8=-3.4817e-13
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_8=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_8=0.0022824
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_8=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_8=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_8=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_8=7.1857e-20
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_8=0.47872
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_8=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_8=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_8=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_8=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_8=-0.017505
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_8=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_8=0.00056754
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_8=-0.037424
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_8=0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 009, W = 1.0, L = 4.0
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_9=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_9=-3.1448e-5
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_9=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_9=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_9=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_9=-0.039057
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_9=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_9=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_9=-1.1637e-12
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_9=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_9=0.0044918
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_9=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_9=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_9=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_9=-1.0967e-19
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_9=0.47982
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_9=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_9=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_9=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_9=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_9=-0.01097
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_9=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_9=-0.028174
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 010, W = 1.0, L = 8.0
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_10=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_10=0.0020684
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_10=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_10=0.00054307
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_10=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_10=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_10=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_10=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_10=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_10=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_10=-0.014456
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_10=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_10=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_10=-0.026085
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_10=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_10=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_10=-0.012853
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_10=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_10=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_10=0.58337
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_10=-1.0424e-12
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_10=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_10=6.9348e-20
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 011, W = 1.0, L = 0.5
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_11=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_11=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_11=5.8398e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_11=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_11=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_11=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_11=0.00087252
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_11=-11273.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_11=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_11=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_11=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_11=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_11=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_11=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_11=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_11=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_11=-0.098283
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_11=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_11=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_11=0.009725
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_11=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_11=0.64332
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_11=5.7181e-12
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 012, W = 1.0, L = 0.6
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_12=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_12=0.56622
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_12=2.5824e-13
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_12=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_12=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_12=2.189e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_12=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_12=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_12=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_12=0.0013169
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_12=-12347.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_12=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_12=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_12=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_12=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_12=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_12=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_12=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_12=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_12=-0.078832
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_12=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_12=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_12=-6.4922e-5
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 013, W = 1.0, L = 0.8
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_13=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_13=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_13=-0.0037695
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_13=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_13=0.48453
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_13=1.0279e-12
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_13=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_13=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_13=1.6812e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_13=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_13=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_13=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_13=0.00063843
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_13=-10586.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_13=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_13=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_13=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_13=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_13=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_13=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_13=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_13=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_13=-0.040366
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 014, W = 20.0, L = 1.0
* -------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_14=-0.030427
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_14=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_14=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_14=0.0052638
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_14=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_14=0.23489
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_14=-1.5158e-12
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_14=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_14=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_14=-5.2955e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_14=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_14=0.015139
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_14=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_14=0.00080727
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_14=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_14=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_14=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_14=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_14=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_14=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_14=-0.035603
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_14=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_14=0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 015, W = 20.0, L = 0.5
* -------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_15=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_15=-0.077885
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_15=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_15=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_15=-0.00642
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_15=-0.0080405
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_15=-3.4099e-12
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_15=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_15=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_15=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_15=-1.0702e-18
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_15=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_15=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_15=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_15=0.00091931
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_15=-9206.5
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_15=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_15=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_15=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_15=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_15=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_15=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_15=0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 016, W = 3.0, L = 1.0
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_16=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_16=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_16=-0.041274
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_16=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_16=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_16=-0.0037619
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_16=0.31557
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_16=1.7658e-12
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_16=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_16=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_16=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_16=-2.2493e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_16=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_16=0.020382
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_16=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_16=-0.0014343
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_16=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_16=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_16=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_16=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_16=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_16=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_16=-0.065114
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 017, W = 3.0, L = 2.0
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_17=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_17=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_17=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_17=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_17=-0.031553
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_17=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_17=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_17=-0.03465
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_17=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_17=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_17=-0.012842
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_17=0.31329
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_17=9.6403e-13
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_17=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_17=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_17=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_17=-1.9267e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_17=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_17=0.0035437
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_17=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_17=-0.0010807
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_17=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_17=0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 018, W = 3.0, L = 4.0
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_18=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_18=-0.0010212
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_18=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_18=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_18=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_18=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_18=-0.0060841
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_18=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_18=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_18=-0.026041
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_18=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_18=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_18=-0.017484
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_18=0.38531
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_18=7.0524e-13
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_18=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_18=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_18=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_18=-1.7595e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_18=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_18=-0.00075152
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_18=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_18=0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 019, W = 3.0, L = 8.0
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_19=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_19=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_19=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_19=-0.00069241
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_19=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_19=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_19=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_19=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_19=-0.0036221
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_19=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_19=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_19=-0.027928
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_19=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_19=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_19=-0.019581
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_19=0.42719
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_19=7.685e-13
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_19=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_19=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_19=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_19=-7.8066e-20
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_19=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_19=-0.00099191
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 020, W = 3.0, L = 0.5
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_20=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_20=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_20=0.0013
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_20=-7459.6
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_20=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_20=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_20=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_20=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_20=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_20=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_20=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_20=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_20=-0.083823
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_20=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_20=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_20=0.00020718
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_20=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_20=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_20=0.37831
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_20=1.0967e-12
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_20=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_20=3.1912e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_20=0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 021, W = 3.0, L = 0.6
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_21=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_21=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_21=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_21=0.0016329
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_21=-8092.6
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_21=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_21=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_21=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_21=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_21=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_21=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_21=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_21=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_21=-0.046029
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_21=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_21=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_21=-0.0043173
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_21=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_21=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_21=0.29359
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_21=4.4953e-13
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_21=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_21=3.6335e-19
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 022, W = 5.0, L = 1.0
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_22=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_22=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_22=-2.0321e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_22=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_22=0.01461
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_22=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_22=-0.00057883
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_22=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_22=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_22=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_22=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_22=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_22=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_22=-0.052098
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_22=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_22=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_22=-0.042799
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_22=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_22=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_22=0.0070137
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_22=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_22=0.2603
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_22=5.116e-13
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 023, W = 5.0, L = 2.0
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_23=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_23=0.31947
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_23=2.5465e-12
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_23=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_23=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_23=-2.8995e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_23=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_23=-0.0029884
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_23=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_23=-0.0020677
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_23=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_23=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_23=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_23=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_23=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_23=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_23=-0.0011022
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_23=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_23=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_23=-0.032747
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_23=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_23=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_23=-0.003602
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 024, W = 5.0, L = 4.0
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_24=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_24=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_24=-0.0074643
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_24=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_24=0.37028
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_24=2.221e-12
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_24=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_24=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_24=-3.6366e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_24=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_24=-0.0010324
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_24=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_24=-0.0022597
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_24=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_24=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_24=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_24=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_24=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_24=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_24=-0.0052798
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_24=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_24=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_24=-0.027581
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 025, W = 5.0, L = 8.0
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_25=-0.022259
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_25=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_25=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_25=-0.010119
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_25=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_25=0.41609
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_25=2.2767e-12
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_25=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_25=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_25=-2.7467e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_25=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_25=-0.0009647
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_25=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_25=-0.0020508
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_25=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_25=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_25=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_25=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_25=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_25=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_25=0.00032626
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_25=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_25=0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 026, W = 5.0, L = 0.5
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_26=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_26=-0.086548
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_26=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_26=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_26=-0.0050158
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_26=0.2557
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_26=-1.161e-12
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_26=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_26=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_26=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_26=3.2723e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_26=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_26=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_26=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_26=0.0021239
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_26=-6995.1
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_26=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_26=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_26=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_26=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_26=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_26=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_26=0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 027, W = 5.0, L = 0.6
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_27=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_27=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_27=-0.038139
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_27=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_27=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_27=0.0032747
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_27=0.25608
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_27=-1.5018e-12
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_27=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_27=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_27=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_27=3.0302e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_27=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_27=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_27=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_27=0.0020646
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_27=-6597.3
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_27=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_27=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_27=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_27=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_27=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_27=0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 028, W = 5.0, L = 0.8
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_28=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_28=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_28=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_28=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_28=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_28=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_28=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_28=-0.044634
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_28=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_28=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_28=0.0096143
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_28=0.25408
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_28=-9.9611e-14
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_28=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_28=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_28=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_28=-6.4691e-20
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_28=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_28=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_28=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_28=-2.5118e-5
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_28=-6227.3
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_28=0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 029, W = 7.0, L = 1.0
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_29=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_29=-0.0018504
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_29=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_29=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_29=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_29=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_29=-0.05638
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_29=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_29=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_29=-0.044064
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_29=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_29=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_29=0.0063314
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_29=0.25044
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_29=1.2724e-12
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_29=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_29=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_29=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_29=-3.9876e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_29=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_29=0.014604
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_29=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_29=0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 030, W = 7.0, L = 2.0
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_30=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_30=-0.002852
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_30=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_30=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_30=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_30=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_30=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_30=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_30=-0.010921
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_30=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_30=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_30=-0.033936
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_30=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_30=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_30=-0.0035423
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_30=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_30=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_30=0.30296
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_30=2.8109e-12
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_30=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_30=-4.8973e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_30=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_30=-0.00078965
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 031, W = 7.0, L = 4.0
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_31=-0.00046676
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_31=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_31=-0.0024131
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_31=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_31=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_31=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_31=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_31=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_31=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_31=-0.0083154
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_31=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_31=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_31=-0.028874
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_31=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_31=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_31=-0.008373
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_31=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_31=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_31=0.3483
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_31=2.1907e-12
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_31=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_31=-4.138e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_31=0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 032, W = 7.0, L = 8.0
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_32=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_32=-0.0012569
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_32=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_32=-0.0023959
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_32=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_32=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_32=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_32=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_32=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_32=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_32=-0.0013673
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_32=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_32=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_32=-0.025062
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_32=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_32=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_32=-0.0096443
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_32=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_32=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_32=0.38967
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_32=2.6931e-12
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_32=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_32=-3.5024e-19
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 033, W = 7.0, L = 0.5
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_33=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_33=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_33=3.7315e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_33=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_33=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_33=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_33=0.0029548
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_33=-4708.3
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_33=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_33=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_33=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_33=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_33=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_33=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_33=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_33=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_33=-0.087831
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_33=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_33=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_33=-0.0049325
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_33=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_33=0.13655
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_33=-2.4379e-12
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 034, W = 7.0, L = 0.8
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_34=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_34=0.24119
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_34=7.0668e-14
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_34=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_34=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_34=-3.9044e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_34=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_34=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_34=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_34=-0.0014463
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_34=-8550.4
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_34=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_34=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_34=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_34=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_34=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_34=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_34=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_34=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_34=-0.041196
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_34=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_34=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_34=0.0089142
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 035, W = 0.42, L = 1.0
* -------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_35=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_35=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_35=-0.010696
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_35=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_35=0.34258
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_35=3.9893e-12
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_35=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_35=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_35=2.8144e-20
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_35=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_35=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_35=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_35=-0.00078634
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_35=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_35=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_35=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_35=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_35=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_35=1.6359e-7
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_35=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_35=3.2317e-9
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_35=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_35=-0.0987
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 036, W = 0.42, L = 20.0
* --------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_36=-0.050867
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_36=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_36=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_36=-0.014717
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_36=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_36=0.84261
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_36=4.2528e-12
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_36=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_36=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_36=-1.3575e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_36=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_36=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_36=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_36=-0.0017002
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_36=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_36=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_36=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_36=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_36=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_36=4.3021e-8
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_36=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_36=1.6373e-8
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_36=0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 037, W = 0.42, L = 2.0
* -------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_37=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_37=-0.054153
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_37=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_37=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_37=-0.015653
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_37=0.46203
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_37=6.6845e-13
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_37=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_37=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_37=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_37=-8.5678e-20
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_37=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_37=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_37=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_37=-0.00033292
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_37=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_37=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_37=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_37=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_37=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_37=5.2233e-8
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_37=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_37=1.0156e-8
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 038, W = 0.42, L = 4.0
* -------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_38=1.6953e-9
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_38=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_38=-0.056807
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_38=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_38=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_38=-0.012851
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_38=0.51933
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_38=5.1331e-12
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_38=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_38=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_38=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_38=-1.2021e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_38=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_38=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_38=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_38=-0.0020417
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_38=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_38=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_38=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_38=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_38=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_38=2.3908e-8
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_38=0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 039, W = 0.42, L = 8.0
* -------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_39=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_39=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_39=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_39=3.1542e-8
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_39=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_39=2.0388e-11
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_39=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_39=-0.056058
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_39=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_39=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_39=-0.016471
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_39=0.66375
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_39=3.7681e-12
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_39=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_39=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_39=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_39=-3.1135e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_39=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_39=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_39=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_39=-0.0020927
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_39=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_39=0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 040, W = 0.42, L = 0.5
* -------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_40=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_40=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_40=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_40=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_40=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_40=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_40=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_40=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_40=-0.10791
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_40=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_40=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_40=0.00018191
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_40=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_40=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_40=0.56496
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_40=-6.008e-13
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_40=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_40=1.1662e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_40=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_40=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_40=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_40=0.00080213
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_40=-15876.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 041, W = 0.42, L = 0.6
* -------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_41=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_41=0.00068511
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_41=-14626.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_41=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_41=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_41=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_41=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_41=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_41=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_41=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_41=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_41=-0.10296
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_41=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_41=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_41=-0.013171
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_41=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_41=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_41=0.43908
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_41=-2.223e-13
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_41=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_41=2.9418e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_41=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_41=0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 042, W = 0.42, L = 0.8
* -------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_42=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_42=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_42=0.00071959
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_42=-10576.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_42=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_42=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_42=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_42=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_42=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_42=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_42=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_42=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_42=-0.11458
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_42=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_42=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_42=-0.019163
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_42=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_42=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_42=0.41785
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_42=3.1011e-13
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_42=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_42=1.4931e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_42=0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 043, W = 0.75, L = 1.0
* -------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_43=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_43=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_43=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_43=0.00031538
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_43=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_43=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_43=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_43=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_43=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_43=1.1826e-7
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_43=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_43=3.1376e-10
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_43=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_43=-0.045571
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_43=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_43=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_43=-0.0033931
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_43=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_43=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_43=0.4774
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_43=7.6428e-13
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_43=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_43=9.6791e-20
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 044, W = 0.75, L = 2.0
* -------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_44=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_44=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_44=4.1633e-20
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_44=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_44=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_44=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_44=0.00052743
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_44=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_44=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_44=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_44=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_44=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_44=6.66e-8
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_44=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_44=3.5282e-11
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_44=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_44=-0.056435
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_44=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_44=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_44=-0.011972
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_44=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_44=0.4896
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_44=-8.2831e-14
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 045, W = 0.75, L = 4.0
* -------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_45=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_45=0.56435
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_45=-6.1055e-13
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_45=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_45=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_45=-1.8313e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_45=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_45=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_45=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_45=-0.00062318
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_45=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_45=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_45=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_45=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_45=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_45=1.133e-7
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_45=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_45=-3.2543e-11
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_45=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_45=-0.033666
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_45=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_45=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_45=-0.016427
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 046, W = 0.75, L = 0.5
* -------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_46=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_46=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_46=0.0018396
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_46=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_46=0.6137
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_46=4.3681e-12
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_46=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_46=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_46=5.9892e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_46=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_46=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_46=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_46=0.0014762
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_46=-11740.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_46=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_46=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_46=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_46=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_46=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_46=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_46=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_46=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_46=-0.097457
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 047, W = 0.75, L = 0.8
* -------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_47=-0.051222
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_47=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_47=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_47=-0.00044726
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_47=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_47=0.54901
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_47=-2.612e-13
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_47=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_47=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_47=8.7859e-20
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_47=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_47=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_47=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_47=0.00080669
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_47=-12361.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_47=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_47=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_47=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_47=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_47=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_47=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_47=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_47=0.0
*
* sky130_fd_pr__nfet_g5v0d10v5, Bin 048, W = 0.7, L = 0.6
* ------------------------------
+  sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_48=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_48=-0.076516
+  sky130_fd_pr__nfet_g5v0d10v5__keta_diff_48=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_48=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__k2_diff_48=0.00055257
+  sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_48=0.6225
+  sky130_fd_pr__nfet_g5v0d10v5__ua_diff_48=1.8742e-12
+  sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_48=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_48=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_48=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ub_diff_48=1.945e-19
+  sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_48=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__a0_diff_48=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_48=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__u0_diff_48=0.00058111
+  sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_48=-14997.0
+  sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_48=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_48=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_48=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__voff_diff_48=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b0_diff_48=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__ags_diff_48=0.0
+  sky130_fd_pr__nfet_g5v0d10v5__b1_diff_48=0.0
.include "sky130_fd_pr__nfet_g5v0d10v5.pm3.spice"
