* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* statistics {
*   mismatch {
*   }
* }
.subckt sky130_fd_pr__cap_vpp_08p6x07p8_m1m2_noshield c0 c1 b
.param mult=1 presim_flag=0.0
+  lvpp=7.06 wm1=0.14 wm2=0.14
+  ctot_a={35.0e-15*cvpp3_cor+0.0283/sqrt(7.84*8.58*2*mult)*35.0e-15*cvpp3_cor*sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_noshield_o1__generic_slope}
+  rat_m2=0.5767
+  rat_m1=0.4233
+  cap_m2={rat_m2*ctot_a}
+  cap_m1={rat_m1*ctot_a}
+  caps_m1={(1.65+presim_flag*0.19)*1e-15*cli2s_vpp}
+  nvia=47.0
+  nf=14.0
rm21 c0 a1 r={2*rm2*lvpp/wm2*(1/3)*(1/nf)}
ccmvpp3 a1 c1 c={cap_m2}
rvia1 c0 d0 r={rcvia/nvia}
rvia2 c1 d1 r={rcvia/nvia}
rm11 d0 b1 r={2*rm1*lvpp/wm1*(1/3)*(1/nf)}
cm1 b1 d1 c={cap_m1}
csli1 d0 b c={caps_m1}
csli2 d1 b c={caps_m1}
.ends sky130_fd_pr__cap_vpp_08p6x07p8_m1m2_noshield
