* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 8
.param
+  sky130_fd_pr__rf_pfet_01v8_b__toxe_mult=1.0365
+  sky130_fd_pr__rf_pfet_01v8_b__rbpb_mult=1.2
+  sky130_fd_pr__rf_pfet_01v8_b__overlap_mult=1.1043
+  sky130_fd_pr__rf_pfet_01v8_b__ajunction_mult=1.0625
+  sky130_fd_pr__rf_pfet_01v8_b__pjunction_mult=1.0675
+  sky130_fd_pr__rf_pfet_01v8_b__lint_diff=-1.21275e-8
+  sky130_fd_pr__rf_pfet_01v8_b__wint_diff=2.252e-8
+  sky130_fd_pr__rf_pfet_01v8_b__rshg_diff=7.0
+  sky130_fd_pr__rf_pfet_01v8_b__dlc_diff=-1.21275e-8
+  sky130_fd_pr__rf_pfet_01v8_b__dwc_diff=0.0
+  sky130_fd_pr__rf_pfet_01v8_b__xgw_diff=4.504e-8
+  sky130_fd_pr__rf_pfet_01v8__aw_cap_mult=1.1125
+  sky130_fd_pr__rf_pfet_01v8__aw_rgate_dist_mult=1.315
+  sky130_fd_pr__rf_pfet_01v8__aw_rgate_stub_mult=1.315
+  sky130_fd_pr__rf_pfet_01v8__aw_cap_mult_2=1.1125
+  sky130_fd_pr__rf_pfet_01v8__aw_rgate_dist_mult_2=1.21
+  sky130_fd_pr__rf_pfet_01v8__aw_rgate_stub_mult_2=1.21
+  sky130_fd_pr__rf_pfet_01v8__aw_rd_mult=1.0
+  sky130_fd_pr__rf_pfet_01v8__aw_rs_mult=1.0
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 000, W = 1.65, L = 0.15
* ------------------------------------------------
+  sky130_fd_pr__rf_pfet_01v8_bM02__rdsw_diff_0=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__ua_diff_0=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_0=-0.025683
+  sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_0=-0.00046629
+  sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_0=0.036263
+  sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_0=-4705.4
+  sky130_fd_pr__rf_pfet_01v8_bM02__b1_diff_0=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__kt1_diff_0=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__nfactor_diff_0=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__ub_diff_0=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__voff_diff_0=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__ags_diff_0=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__a0_diff_0=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__b0_diff_0=0.0
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 001, W = 1.65, L = 0.18
* ------------------------------------------------
+  sky130_fd_pr__rf_pfet_01v8_bM02__b0_diff_1=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__rdsw_diff_1=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__ua_diff_1=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_1=-0.0096007
+  sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_1=-0.00041939
+  sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_1=0.036542
+  sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_1=-19320.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__b1_diff_1=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__kt1_diff_1=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__nfactor_diff_1=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__ub_diff_1=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__voff_diff_1=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__ags_diff_1=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__a0_diff_1=0.0
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 002, W = 1.65, L = 0.25
* ------------------------------------------------
+  sky130_fd_pr__rf_pfet_01v8_bM02__voff_diff_2=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__ags_diff_2=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__a0_diff_2=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__b0_diff_2=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__ua_diff_2=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__rdsw_diff_2=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_2=-0.00361
+  sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_2=-0.000495
+  sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_2=0.022214
+  sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_2=-19622.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__b1_diff_2=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__kt1_diff_2=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__nfactor_diff_2=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__ub_diff_2=0.0
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 003, W = 3.01, L = 0.15
* ------------------------------------------------
+  sky130_fd_pr__rf_pfet_01v8_bM02__rdsw_diff_3=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__ua_diff_3=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_3=-0.02462
+  sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_3=-0.0008663
+  sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_3=0.054438
+  sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_3=-17486.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__b1_diff_3=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__kt1_diff_3=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__nfactor_diff_3=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__ub_diff_3=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__voff_diff_3=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__ags_diff_3=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__a0_diff_3=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__b0_diff_3=0.0
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 004, W = 3.01, L = 0.18
* ------------------------------------------------
+  sky130_fd_pr__rf_pfet_01v8_bM02__kt1_diff_4=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__nfactor_diff_4=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__ub_diff_4=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__voff_diff_4=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__ags_diff_4=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__a0_diff_4=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__b0_diff_4=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__ua_diff_4=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__rdsw_diff_4=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_4=-0.018152
+  sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_4=-0.00068712
+  sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_4=0.046452
+  sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_4=-11488.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__b1_diff_4=0.0
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 005, W = 3.01, L = 0.25
* ------------------------------------------------
+  sky130_fd_pr__rf_pfet_01v8_bM02__kt1_diff_5=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__nfactor_diff_5=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__ub_diff_5=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__ags_diff_5=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__a0_diff_5=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__voff_diff_5=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__b0_diff_5=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__ua_diff_5=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__rdsw_diff_5=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_5=-0.016536
+  sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_5=-0.00054677
+  sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_5=0.022396
+  sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_5=-14168.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__b1_diff_5=0.0
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 006, W = 5.05, L = 0.15
* ------------------------------------------------
+  sky130_fd_pr__rf_pfet_01v8_bM02__b1_diff_6=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__kt1_diff_6=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__nfactor_diff_6=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__ub_diff_6=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__ags_diff_6=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__a0_diff_6=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__voff_diff_6=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__b0_diff_6=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__ua_diff_6=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__rdsw_diff_6=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_6=-0.025252
+  sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_6=-0.0012477
+  sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_6=0.074957
+  sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_6=-15388.0
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 007, W = 5.05, L = 0.18
* ------------------------------------------------
+  sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_7=-0.0006238
+  sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_7=-19606.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__b1_diff_7=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__kt1_diff_7=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__ub_diff_7=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__nfactor_diff_7=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__ags_diff_7=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__a0_diff_7=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__voff_diff_7=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__b0_diff_7=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__ua_diff_7=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__rdsw_diff_7=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_7=-0.013565
+  sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_7=0.045593
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 008, W = 5.05, L = 0.25
* ------------------------------------------------
+  sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_8=0.026563
+  sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_8=-0.0006639
+  sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_8=-20194.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__b1_diff_8=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__kt1_diff_8=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__ub_diff_8=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__nfactor_diff_8=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__ags_diff_8=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__a0_diff_8=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__voff_diff_8=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__b0_diff_8=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__ua_diff_8=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__rdsw_diff_8=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_8=-0.013354
*
* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 000, W = 1.65, L = 0.15
* ------------------------------------------------
+  sky130_fd_pr__rf_pfet_01v8_bM04__b1_diff_0=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__ub_diff_0=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__rdsw_diff_0=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_0=-0.024438
+  sky130_fd_pr__rf_pfet_01v8_bM04__kt1_diff_0=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__nfactor_diff_0=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__voff_diff_0=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__ags_diff_0=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__a0_diff_0=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__b0_diff_0=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_0=-0.00066296
+  sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_0=0.049452
+  sky130_fd_pr__rf_pfet_01v8_bM04__ua_diff_0=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_0=-8761.9
*
* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 001, W = 1.65, L = 0.18
* ------------------------------------------------
+  sky130_fd_pr__rf_pfet_01v8_bM04__b1_diff_1=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__ub_diff_1=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__rdsw_diff_1=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_1=-0.0094416
+  sky130_fd_pr__rf_pfet_01v8_bM04__kt1_diff_1=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__nfactor_diff_1=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__voff_diff_1=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__ags_diff_1=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__a0_diff_1=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__b0_diff_1=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_1=-0.00051496
+  sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_1=0.050655
+  sky130_fd_pr__rf_pfet_01v8_bM04__ua_diff_1=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_1=-10144.0
*
* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 002, W = 1.65, L = 0.25
* ------------------------------------------------
+  sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_2=-0.00053393
+  sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_2=0.029231
+  sky130_fd_pr__rf_pfet_01v8_bM04__ua_diff_2=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_2=-14879.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__b1_diff_2=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__ub_diff_2=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__rdsw_diff_2=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_2=-0.0049051
+  sky130_fd_pr__rf_pfet_01v8_bM04__kt1_diff_2=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__nfactor_diff_2=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__voff_diff_2=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__ags_diff_2=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__a0_diff_2=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__b0_diff_2=0.0
*
* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 003, W = 3.01, L = 0.15
* ------------------------------------------------
+  sky130_fd_pr__rf_pfet_01v8_bM04__b1_diff_3=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__ub_diff_3=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__rdsw_diff_3=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_3=-0.022453
+  sky130_fd_pr__rf_pfet_01v8_bM04__kt1_diff_3=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__nfactor_diff_3=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__voff_diff_3=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__ags_diff_3=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__a0_diff_3=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__b0_diff_3=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_3=-0.00092315
+  sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_3=0.053737
+  sky130_fd_pr__rf_pfet_01v8_bM04__ua_diff_3=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_3=-16685.0
*
* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 004, W = 3.01, L = 0.18
* ------------------------------------------------
+  sky130_fd_pr__rf_pfet_01v8_bM04__ags_diff_4=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__a0_diff_4=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__voff_diff_4=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__b0_diff_4=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_4=-0.00093397
+  sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_4=0.059286
+  sky130_fd_pr__rf_pfet_01v8_bM04__ua_diff_4=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_4=-15584.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__b1_diff_4=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__ub_diff_4=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__rdsw_diff_4=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_4=-0.014614
+  sky130_fd_pr__rf_pfet_01v8_bM04__kt1_diff_4=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__nfactor_diff_4=0.0
*
* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 005, W = 3.01, L = 0.25
* ------------------------------------------------
+  sky130_fd_pr__rf_pfet_01v8_bM04__ags_diff_5=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__a0_diff_5=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__voff_diff_5=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__b0_diff_5=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_5=0.029916
+  sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_5=-0.00065774
+  sky130_fd_pr__rf_pfet_01v8_bM04__ua_diff_5=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_5=-21301.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__b1_diff_5=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__ub_diff_5=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__rdsw_diff_5=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_5=-0.0167
+  sky130_fd_pr__rf_pfet_01v8_bM04__kt1_diff_5=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__nfactor_diff_5=0.0
*
* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 006, W = 5.05, L = 0.15
* ------------------------------------------------
+  sky130_fd_pr__rf_pfet_01v8_bM04__kt1_diff_6=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__nfactor_diff_6=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__ags_diff_6=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__a0_diff_6=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__voff_diff_6=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__b0_diff_6=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_6=0.078414
+  sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_6=-0.0011357
+  sky130_fd_pr__rf_pfet_01v8_bM04__ua_diff_6=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_6=-13899.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__b1_diff_6=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__ub_diff_6=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__rdsw_diff_6=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_6=-0.024399
*
* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 007, W = 5.05, L = 0.18
* ------------------------------------------------
+  sky130_fd_pr__rf_pfet_01v8_bM04__rdsw_diff_7=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_7=-0.010627
+  sky130_fd_pr__rf_pfet_01v8_bM04__kt1_diff_7=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__nfactor_diff_7=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__ags_diff_7=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__a0_diff_7=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__voff_diff_7=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__b0_diff_7=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_7=0.049986
+  sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_7=-0.00088539
+  sky130_fd_pr__rf_pfet_01v8_bM04__ua_diff_7=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_7=-18591.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__b1_diff_7=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__ub_diff_7=0.0
*
* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 008, W = 5.05, L = 0.25
* ------------------------------------------------
+  sky130_fd_pr__rf_pfet_01v8_bM04__rdsw_diff_8=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_8=-0.012274
+  sky130_fd_pr__rf_pfet_01v8_bM04__kt1_diff_8=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__nfactor_diff_8=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__ags_diff_8=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__a0_diff_8=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__voff_diff_8=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__b0_diff_8=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_8=0.038873
+  sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_8=-0.000789
+  sky130_fd_pr__rf_pfet_01v8_bM04__ua_diff_8=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_8=-17257.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__b1_diff_8=0.0
+  sky130_fd_pr__rf_pfet_01v8_bM04__ub_diff_8=0.0
.include "sky130_fd_pr__rf_pfet_01v8_b.pm3.spice"
