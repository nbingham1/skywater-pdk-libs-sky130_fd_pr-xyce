* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 2
.param
+  sky130_fd_pr__rf_nfet_g5v0d10v5_b__toxe_mult=1.042
+  sky130_fd_pr__rf_nfet_g5v0d10v5_b__rbpb_mult=1.2
+  sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult=0.99758
+  sky130_fd_pr__rf_nfet_g5v0d10v5_b__ajunction_mult=1.1193
+  sky130_fd_pr__rf_nfet_g5v0d10v5_b__pjunction_mult=1.1801
+  sky130_fd_pr__rf_nfet_g5v0d10v5_b__lint_diff=-1.21275e-8
+  sky130_fd_pr__rf_nfet_g5v0d10v5_b__wint_diff=2.252e-8
+  sky130_fd_pr__rf_nfet_g5v0d10v5_b__rshg_diff=7.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_b__dlc_diff=-1.21275e-8
+  sky130_fd_pr__rf_nfet_g5v0d10v5_b__dwc_diff=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_b__xgw_diff=4.504e-8
*
* sky130_fd_pr__rf_nfet_g5v0d10v5_bM02, Bin 000, W = 3.01, L = 0.5
* --------------------------------------------
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__voff_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__ub_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__vth0_diff_0=0.037892
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__nfactor_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__ua_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__vsat_diff_0=-7490.2
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__a0_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__rdsw_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__b0_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__ags_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__k2_diff_0=0.0061192
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__kt1_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__pclm_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__u0_diff_0=-0.0068374
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__b1_diff_0=0.0
*
* sky130_fd_pr__rf_nfet_g5v0d10v5_bM02, Bin 001, W = 5.05, L = 0.5
* --------------------------------------------
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__voff_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__ub_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__vth0_diff_1=0.042869
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__nfactor_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__ua_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__vsat_diff_1=-5260.5
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__a0_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__rdsw_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__b0_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__ags_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__k2_diff_1=0.0082977
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__kt1_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__pclm_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__u0_diff_1=-0.0034898
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02__b1_diff_1=0.0
*
* sky130_fd_pr__rf_nfet_g5v0d10v5_bM04, Bin 000, W = 3.01, L = 0.5
* --------------------------------------------
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__nfactor_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__vsat_diff_0=-7602.3
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__vth0_diff_0=0.028278
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__a0_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__b0_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__k2_diff_0=0.0058947
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__u0_diff_0=-0.0070921
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__b1_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__ags_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__kt1_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__voff_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__pclm_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__ub_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__ua_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__rdsw_diff_0=0.0
*
* sky130_fd_pr__rf_nfet_g5v0d10v5_bM04, Bin 001, W = 5.05, L = 0.5
* --------------------------------------------
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__nfactor_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__vsat_diff_1=-7404.4
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__vth0_diff_1=0.035525
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__a0_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__b0_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__k2_diff_1=0.0078725
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__u0_diff_1=-0.0038822
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__b1_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__ags_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__kt1_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__voff_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__pclm_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__ub_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__ua_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__rdsw_diff_1=0.0
*
* sky130_fd_pr__rf_nfet_g5v0d10v5_bM04, Bin 002, W = 7.09, L = 0.5
* --------------------------------------------
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__rdsw_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__nfactor_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__vsat_diff_2=-8487.7
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__vth0_diff_2=0.039934
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__a0_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__b0_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__k2_diff_2=0.0052827
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__u0_diff_2=-0.0061567
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__b1_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__ags_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__kt1_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__voff_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__pclm_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__ub_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04__ua_diff_2=0.0
*
* sky130_fd_pr__rf_nfet_g5v0d10v5_bM10, Bin 000, W = 3.01, L = 0.5
* ---------------------------------------------
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__ags_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__ua_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__rdsw_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__k2_diff_0=0.0053572
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__kt1_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__pclm_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__u0_diff_0=-0.0056999
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__b1_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__voff_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__nfactor_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__ub_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__vth0_diff_0=0.037862
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__vsat_diff_0=86.018
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__a0_diff_0=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__b0_diff_0=0.0
*
* sky130_fd_pr__rf_nfet_g5v0d10v5_bM10, Bin 001, W = 5.05, L = 0.5
* ---------------------------------------------
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__b0_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__ags_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__ua_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__rdsw_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__k2_diff_1=0.001022
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__kt1_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__pclm_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__u0_diff_1=-0.0060669
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__b1_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__voff_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__nfactor_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__ub_diff_1=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__vth0_diff_1=0.032656
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__vsat_diff_1=-8977.1
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__a0_diff_1=0.0
*
* sky130_fd_pr__rf_nfet_g5v0d10v5_bM10, Bin 002, W = 7.09, L = 0.5
* ---------------------------------------------
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__a0_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__b0_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__ua_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__ags_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__rdsw_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__k2_diff_2=0.0043107
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__kt1_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__pclm_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__u0_diff_2=-0.011734
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__b1_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__voff_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__nfactor_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__ub_diff_2=0.0
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__vth0_diff_2=0.025004
+  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10__vsat_diff_2=-884.49
.include "sky130_fd_pr__rf_nfet_g5v0d10v5_b.pm3.spice"
