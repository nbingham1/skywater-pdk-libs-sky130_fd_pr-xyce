* SKY130 Spice File.
.param globalk=1
.param localkswitch=1
.param capunits='1.0*1e-6'
.param
+  mcp1f_ca_w_0_150_s_0_210=8.67e-05 mcp1f_cc_w_0_150_s_0_210=6.82e-11 mcp1f_cf_w_0_150_s_0_210=9.08e-12
+  mcp1f_ca_w_0_150_s_0_263=8.67e-05 mcp1f_cc_w_0_150_s_0_263=5.67e-11 mcp1f_cf_w_0_150_s_0_263=1.09e-11
+  mcp1f_ca_w_0_150_s_0_315=8.67e-05 mcp1f_cc_w_0_150_s_0_315=4.92e-11 mcp1f_cf_w_0_150_s_0_315=1.26e-11
+  mcp1f_ca_w_0_150_s_0_420=8.67e-05 mcp1f_cc_w_0_150_s_0_420=3.84e-11 mcp1f_cf_w_0_150_s_0_420=1.60e-11
+  mcp1f_ca_w_0_150_s_0_525=8.67e-05 mcp1f_cc_w_0_150_s_0_525=3.18e-11 mcp1f_cf_w_0_150_s_0_525=1.89e-11
+  mcp1f_ca_w_0_150_s_0_630=8.67e-05 mcp1f_cc_w_0_150_s_0_630=2.70e-11 mcp1f_cf_w_0_150_s_0_630=2.14e-11
+  mcp1f_ca_w_0_150_s_0_840=8.67e-05 mcp1f_cc_w_0_150_s_0_840=2.01e-11 mcp1f_cf_w_0_150_s_0_840=2.57e-11
+  mcp1f_ca_w_0_150_s_1_260=8.67e-05 mcp1f_cc_w_0_150_s_1_260=1.20e-11 mcp1f_cf_w_0_150_s_1_260=3.22e-11
+  mcp1f_ca_w_0_150_s_2_310=8.67e-05 mcp1f_cc_w_0_150_s_2_310=5.31e-12 mcp1f_cf_w_0_150_s_2_310=3.82e-11
+  mcp1f_ca_w_0_150_s_5_250=8.67e-05 mcp1f_cc_w_0_150_s_5_250=1.24e-12 mcp1f_cf_w_0_150_s_5_250=4.23e-11
+  mcp1f_ca_w_1_200_s_0_210=8.67e-05 mcp1f_cc_w_1_200_s_0_210=8.65e-11 mcp1f_cf_w_1_200_s_0_210=9.01e-12
+  mcp1f_ca_w_1_200_s_0_263=8.67e-05 mcp1f_cc_w_1_200_s_0_263=7.39e-11 mcp1f_cf_w_1_200_s_0_263=1.09e-11
+  mcp1f_ca_w_1_200_s_0_315=8.67e-05 mcp1f_cc_w_1_200_s_0_315=6.50e-11 mcp1f_cf_w_1_200_s_0_315=1.27e-11
+  mcp1f_ca_w_1_200_s_0_420=8.67e-05 mcp1f_cc_w_1_200_s_0_420=5.30e-11 mcp1f_cf_w_1_200_s_0_420=1.60e-11
+  mcp1f_ca_w_1_200_s_0_525=8.67e-05 mcp1f_cc_w_1_200_s_0_525=4.49e-11 mcp1f_cf_w_1_200_s_0_525=1.90e-11
+  mcp1f_ca_w_1_200_s_0_630=8.67e-05 mcp1f_cc_w_1_200_s_0_630=3.92e-11 mcp1f_cf_w_1_200_s_0_630=2.17e-11
+  mcp1f_ca_w_1_200_s_0_840=8.67e-05 mcp1f_cc_w_1_200_s_0_840=3.10e-11 mcp1f_cf_w_1_200_s_0_840=2.63e-11
+  mcp1f_ca_w_1_200_s_1_260=8.67e-05 mcp1f_cc_w_1_200_s_1_260=2.15e-11 mcp1f_cf_w_1_200_s_1_260=3.31e-11
+  mcp1f_ca_w_1_200_s_2_310=8.67e-05 mcp1f_cc_w_1_200_s_2_310=1.10e-11 mcp1f_cf_w_1_200_s_2_310=4.22e-11
+  mcp1f_ca_w_1_200_s_5_250=8.67e-05 mcp1f_cc_w_1_200_s_5_250=3.55e-12 mcp1f_cf_w_1_200_s_5_250=4.94e-11
+  mcl1f_ca_w_0_170_s_0_180=3.12e-05 mcl1f_cc_w_0_170_s_0_180=6.92e-11 mcl1f_cf_w_0_170_s_0_180=3.11e-12
+  mcl1f_ca_w_0_170_s_0_225=3.12e-05 mcl1f_cc_w_0_170_s_0_225=6.05e-11 mcl1f_cf_w_0_170_s_0_225=3.78e-12
+  mcl1f_ca_w_0_170_s_0_270=3.12e-05 mcl1f_cc_w_0_170_s_0_270=5.48e-11 mcl1f_cf_w_0_170_s_0_270=4.43e-12
+  mcl1f_ca_w_0_170_s_0_360=3.12e-05 mcl1f_cc_w_0_170_s_0_360=4.57e-11 mcl1f_cf_w_0_170_s_0_360=5.88e-12
+  mcl1f_ca_w_0_170_s_0_450=3.12e-05 mcl1f_cc_w_0_170_s_0_450=4.02e-11 mcl1f_cf_w_0_170_s_0_450=6.93e-12
+  mcl1f_ca_w_0_170_s_0_540=3.12e-05 mcl1f_cc_w_0_170_s_0_540=3.54e-11 mcl1f_cf_w_0_170_s_0_540=8.34e-12
+  mcl1f_ca_w_0_170_s_0_720=3.12e-05 mcl1f_cc_w_0_170_s_0_720=2.90e-11 mcl1f_cf_w_0_170_s_0_720=1.06e-11
+  mcl1f_ca_w_0_170_s_1_080=3.12e-05 mcl1f_cc_w_0_170_s_1_080=2.11e-11 mcl1f_cf_w_0_170_s_1_080=1.45e-11
+  mcl1f_ca_w_0_170_s_1_980=3.12e-05 mcl1f_cc_w_0_170_s_1_980=1.19e-11 mcl1f_cf_w_0_170_s_1_980=2.09e-11
+  mcl1f_ca_w_0_170_s_4_500=3.12e-05 mcl1f_cc_w_0_170_s_4_500=3.77e-12 mcl1f_cf_w_0_170_s_4_500=2.82e-11
+  mcl1f_ca_w_1_360_s_0_180=3.12e-05 mcl1f_cc_w_1_360_s_0_180=9.22e-11 mcl1f_cf_w_1_360_s_0_180=3.11e-12
+  mcl1f_ca_w_1_360_s_0_225=3.12e-05 mcl1f_cc_w_1_360_s_0_225=8.24e-11 mcl1f_cf_w_1_360_s_0_225=3.78e-12
+  mcl1f_ca_w_1_360_s_0_270=3.12e-05 mcl1f_cc_w_1_360_s_0_270=7.49e-11 mcl1f_cf_w_1_360_s_0_270=4.44e-12
+  mcl1f_ca_w_1_360_s_0_360=3.12e-05 mcl1f_cc_w_1_360_s_0_360=6.41e-11 mcl1f_cf_w_1_360_s_0_360=5.74e-12
+  mcl1f_ca_w_1_360_s_0_450=3.12e-05 mcl1f_cc_w_1_360_s_0_450=5.67e-11 mcl1f_cf_w_1_360_s_0_450=7.00e-12
+  mcl1f_ca_w_1_360_s_0_540=3.12e-05 mcl1f_cc_w_1_360_s_0_540=5.10e-11 mcl1f_cf_w_1_360_s_0_540=8.21e-12
+  mcl1f_ca_w_1_360_s_0_720=3.12e-05 mcl1f_cc_w_1_360_s_0_720=4.29e-11 mcl1f_cf_w_1_360_s_0_720=1.05e-11
+  mcl1f_ca_w_1_360_s_1_080=3.12e-05 mcl1f_cc_w_1_360_s_1_080=3.28e-11 mcl1f_cf_w_1_360_s_1_080=1.47e-11
+  mcl1f_ca_w_1_360_s_1_980=3.12e-05 mcl1f_cc_w_1_360_s_1_980=1.99e-11 mcl1f_cf_w_1_360_s_1_980=2.26e-11
+  mcl1f_ca_w_1_360_s_4_500=3.12e-05 mcl1f_cc_w_1_360_s_4_500=7.70e-12 mcl1f_cf_w_1_360_s_4_500=3.30e-11
+  mcl1d_ca_w_0_170_s_0_180=4.77e-05 mcl1d_cc_w_0_170_s_0_180=6.69e-11 mcl1d_cf_w_0_170_s_0_180=4.71e-12
+  mcl1d_ca_w_0_170_s_0_225=4.77e-05 mcl1d_cc_w_0_170_s_0_225=5.81e-11 mcl1d_cf_w_0_170_s_0_225=5.71e-12
+  mcl1d_ca_w_0_170_s_0_270=4.77e-05 mcl1d_cc_w_0_170_s_0_270=5.21e-11 mcl1d_cf_w_0_170_s_0_270=6.65e-12
+  mcl1d_ca_w_0_170_s_0_360=4.77e-05 mcl1d_cc_w_0_170_s_0_360=4.28e-11 mcl1d_cf_w_0_170_s_0_360=8.74e-12
+  mcl1d_ca_w_0_170_s_0_450=4.77e-05 mcl1d_cc_w_0_170_s_0_450=3.71e-11 mcl1d_cf_w_0_170_s_0_450=1.03e-11
+  mcl1d_ca_w_0_170_s_0_540=4.77e-05 mcl1d_cc_w_0_170_s_0_540=3.21e-11 mcl1d_cf_w_0_170_s_0_540=1.22e-11
+  mcl1d_ca_w_0_170_s_0_720=4.77e-05 mcl1d_cc_w_0_170_s_0_720=2.54e-11 mcl1d_cf_w_0_170_s_0_720=1.53e-11
+  mcl1d_ca_w_0_170_s_1_080=4.77e-05 mcl1d_cc_w_0_170_s_1_080=1.74e-11 mcl1d_cf_w_0_170_s_1_080=2.03e-11
+  mcl1d_ca_w_0_170_s_1_980=4.77e-05 mcl1d_cc_w_0_170_s_1_980=8.68e-12 mcl1d_cf_w_0_170_s_1_980=2.72e-11
+  mcl1d_ca_w_0_170_s_4_500=4.77e-05 mcl1d_cc_w_0_170_s_4_500=2.43e-12 mcl1d_cf_w_0_170_s_4_500=3.32e-11
+  mcl1d_ca_w_1_360_s_0_180=4.77e-05 mcl1d_cc_w_1_360_s_0_180=8.77e-11 mcl1d_cf_w_1_360_s_0_180=4.71e-12
+  mcl1d_ca_w_1_360_s_0_225=4.77e-05 mcl1d_cc_w_1_360_s_0_225=7.78e-11 mcl1d_cf_w_1_360_s_0_225=5.70e-12
+  mcl1d_ca_w_1_360_s_0_270=4.77e-05 mcl1d_cc_w_1_360_s_0_270=7.03e-11 mcl1d_cf_w_1_360_s_0_270=6.68e-12
+  mcl1d_ca_w_1_360_s_0_360=4.77e-05 mcl1d_cc_w_1_360_s_0_360=5.95e-11 mcl1d_cf_w_1_360_s_0_360=8.57e-12
+  mcl1d_ca_w_1_360_s_0_450=4.77e-05 mcl1d_cc_w_1_360_s_0_450=5.21e-11 mcl1d_cf_w_1_360_s_0_450=1.04e-11
+  mcl1d_ca_w_1_360_s_0_540=4.77e-05 mcl1d_cc_w_1_360_s_0_540=4.65e-11 mcl1d_cf_w_1_360_s_0_540=1.21e-11
+  mcl1d_ca_w_1_360_s_0_720=4.77e-05 mcl1d_cc_w_1_360_s_0_720=3.83e-11 mcl1d_cf_w_1_360_s_0_720=1.53e-11
+  mcl1d_ca_w_1_360_s_1_080=4.77e-05 mcl1d_cc_w_1_360_s_1_080=2.83e-11 mcl1d_cf_w_1_360_s_1_080=2.07e-11
+  mcl1d_ca_w_1_360_s_1_980=4.77e-05 mcl1d_cc_w_1_360_s_1_980=1.60e-11 mcl1d_cf_w_1_360_s_1_980=2.97e-11
+  mcl1d_ca_w_1_360_s_4_500=4.77e-05 mcl1d_cc_w_1_360_s_4_500=5.70e-12 mcl1d_cf_w_1_360_s_4_500=3.92e-11
+  mcl1p1_ca_w_0_170_s_0_180=7.09e-05 mcl1p1_cc_w_0_170_s_0_180=6.41e-11 mcl1p1_cf_w_0_170_s_0_180=6.89e-12
+  mcl1p1_ca_w_0_170_s_0_225=7.09e-05 mcl1p1_cc_w_0_170_s_0_225=5.51e-11 mcl1p1_cf_w_0_170_s_0_225=8.32e-12
+  mcl1p1_ca_w_0_170_s_0_270=7.09e-05 mcl1p1_cc_w_0_170_s_0_270=4.90e-11 mcl1p1_cf_w_0_170_s_0_270=9.65e-12
+  mcl1p1_ca_w_0_170_s_0_360=7.09e-05 mcl1p1_cc_w_0_170_s_0_360=3.94e-11 mcl1p1_cf_w_0_170_s_0_360=1.25e-11
+  mcl1p1_ca_w_0_170_s_0_450=7.09e-05 mcl1p1_cc_w_0_170_s_0_450=3.36e-11 mcl1p1_cf_w_0_170_s_0_450=1.46e-11
+  mcl1p1_ca_w_0_170_s_0_540=7.09e-05 mcl1p1_cc_w_0_170_s_0_540=2.84e-11 mcl1p1_cf_w_0_170_s_0_540=1.72e-11
+  mcl1p1_ca_w_0_170_s_0_720=7.09e-05 mcl1p1_cc_w_0_170_s_0_720=2.17e-11 mcl1p1_cf_w_0_170_s_0_720=2.11e-11
+  mcl1p1_ca_w_0_170_s_1_080=7.09e-05 mcl1p1_cc_w_0_170_s_1_080=1.38e-11 mcl1p1_cf_w_0_170_s_1_080=2.68e-11
+  mcl1p1_ca_w_0_170_s_1_980=7.09e-05 mcl1p1_cc_w_0_170_s_1_980=6.23e-12 mcl1p1_cf_w_0_170_s_1_980=3.35e-11
+  mcl1p1_ca_w_0_170_s_4_500=7.09e-05 mcl1p1_cc_w_0_170_s_4_500=1.61e-12 mcl1p1_cf_w_0_170_s_4_500=3.80e-11
+  mcl1p1_ca_w_1_360_s_0_180=7.09e-05 mcl1p1_cc_w_1_360_s_0_180=8.32e-11 mcl1p1_cf_w_1_360_s_0_180=6.92e-12
+  mcl1p1_ca_w_1_360_s_0_225=7.09e-05 mcl1p1_cc_w_1_360_s_0_225=7.34e-11 mcl1p1_cf_w_1_360_s_0_225=8.35e-12
+  mcl1p1_ca_w_1_360_s_0_270=7.09e-05 mcl1p1_cc_w_1_360_s_0_270=6.59e-11 mcl1p1_cf_w_1_360_s_0_270=9.73e-12
+  mcl1p1_ca_w_1_360_s_0_360=7.09e-05 mcl1p1_cc_w_1_360_s_0_360=5.51e-11 mcl1p1_cf_w_1_360_s_0_360=1.24e-11
+  mcl1p1_ca_w_1_360_s_0_450=7.09e-05 mcl1p1_cc_w_1_360_s_0_450=4.78e-11 mcl1p1_cf_w_1_360_s_0_450=1.48e-11
+  mcl1p1_ca_w_1_360_s_0_540=7.09e-05 mcl1p1_cc_w_1_360_s_0_540=4.22e-11 mcl1p1_cf_w_1_360_s_0_540=1.71e-11
+  mcl1p1_ca_w_1_360_s_0_720=7.09e-05 mcl1p1_cc_w_1_360_s_0_720=3.41e-11 mcl1p1_cf_w_1_360_s_0_720=2.12e-11
+  mcl1p1_ca_w_1_360_s_1_080=7.09e-05 mcl1p1_cc_w_1_360_s_1_080=2.44e-11 mcl1p1_cf_w_1_360_s_1_080=2.76e-11
+  mcl1p1_ca_w_1_360_s_1_980=7.09e-05 mcl1p1_cc_w_1_360_s_1_980=1.30e-11 mcl1p1_cf_w_1_360_s_1_980=3.70e-11
+  mcl1p1_ca_w_1_360_s_4_500=7.09e-05 mcl1p1_cc_w_1_360_s_4_500=4.40e-12 mcl1p1_cf_w_1_360_s_4_500=4.53e-11
+  mcm1f_ca_w_0_140_s_0_140=2.17e-05 mcm1f_cc_w_0_140_s_0_140=9.19e-11 mcm1f_cf_w_0_140_s_0_140=1.73e-12
+  mcm1f_ca_w_0_140_s_0_175=2.17e-05 mcm1f_cc_w_0_140_s_0_175=9.15e-11 mcm1f_cf_w_0_140_s_0_175=2.11e-12
+  mcm1f_ca_w_0_140_s_0_210=2.17e-05 mcm1f_cc_w_0_140_s_0_210=8.72e-11 mcm1f_cf_w_0_140_s_0_210=2.49e-12
+  mcm1f_ca_w_0_140_s_0_280=2.17e-05 mcm1f_cc_w_0_140_s_0_280=7.94e-11 mcm1f_cf_w_0_140_s_0_280=3.23e-12
+  mcm1f_ca_w_0_140_s_0_350=2.17e-05 mcm1f_cc_w_0_140_s_0_350=7.00e-11 mcm1f_cf_w_0_140_s_0_350=3.95e-12
+  mcm1f_ca_w_0_140_s_0_420=2.17e-05 mcm1f_cc_w_0_140_s_0_420=6.21e-11 mcm1f_cf_w_0_140_s_0_420=4.72e-12
+  mcm1f_ca_w_0_140_s_0_560=2.17e-05 mcm1f_cc_w_0_140_s_0_560=5.17e-11 mcm1f_cf_w_0_140_s_0_560=6.07e-12
+  mcm1f_ca_w_0_140_s_0_840=2.17e-05 mcm1f_cc_w_0_140_s_0_840=3.93e-11 mcm1f_cf_w_0_140_s_0_840=8.70e-12
+  mcm1f_ca_w_0_140_s_1_540=2.17e-05 mcm1f_cc_w_0_140_s_1_540=2.48e-11 mcm1f_cf_w_0_140_s_1_540=1.44e-11
+  mcm1f_ca_w_0_140_s_3_500=2.17e-05 mcm1f_cc_w_0_140_s_3_500=1.07e-11 mcm1f_cf_w_0_140_s_3_500=2.41e-11
+  mcm1f_ca_w_1_120_s_0_140=2.17e-05 mcm1f_cc_w_1_120_s_0_140=1.19e-10 mcm1f_cf_w_1_120_s_0_140=1.76e-12
+  mcm1f_ca_w_1_120_s_0_175=2.17e-05 mcm1f_cc_w_1_120_s_0_175=1.16e-10 mcm1f_cf_w_1_120_s_0_175=2.14e-12
+  mcm1f_ca_w_1_120_s_0_210=2.17e-05 mcm1f_cc_w_1_120_s_0_210=1.11e-10 mcm1f_cf_w_1_120_s_0_210=2.51e-12
+  mcm1f_ca_w_1_120_s_0_280=2.17e-05 mcm1f_cc_w_1_120_s_0_280=1.00e-10 mcm1f_cf_w_1_120_s_0_280=3.26e-12
+  mcm1f_ca_w_1_120_s_0_350=2.17e-05 mcm1f_cc_w_1_120_s_0_350=8.94e-11 mcm1f_cf_w_1_120_s_0_350=4.00e-12
+  mcm1f_ca_w_1_120_s_0_420=2.17e-05 mcm1f_cc_w_1_120_s_0_420=8.02e-11 mcm1f_cf_w_1_120_s_0_420=4.72e-12
+  mcm1f_ca_w_1_120_s_0_560=2.17e-05 mcm1f_cc_w_1_120_s_0_560=6.69e-11 mcm1f_cf_w_1_120_s_0_560=6.12e-12
+  mcm1f_ca_w_1_120_s_0_840=2.17e-05 mcm1f_cc_w_1_120_s_0_840=5.15e-11 mcm1f_cf_w_1_120_s_0_840=8.79e-12
+  mcm1f_ca_w_1_120_s_1_540=2.17e-05 mcm1f_cc_w_1_120_s_1_540=3.35e-11 mcm1f_cf_w_1_120_s_1_540=1.47e-11
+  mcm1f_ca_w_1_120_s_3_500=2.17e-05 mcm1f_cc_w_1_120_s_3_500=1.57e-11 mcm1f_cf_w_1_120_s_3_500=2.57e-11
+  mcm1d_ca_w_0_140_s_0_140=2.86e-05 mcm1d_cc_w_0_140_s_0_140=9.11e-11 mcm1d_cf_w_0_140_s_0_140=2.27e-12
+  mcm1d_ca_w_0_140_s_0_175=2.86e-05 mcm1d_cc_w_0_140_s_0_175=9.07e-11 mcm1d_cf_w_0_140_s_0_175=2.77e-12
+  mcm1d_ca_w_0_140_s_0_210=2.86e-05 mcm1d_cc_w_0_140_s_0_210=8.67e-11 mcm1d_cf_w_0_140_s_0_210=3.27e-12
+  mcm1d_ca_w_0_140_s_0_280=2.86e-05 mcm1d_cc_w_0_140_s_0_280=7.80e-11 mcm1d_cf_w_0_140_s_0_280=4.24e-12
+  mcm1d_ca_w_0_140_s_0_350=2.86e-05 mcm1d_cc_w_0_140_s_0_350=6.88e-11 mcm1d_cf_w_0_140_s_0_350=5.17e-12
+  mcm1d_ca_w_0_140_s_0_420=2.86e-05 mcm1d_cc_w_0_140_s_0_420=6.09e-11 mcm1d_cf_w_0_140_s_0_420=6.16e-12
+  mcm1d_ca_w_0_140_s_0_560=2.86e-05 mcm1d_cc_w_0_140_s_0_560=4.99e-11 mcm1d_cf_w_0_140_s_0_560=7.90e-12
+  mcm1d_ca_w_0_140_s_0_840=2.86e-05 mcm1d_cc_w_0_140_s_0_840=3.73e-11 mcm1d_cf_w_0_140_s_0_840=1.12e-11
+  mcm1d_ca_w_0_140_s_1_540=2.86e-05 mcm1d_cc_w_0_140_s_1_540=2.24e-11 mcm1d_cf_w_0_140_s_1_540=1.81e-11
+  mcm1d_ca_w_0_140_s_3_500=2.86e-05 mcm1d_cc_w_0_140_s_3_500=8.78e-12 mcm1d_cf_w_0_140_s_3_500=2.84e-11
+  mcm1d_ca_w_1_120_s_0_140=2.86e-05 mcm1d_cc_w_1_120_s_0_140=1.16e-10 mcm1d_cf_w_1_120_s_0_140=2.32e-12
+  mcm1d_ca_w_1_120_s_0_175=2.86e-05 mcm1d_cc_w_1_120_s_0_175=1.13e-10 mcm1d_cf_w_1_120_s_0_175=2.82e-12
+  mcm1d_ca_w_1_120_s_0_210=2.86e-05 mcm1d_cc_w_1_120_s_0_210=1.09e-10 mcm1d_cf_w_1_120_s_0_210=3.31e-12
+  mcm1d_ca_w_1_120_s_0_280=2.86e-05 mcm1d_cc_w_1_120_s_0_280=9.74e-11 mcm1d_cf_w_1_120_s_0_280=4.29e-12
+  mcm1d_ca_w_1_120_s_0_350=2.86e-05 mcm1d_cc_w_1_120_s_0_350=8.66e-11 mcm1d_cf_w_1_120_s_0_350=5.25e-12
+  mcm1d_ca_w_1_120_s_0_420=2.86e-05 mcm1d_cc_w_1_120_s_0_420=7.74e-11 mcm1d_cf_w_1_120_s_0_420=6.18e-12
+  mcm1d_ca_w_1_120_s_0_560=2.86e-05 mcm1d_cc_w_1_120_s_0_560=6.42e-11 mcm1d_cf_w_1_120_s_0_560=7.98e-12
+  mcm1d_ca_w_1_120_s_0_840=2.86e-05 mcm1d_cc_w_1_120_s_0_840=4.85e-11 mcm1d_cf_w_1_120_s_0_840=1.14e-11
+  mcm1d_ca_w_1_120_s_1_540=2.86e-05 mcm1d_cc_w_1_120_s_1_540=3.06e-11 mcm1d_cf_w_1_120_s_1_540=1.85e-11
+  mcm1d_ca_w_1_120_s_3_500=2.86e-05 mcm1d_cc_w_1_120_s_3_500=1.34e-11 mcm1d_cf_w_1_120_s_3_500=3.06e-11
+  mcm1p1_ca_w_0_140_s_0_140=3.55e-05 mcm1p1_cc_w_0_140_s_0_140=9.03e-11 mcm1p1_cf_w_0_140_s_0_140=2.82e-12
+  mcm1p1_ca_w_0_140_s_0_175=3.55e-05 mcm1p1_cc_w_0_140_s_0_175=8.93e-11 mcm1p1_cf_w_0_140_s_0_175=3.44e-12
+  mcm1p1_ca_w_0_140_s_0_210=3.55e-05 mcm1p1_cc_w_0_140_s_0_210=8.60e-11 mcm1p1_cf_w_0_140_s_0_210=4.05e-12
+  mcm1p1_ca_w_0_140_s_0_280=3.55e-05 mcm1p1_cc_w_0_140_s_0_280=7.65e-11 mcm1p1_cf_w_0_140_s_0_280=5.25e-12
+  mcm1p1_ca_w_0_140_s_0_350=3.55e-05 mcm1p1_cc_w_0_140_s_0_350=6.73e-11 mcm1p1_cf_w_0_140_s_0_350=6.41e-12
+  mcm1p1_ca_w_0_140_s_0_420=3.55e-05 mcm1p1_cc_w_0_140_s_0_420=5.96e-11 mcm1p1_cf_w_0_140_s_0_420=7.61e-12
+  mcm1p1_ca_w_0_140_s_0_560=3.55e-05 mcm1p1_cc_w_0_140_s_0_560=4.83e-11 mcm1p1_cf_w_0_140_s_0_560=9.73e-12
+  mcm1p1_ca_w_0_140_s_0_840=3.55e-05 mcm1p1_cc_w_0_140_s_0_840=3.54e-11 mcm1p1_cf_w_0_140_s_0_840=1.37e-11
+  mcm1p1_ca_w_0_140_s_1_540=3.55e-05 mcm1p1_cc_w_0_140_s_1_540=2.04e-11 mcm1p1_cf_w_0_140_s_1_540=2.15e-11
+  mcm1p1_ca_w_0_140_s_3_500=3.55e-05 mcm1p1_cc_w_0_140_s_3_500=7.39e-12 mcm1p1_cf_w_0_140_s_3_500=3.21e-11
+  mcm1p1_ca_w_1_120_s_0_140=3.55e-05 mcm1p1_cc_w_1_120_s_0_140=1.14e-10 mcm1p1_cf_w_1_120_s_0_140=2.91e-12
+  mcm1p1_ca_w_1_120_s_0_175=3.55e-05 mcm1p1_cc_w_1_120_s_0_175=1.11e-10 mcm1p1_cf_w_1_120_s_0_175=3.53e-12
+  mcm1p1_ca_w_1_120_s_0_210=3.55e-05 mcm1p1_cc_w_1_120_s_0_210=1.06e-10 mcm1p1_cf_w_1_120_s_0_210=4.13e-12
+  mcm1p1_ca_w_1_120_s_0_280=3.55e-05 mcm1p1_cc_w_1_120_s_0_280=9.50e-11 mcm1p1_cf_w_1_120_s_0_280=5.34e-12
+  mcm1p1_ca_w_1_120_s_0_350=3.55e-05 mcm1p1_cc_w_1_120_s_0_350=8.43e-11 mcm1p1_cf_w_1_120_s_0_350=6.52e-12
+  mcm1p1_ca_w_1_120_s_0_420=3.55e-05 mcm1p1_cc_w_1_120_s_0_420=7.52e-11 mcm1p1_cf_w_1_120_s_0_420=7.66e-12
+  mcm1p1_ca_w_1_120_s_0_560=3.55e-05 mcm1p1_cc_w_1_120_s_0_560=6.17e-11 mcm1p1_cf_w_1_120_s_0_560=9.84e-12
+  mcm1p1_ca_w_1_120_s_0_840=3.55e-05 mcm1p1_cc_w_1_120_s_0_840=4.62e-11 mcm1p1_cf_w_1_120_s_0_840=1.39e-11
+  mcm1p1_ca_w_1_120_s_1_540=3.55e-05 mcm1p1_cc_w_1_120_s_1_540=2.83e-11 mcm1p1_cf_w_1_120_s_1_540=2.21e-11
+  mcm1p1_ca_w_1_120_s_3_500=3.55e-05 mcm1p1_cc_w_1_120_s_3_500=1.18e-11 mcm1p1_cf_w_1_120_s_3_500=3.46e-11
+  mcm1l1_ca_w_0_140_s_0_140=8.73e-05 mcm1l1_cc_w_0_140_s_0_140=8.54e-11 mcm1l1_cf_w_0_140_s_0_140=6.63e-12
+  mcm1l1_ca_w_0_140_s_0_175=8.73e-05 mcm1l1_cc_w_0_140_s_0_175=8.41e-11 mcm1l1_cf_w_0_140_s_0_175=8.14e-12
+  mcm1l1_ca_w_0_140_s_0_210=8.73e-05 mcm1l1_cc_w_0_140_s_0_210=7.97e-11 mcm1l1_cf_w_0_140_s_0_210=9.58e-12
+  mcm1l1_ca_w_0_140_s_0_280=8.73e-05 mcm1l1_cc_w_0_140_s_0_280=7.00e-11 mcm1l1_cf_w_0_140_s_0_280=1.24e-11
+  mcm1l1_ca_w_0_140_s_0_350=8.73e-05 mcm1l1_cc_w_0_140_s_0_350=6.04e-11 mcm1l1_cf_w_0_140_s_0_350=1.50e-11
+  mcm1l1_ca_w_0_140_s_0_420=8.73e-05 mcm1l1_cc_w_0_140_s_0_420=5.18e-11 mcm1l1_cf_w_0_140_s_0_420=1.75e-11
+  mcm1l1_ca_w_0_140_s_0_560=8.73e-05 mcm1l1_cc_w_0_140_s_0_560=4.01e-11 mcm1l1_cf_w_0_140_s_0_560=2.18e-11
+  mcm1l1_ca_w_0_140_s_0_840=8.73e-05 mcm1l1_cc_w_0_140_s_0_840=2.71e-11 mcm1l1_cf_w_0_140_s_0_840=2.89e-11
+  mcm1l1_ca_w_0_140_s_1_540=8.73e-05 mcm1l1_cc_w_0_140_s_1_540=1.30e-11 mcm1l1_cf_w_0_140_s_1_540=3.96e-11
+  mcm1l1_ca_w_0_140_s_3_500=8.73e-05 mcm1l1_cc_w_0_140_s_3_500=3.75e-12 mcm1l1_cf_w_0_140_s_3_500=4.85e-11
+  mcm1l1_ca_w_1_120_s_0_140=8.73e-05 mcm1l1_cc_w_1_120_s_0_140=1.04e-10 mcm1l1_cf_w_1_120_s_0_140=6.71e-12
+  mcm1l1_ca_w_1_120_s_0_175=8.73e-05 mcm1l1_cc_w_1_120_s_0_175=1.02e-10 mcm1l1_cf_w_1_120_s_0_175=8.23e-12
+  mcm1l1_ca_w_1_120_s_0_210=8.73e-05 mcm1l1_cc_w_1_120_s_0_210=9.63e-11 mcm1l1_cf_w_1_120_s_0_210=9.67e-12
+  mcm1l1_ca_w_1_120_s_0_280=8.73e-05 mcm1l1_cc_w_1_120_s_0_280=8.48e-11 mcm1l1_cf_w_1_120_s_0_280=1.24e-11
+  mcm1l1_ca_w_1_120_s_0_350=8.73e-05 mcm1l1_cc_w_1_120_s_0_350=7.40e-11 mcm1l1_cf_w_1_120_s_0_350=1.50e-11
+  mcm1l1_ca_w_1_120_s_0_420=8.73e-05 mcm1l1_cc_w_1_120_s_0_420=6.50e-11 mcm1l1_cf_w_1_120_s_0_420=1.75e-11
+  mcm1l1_ca_w_1_120_s_0_560=8.73e-05 mcm1l1_cc_w_1_120_s_0_560=5.17e-11 mcm1l1_cf_w_1_120_s_0_560=2.19e-11
+  mcm1l1_ca_w_1_120_s_0_840=8.73e-05 mcm1l1_cc_w_1_120_s_0_840=3.68e-11 mcm1l1_cf_w_1_120_s_0_840=2.91e-11
+  mcm1l1_ca_w_1_120_s_1_540=8.73e-05 mcm1l1_cc_w_1_120_s_1_540=2.04e-11 mcm1l1_cf_w_1_120_s_1_540=4.07e-11
+  mcm1l1_ca_w_1_120_s_3_500=8.73e-05 mcm1l1_cc_w_1_120_s_3_500=7.40e-12 mcm1l1_cf_w_1_120_s_3_500=5.25e-11
+  mcm2f_ca_w_0_140_s_0_140=1.49e-05 mcm2f_cc_w_0_140_s_0_140=9.27e-11 mcm2f_cf_w_0_140_s_0_140=1.20e-12
+  mcm2f_ca_w_0_140_s_0_175=1.49e-05 mcm2f_cc_w_0_140_s_0_175=9.17e-11 mcm2f_cf_w_0_140_s_0_175=1.46e-12
+  mcm2f_ca_w_0_140_s_0_210=1.49e-05 mcm2f_cc_w_0_140_s_0_210=8.82e-11 mcm2f_cf_w_0_140_s_0_210=1.72e-12
+  mcm2f_ca_w_0_140_s_0_280=1.49e-05 mcm2f_cc_w_0_140_s_0_280=8.06e-11 mcm2f_cf_w_0_140_s_0_280=2.24e-12
+  mcm2f_ca_w_0_140_s_0_350=1.49e-05 mcm2f_cc_w_0_140_s_0_350=7.12e-11 mcm2f_cf_w_0_140_s_0_350=2.74e-12
+  mcm2f_ca_w_0_140_s_0_420=1.49e-05 mcm2f_cc_w_0_140_s_0_420=6.34e-11 mcm2f_cf_w_0_140_s_0_420=3.28e-12
+  mcm2f_ca_w_0_140_s_0_560=1.49e-05 mcm2f_cc_w_0_140_s_0_560=5.30e-11 mcm2f_cf_w_0_140_s_0_560=4.23e-12
+  mcm2f_ca_w_0_140_s_0_840=1.49e-05 mcm2f_cc_w_0_140_s_0_840=4.13e-11 mcm2f_cf_w_0_140_s_0_840=6.12e-12
+  mcm2f_ca_w_0_140_s_1_540=1.49e-05 mcm2f_cc_w_0_140_s_1_540=2.73e-11 mcm2f_cf_w_0_140_s_1_540=1.04e-11
+  mcm2f_ca_w_0_140_s_3_500=1.49e-05 mcm2f_cc_w_0_140_s_3_500=1.33e-11 mcm2f_cf_w_0_140_s_3_500=1.87e-11
+  mcm2f_ca_w_1_120_s_0_140=1.49e-05 mcm2f_cc_w_1_120_s_0_140=1.21e-10 mcm2f_cf_w_1_120_s_0_140=1.22e-12
+  mcm2f_ca_w_1_120_s_0_175=1.49e-05 mcm2f_cc_w_1_120_s_0_175=1.18e-10 mcm2f_cf_w_1_120_s_0_175=1.48e-12
+  mcm2f_ca_w_1_120_s_0_210=1.49e-05 mcm2f_cc_w_1_120_s_0_210=1.14e-10 mcm2f_cf_w_1_120_s_0_210=1.74e-12
+  mcm2f_ca_w_1_120_s_0_280=1.49e-05 mcm2f_cc_w_1_120_s_0_280=1.03e-10 mcm2f_cf_w_1_120_s_0_280=2.26e-12
+  mcm2f_ca_w_1_120_s_0_350=1.49e-05 mcm2f_cc_w_1_120_s_0_350=9.18e-11 mcm2f_cf_w_1_120_s_0_350=2.77e-12
+  mcm2f_ca_w_1_120_s_0_420=1.49e-05 mcm2f_cc_w_1_120_s_0_420=8.29e-11 mcm2f_cf_w_1_120_s_0_420=3.27e-12
+  mcm2f_ca_w_1_120_s_0_560=1.49e-05 mcm2f_cc_w_1_120_s_0_560=6.95e-11 mcm2f_cf_w_1_120_s_0_560=4.27e-12
+  mcm2f_ca_w_1_120_s_0_840=1.49e-05 mcm2f_cc_w_1_120_s_0_840=5.44e-11 mcm2f_cf_w_1_120_s_0_840=6.18e-12
+  mcm2f_ca_w_1_120_s_1_540=1.49e-05 mcm2f_cc_w_1_120_s_1_540=3.66e-11 mcm2f_cf_w_1_120_s_1_540=1.06e-11
+  mcm2f_ca_w_1_120_s_3_500=1.49e-05 mcm2f_cc_w_1_120_s_3_500=1.89e-11 mcm2f_cf_w_1_120_s_3_500=1.98e-11
+  mcm2d_ca_w_0_140_s_0_140=1.79e-05 mcm2d_cc_w_0_140_s_0_140=9.24e-11 mcm2d_cf_w_0_140_s_0_140=1.44e-12
+  mcm2d_ca_w_0_140_s_0_175=1.79e-05 mcm2d_cc_w_0_140_s_0_175=9.15e-11 mcm2d_cf_w_0_140_s_0_175=1.75e-12
+  mcm2d_ca_w_0_140_s_0_210=1.79e-05 mcm2d_cc_w_0_140_s_0_210=8.76e-11 mcm2d_cf_w_0_140_s_0_210=2.06e-12
+  mcm2d_ca_w_0_140_s_0_280=1.79e-05 mcm2d_cc_w_0_140_s_0_280=7.97e-11 mcm2d_cf_w_0_140_s_0_280=2.67e-12
+  mcm2d_ca_w_0_140_s_0_350=1.79e-05 mcm2d_cc_w_0_140_s_0_350=7.06e-11 mcm2d_cf_w_0_140_s_0_350=3.27e-12
+  mcm2d_ca_w_0_140_s_0_420=1.79e-05 mcm2d_cc_w_0_140_s_0_420=6.26e-11 mcm2d_cf_w_0_140_s_0_420=3.91e-12
+  mcm2d_ca_w_0_140_s_0_560=1.79e-05 mcm2d_cc_w_0_140_s_0_560=5.23e-11 mcm2d_cf_w_0_140_s_0_560=5.05e-12
+  mcm2d_ca_w_0_140_s_0_840=1.79e-05 mcm2d_cc_w_0_140_s_0_840=4.02e-11 mcm2d_cf_w_0_140_s_0_840=7.27e-12
+  mcm2d_ca_w_0_140_s_1_540=1.79e-05 mcm2d_cc_w_0_140_s_1_540=2.60e-11 mcm2d_cf_w_0_140_s_1_540=1.22e-11
+  mcm2d_ca_w_0_140_s_3_500=1.79e-05 mcm2d_cc_w_0_140_s_3_500=1.20e-11 mcm2d_cf_w_0_140_s_3_500=2.12e-11
+  mcm2d_ca_w_1_120_s_0_140=1.79e-05 mcm2d_cc_w_1_120_s_0_140=1.20e-10 mcm2d_cf_w_1_120_s_0_140=1.46e-12
+  mcm2d_ca_w_1_120_s_0_175=1.79e-05 mcm2d_cc_w_1_120_s_0_175=1.17e-10 mcm2d_cf_w_1_120_s_0_175=1.78e-12
+  mcm2d_ca_w_1_120_s_0_210=1.79e-05 mcm2d_cc_w_1_120_s_0_210=1.12e-10 mcm2d_cf_w_1_120_s_0_210=2.09e-12
+  mcm2d_ca_w_1_120_s_0_280=1.79e-05 mcm2d_cc_w_1_120_s_0_280=1.01e-10 mcm2d_cf_w_1_120_s_0_280=2.70e-12
+  mcm2d_ca_w_1_120_s_0_350=1.79e-05 mcm2d_cc_w_1_120_s_0_350=9.03e-11 mcm2d_cf_w_1_120_s_0_350=3.31e-12
+  mcm2d_ca_w_1_120_s_0_420=1.79e-05 mcm2d_cc_w_1_120_s_0_420=8.13e-11 mcm2d_cf_w_1_120_s_0_420=3.91e-12
+  mcm2d_ca_w_1_120_s_0_560=1.79e-05 mcm2d_cc_w_1_120_s_0_560=6.80e-11 mcm2d_cf_w_1_120_s_0_560=5.09e-12
+  mcm2d_ca_w_1_120_s_0_840=1.79e-05 mcm2d_cc_w_1_120_s_0_840=5.27e-11 mcm2d_cf_w_1_120_s_0_840=7.34e-12
+  mcm2d_ca_w_1_120_s_1_540=1.79e-05 mcm2d_cc_w_1_120_s_1_540=3.49e-11 mcm2d_cf_w_1_120_s_1_540=1.24e-11
+  mcm2d_ca_w_1_120_s_3_500=1.79e-05 mcm2d_cc_w_1_120_s_3_500=1.71e-11 mcm2d_cf_w_1_120_s_3_500=2.25e-11
+  mcm2p1_ca_w_0_140_s_0_140=2.04e-05 mcm2p1_cc_w_0_140_s_0_140=9.21e-11 mcm2p1_cf_w_0_140_s_0_140=1.64e-12
+  mcm2p1_ca_w_0_140_s_0_175=2.04e-05 mcm2p1_cc_w_0_140_s_0_175=9.12e-11 mcm2p1_cf_w_0_140_s_0_175=2.00e-12
+  mcm2p1_ca_w_0_140_s_0_210=2.04e-05 mcm2p1_cc_w_0_140_s_0_210=8.73e-11 mcm2p1_cf_w_0_140_s_0_210=2.35e-12
+  mcm2p1_ca_w_0_140_s_0_280=2.04e-05 mcm2p1_cc_w_0_140_s_0_280=7.93e-11 mcm2p1_cf_w_0_140_s_0_280=3.05e-12
+  mcm2p1_ca_w_0_140_s_0_350=2.04e-05 mcm2p1_cc_w_0_140_s_0_350=7.00e-11 mcm2p1_cf_w_0_140_s_0_350=3.73e-12
+  mcm2p1_ca_w_0_140_s_0_420=2.04e-05 mcm2p1_cc_w_0_140_s_0_420=6.23e-11 mcm2p1_cf_w_0_140_s_0_420=4.45e-12
+  mcm2p1_ca_w_0_140_s_0_560=2.04e-05 mcm2p1_cc_w_0_140_s_0_560=5.15e-11 mcm2p1_cf_w_0_140_s_0_560=5.73e-12
+  mcm2p1_ca_w_0_140_s_0_840=2.04e-05 mcm2p1_cc_w_0_140_s_0_840=3.94e-11 mcm2p1_cf_w_0_140_s_0_840=8.23e-12
+  mcm2p1_ca_w_0_140_s_1_540=2.04e-05 mcm2p1_cc_w_0_140_s_1_540=2.50e-11 mcm2p1_cf_w_0_140_s_1_540=1.37e-11
+  mcm2p1_ca_w_0_140_s_3_500=2.04e-05 mcm2p1_cc_w_0_140_s_3_500=1.10e-11 mcm2p1_cf_w_0_140_s_3_500=2.31e-11
+  mcm2p1_ca_w_1_120_s_0_140=2.04e-05 mcm2p1_cc_w_1_120_s_0_140=1.19e-10 mcm2p1_cf_w_1_120_s_0_140=1.69e-12
+  mcm2p1_ca_w_1_120_s_0_175=2.04e-05 mcm2p1_cc_w_1_120_s_0_175=1.16e-10 mcm2p1_cf_w_1_120_s_0_175=2.04e-12
+  mcm2p1_ca_w_1_120_s_0_210=2.04e-05 mcm2p1_cc_w_1_120_s_0_210=1.11e-10 mcm2p1_cf_w_1_120_s_0_210=2.39e-12
+  mcm2p1_ca_w_1_120_s_0_280=2.04e-05 mcm2p1_cc_w_1_120_s_0_280=1.00e-10 mcm2p1_cf_w_1_120_s_0_280=3.09e-12
+  mcm2p1_ca_w_1_120_s_0_350=2.04e-05 mcm2p1_cc_w_1_120_s_0_350=8.91e-11 mcm2p1_cf_w_1_120_s_0_350=3.78e-12
+  mcm2p1_ca_w_1_120_s_0_420=2.04e-05 mcm2p1_cc_w_1_120_s_0_420=7.98e-11 mcm2p1_cf_w_1_120_s_0_420=4.46e-12
+  mcm2p1_ca_w_1_120_s_0_560=2.04e-05 mcm2p1_cc_w_1_120_s_0_560=6.68e-11 mcm2p1_cf_w_1_120_s_0_560=5.80e-12
+  mcm2p1_ca_w_1_120_s_0_840=2.04e-05 mcm2p1_cc_w_1_120_s_0_840=5.14e-11 mcm2p1_cf_w_1_120_s_0_840=8.32e-12
+  mcm2p1_ca_w_1_120_s_1_540=2.04e-05 mcm2p1_cc_w_1_120_s_1_540=3.35e-11 mcm2p1_cf_w_1_120_s_1_540=1.39e-11
+  mcm2p1_ca_w_1_120_s_3_500=2.04e-05 mcm2p1_cc_w_1_120_s_3_500=1.59e-11 mcm2p1_cf_w_1_120_s_3_500=2.47e-11
+  mcm2l1_ca_w_0_140_s_0_140=3.10e-05 mcm2l1_cc_w_0_140_s_0_140=9.10e-11 mcm2l1_cf_w_0_140_s_0_140=2.45e-12
+  mcm2l1_ca_w_0_140_s_0_175=3.10e-05 mcm2l1_cc_w_0_140_s_0_175=8.99e-11 mcm2l1_cf_w_0_140_s_0_175=2.98e-12
+  mcm2l1_ca_w_0_140_s_0_210=3.10e-05 mcm2l1_cc_w_0_140_s_0_210=8.63e-11 mcm2l1_cf_w_0_140_s_0_210=3.53e-12
+  mcm2l1_ca_w_0_140_s_0_280=3.10e-05 mcm2l1_cc_w_0_140_s_0_280=7.73e-11 mcm2l1_cf_w_0_140_s_0_280=4.57e-12
+  mcm2l1_ca_w_0_140_s_0_350=3.10e-05 mcm2l1_cc_w_0_140_s_0_350=6.82e-11 mcm2l1_cf_w_0_140_s_0_350=5.60e-12
+  mcm2l1_ca_w_0_140_s_0_420=3.10e-05 mcm2l1_cc_w_0_140_s_0_420=6.01e-11 mcm2l1_cf_w_0_140_s_0_420=6.62e-12
+  mcm2l1_ca_w_0_140_s_0_560=3.10e-05 mcm2l1_cc_w_0_140_s_0_560=4.91e-11 mcm2l1_cf_w_0_140_s_0_560=8.53e-12
+  mcm2l1_ca_w_0_140_s_0_840=3.10e-05 mcm2l1_cc_w_0_140_s_0_840=3.64e-11 mcm2l1_cf_w_0_140_s_0_840=1.20e-11
+  mcm2l1_ca_w_0_140_s_1_540=3.10e-05 mcm2l1_cc_w_0_140_s_1_540=2.14e-11 mcm2l1_cf_w_0_140_s_1_540=1.92e-11
+  mcm2l1_ca_w_0_140_s_3_500=3.10e-05 mcm2l1_cc_w_0_140_s_3_500=8.11e-12 mcm2l1_cf_w_0_140_s_3_500=2.96e-11
+  mcm2l1_ca_w_1_120_s_0_140=3.10e-05 mcm2l1_cc_w_1_120_s_0_140=1.15e-10 mcm2l1_cf_w_1_120_s_0_140=2.48e-12
+  mcm2l1_ca_w_1_120_s_0_175=3.10e-05 mcm2l1_cc_w_1_120_s_0_175=1.13e-10 mcm2l1_cf_w_1_120_s_0_175=3.02e-12
+  mcm2l1_ca_w_1_120_s_0_210=3.10e-05 mcm2l1_cc_w_1_120_s_0_210=1.07e-10 mcm2l1_cf_w_1_120_s_0_210=3.55e-12
+  mcm2l1_ca_w_1_120_s_0_280=3.10e-05 mcm2l1_cc_w_1_120_s_0_280=9.60e-11 mcm2l1_cf_w_1_120_s_0_280=4.60e-12
+  mcm2l1_ca_w_1_120_s_0_350=3.10e-05 mcm2l1_cc_w_1_120_s_0_350=8.53e-11 mcm2l1_cf_w_1_120_s_0_350=5.63e-12
+  mcm2l1_ca_w_1_120_s_0_420=3.10e-05 mcm2l1_cc_w_1_120_s_0_420=7.59e-11 mcm2l1_cf_w_1_120_s_0_420=6.63e-12
+  mcm2l1_ca_w_1_120_s_0_560=3.10e-05 mcm2l1_cc_w_1_120_s_0_560=6.26e-11 mcm2l1_cf_w_1_120_s_0_560=8.56e-12
+  mcm2l1_ca_w_1_120_s_0_840=3.10e-05 mcm2l1_cc_w_1_120_s_0_840=4.72e-11 mcm2l1_cf_w_1_120_s_0_840=1.22e-11
+  mcm2l1_ca_w_1_120_s_1_540=3.10e-05 mcm2l1_cc_w_1_120_s_1_540=2.93e-11 mcm2l1_cf_w_1_120_s_1_540=1.97e-11
+  mcm2l1_ca_w_1_120_s_3_500=3.10e-05 mcm2l1_cc_w_1_120_s_3_500=1.26e-11 mcm2l1_cf_w_1_120_s_3_500=3.17e-11
+  mcm2m1_ca_w_0_140_s_0_140=9.04e-05 mcm2m1_cc_w_0_140_s_0_140=8.52e-11 mcm2m1_cf_w_0_140_s_0_140=6.83e-12
+  mcm2m1_ca_w_0_140_s_0_175=9.04e-05 mcm2m1_cc_w_0_140_s_0_175=8.38e-11 mcm2m1_cf_w_0_140_s_0_175=8.38e-12
+  mcm2m1_ca_w_0_140_s_0_210=9.04e-05 mcm2m1_cc_w_0_140_s_0_210=7.94e-11 mcm2m1_cf_w_0_140_s_0_210=9.88e-12
+  mcm2m1_ca_w_0_140_s_0_280=9.04e-05 mcm2m1_cc_w_0_140_s_0_280=6.97e-11 mcm2m1_cf_w_0_140_s_0_280=1.27e-11
+  mcm2m1_ca_w_0_140_s_0_350=9.04e-05 mcm2m1_cc_w_0_140_s_0_350=6.01e-11 mcm2m1_cf_w_0_140_s_0_350=1.54e-11
+  mcm2m1_ca_w_0_140_s_0_420=9.04e-05 mcm2m1_cc_w_0_140_s_0_420=5.14e-11 mcm2m1_cf_w_0_140_s_0_420=1.80e-11
+  mcm2m1_ca_w_0_140_s_0_560=9.04e-05 mcm2m1_cc_w_0_140_s_0_560=4.00e-11 mcm2m1_cf_w_0_140_s_0_560=2.25e-11
+  mcm2m1_ca_w_0_140_s_0_840=9.04e-05 mcm2m1_cc_w_0_140_s_0_840=2.68e-11 mcm2m1_cf_w_0_140_s_0_840=2.96e-11
+  mcm2m1_ca_w_0_140_s_1_540=9.04e-05 mcm2m1_cc_w_0_140_s_1_540=1.28e-11 mcm2m1_cf_w_0_140_s_1_540=4.04e-11
+  mcm2m1_ca_w_0_140_s_3_500=9.04e-05 mcm2m1_cc_w_0_140_s_3_500=3.70e-12 mcm2m1_cf_w_0_140_s_3_500=4.91e-11
+  mcm2m1_ca_w_1_120_s_0_140=9.04e-05 mcm2m1_cc_w_1_120_s_0_140=1.04e-10 mcm2m1_cf_w_1_120_s_0_140=6.83e-12
+  mcm2m1_ca_w_1_120_s_0_175=9.04e-05 mcm2m1_cc_w_1_120_s_0_175=1.01e-10 mcm2m1_cf_w_1_120_s_0_175=8.40e-12
+  mcm2m1_ca_w_1_120_s_0_210=9.04e-05 mcm2m1_cc_w_1_120_s_0_210=9.61e-11 mcm2m1_cf_w_1_120_s_0_210=9.90e-12
+  mcm2m1_ca_w_1_120_s_0_280=9.04e-05 mcm2m1_cc_w_1_120_s_0_280=8.44e-11 mcm2m1_cf_w_1_120_s_0_280=1.27e-11
+  mcm2m1_ca_w_1_120_s_0_350=9.04e-05 mcm2m1_cc_w_1_120_s_0_350=7.37e-11 mcm2m1_cf_w_1_120_s_0_350=1.54e-11
+  mcm2m1_ca_w_1_120_s_0_420=9.04e-05 mcm2m1_cc_w_1_120_s_0_420=6.46e-11 mcm2m1_cf_w_1_120_s_0_420=1.79e-11
+  mcm2m1_ca_w_1_120_s_0_560=9.04e-05 mcm2m1_cc_w_1_120_s_0_560=5.15e-11 mcm2m1_cf_w_1_120_s_0_560=2.25e-11
+  mcm2m1_ca_w_1_120_s_0_840=9.04e-05 mcm2m1_cc_w_1_120_s_0_840=3.65e-11 mcm2m1_cf_w_1_120_s_0_840=2.98e-11
+  mcm2m1_ca_w_1_120_s_1_540=9.04e-05 mcm2m1_cc_w_1_120_s_1_540=2.01e-11 mcm2m1_cf_w_1_120_s_1_540=4.14e-11
+  mcm2m1_ca_w_1_120_s_3_500=9.04e-05 mcm2m1_cc_w_1_120_s_3_500=7.25e-12 mcm2m1_cf_w_1_120_s_3_500=5.32e-11
+  mcm3f_ca_w_0_300_s_0_300=1.08e-05 mcm3f_cc_w_0_300_s_0_300=9.56e-11 mcm3f_cf_w_0_300_s_0_300=1.78e-12
+  mcm3f_ca_w_0_300_s_0_360=1.08e-05 mcm3f_cc_w_0_300_s_0_360=8.99e-11 mcm3f_cf_w_0_300_s_0_360=2.10e-12
+  mcm3f_ca_w_0_300_s_0_450=1.08e-05 mcm3f_cc_w_0_300_s_0_450=8.19e-11 mcm3f_cf_w_0_300_s_0_450=2.59e-12
+  mcm3f_ca_w_0_300_s_0_600=1.08e-05 mcm3f_cc_w_0_300_s_0_600=7.14e-11 mcm3f_cf_w_0_300_s_0_600=3.39e-12
+  mcm3f_ca_w_0_300_s_0_800=1.08e-05 mcm3f_cc_w_0_300_s_0_800=6.12e-11 mcm3f_cf_w_0_300_s_0_800=4.33e-12
+  mcm3f_ca_w_0_300_s_1_000=1.08e-05 mcm3f_cc_w_0_300_s_1_000=5.32e-11 mcm3f_cf_w_0_300_s_1_000=5.31e-12
+  mcm3f_ca_w_0_300_s_1_200=1.08e-05 mcm3f_cc_w_0_300_s_1_200=4.73e-11 mcm3f_cf_w_0_300_s_1_200=6.25e-12
+  mcm3f_ca_w_0_300_s_2_100=1.08e-05 mcm3f_cc_w_0_300_s_2_100=3.18e-11 mcm3f_cf_w_0_300_s_2_100=1.05e-11
+  mcm3f_ca_w_0_300_s_3_300=1.08e-05 mcm3f_cc_w_0_300_s_3_300=2.26e-11 mcm3f_cf_w_0_300_s_3_300=1.46e-11
+  mcm3f_ca_w_0_300_s_9_000=1.08e-05 mcm3f_cc_w_0_300_s_9_000=7.21e-12 mcm3f_cf_w_0_300_s_9_000=2.58e-11
+  mcm3f_ca_w_2_400_s_0_300=1.08e-05 mcm3f_cc_w_2_400_s_0_300=1.22e-10 mcm3f_cf_w_2_400_s_0_300=1.81e-12
+  mcm3f_ca_w_2_400_s_0_360=1.08e-05 mcm3f_cc_w_2_400_s_0_360=1.14e-10 mcm3f_cf_w_2_400_s_0_360=2.13e-12
+  mcm3f_ca_w_2_400_s_0_450=1.08e-05 mcm3f_cc_w_2_400_s_0_450=1.05e-10 mcm3f_cf_w_2_400_s_0_450=2.60e-12
+  mcm3f_ca_w_2_400_s_0_600=1.08e-05 mcm3f_cc_w_2_400_s_0_600=9.22e-11 mcm3f_cf_w_2_400_s_0_600=3.37e-12
+  mcm3f_ca_w_2_400_s_0_800=1.08e-05 mcm3f_cc_w_2_400_s_0_800=7.94e-11 mcm3f_cf_w_2_400_s_0_800=4.38e-12
+  mcm3f_ca_w_2_400_s_1_000=1.08e-05 mcm3f_cc_w_2_400_s_1_000=6.97e-11 mcm3f_cf_w_2_400_s_1_000=5.37e-12
+  mcm3f_ca_w_2_400_s_1_200=1.08e-05 mcm3f_cc_w_2_400_s_1_200=6.23e-11 mcm3f_cf_w_2_400_s_1_200=6.34e-12
+  mcm3f_ca_w_2_400_s_2_100=1.08e-05 mcm3f_cc_w_2_400_s_2_100=4.33e-11 mcm3f_cf_w_2_400_s_2_100=1.04e-11
+  mcm3f_ca_w_2_400_s_3_300=1.08e-05 mcm3f_cc_w_2_400_s_3_300=3.10e-11 mcm3f_cf_w_2_400_s_3_300=1.51e-11
+  mcm3f_ca_w_2_400_s_9_000=1.08e-05 mcm3f_cc_w_2_400_s_9_000=1.11e-11 mcm3f_cf_w_2_400_s_9_000=2.84e-11
+  mcm3d_ca_w_0_300_s_0_300=1.23e-05 mcm3d_cc_w_0_300_s_0_300=9.52e-11 mcm3d_cf_w_0_300_s_0_300=2.02e-12
+  mcm3d_ca_w_0_300_s_0_360=1.23e-05 mcm3d_cc_w_0_300_s_0_360=8.95e-11 mcm3d_cf_w_0_300_s_0_360=2.38e-12
+  mcm3d_ca_w_0_300_s_0_450=1.23e-05 mcm3d_cc_w_0_300_s_0_450=8.15e-11 mcm3d_cf_w_0_300_s_0_450=2.93e-12
+  mcm3d_ca_w_0_300_s_0_600=1.23e-05 mcm3d_cc_w_0_300_s_0_600=7.08e-11 mcm3d_cf_w_0_300_s_0_600=3.84e-12
+  mcm3d_ca_w_0_300_s_0_800=1.23e-05 mcm3d_cc_w_0_300_s_0_800=6.06e-11 mcm3d_cf_w_0_300_s_0_800=4.90e-12
+  mcm3d_ca_w_0_300_s_1_000=1.23e-05 mcm3d_cc_w_0_300_s_1_000=5.26e-11 mcm3d_cf_w_0_300_s_1_000=6.00e-12
+  mcm3d_ca_w_0_300_s_1_200=1.23e-05 mcm3d_cc_w_0_300_s_1_200=4.64e-11 mcm3d_cf_w_0_300_s_1_200=7.06e-12
+  mcm3d_ca_w_0_300_s_2_100=1.23e-05 mcm3d_cc_w_0_300_s_2_100=3.09e-11 mcm3d_cf_w_0_300_s_2_100=1.17e-11
+  mcm3d_ca_w_0_300_s_3_300=1.23e-05 mcm3d_cc_w_0_300_s_3_300=2.15e-11 mcm3d_cf_w_0_300_s_3_300=1.62e-11
+  mcm3d_ca_w_0_300_s_9_000=1.23e-05 mcm3d_cc_w_0_300_s_9_000=6.51e-12 mcm3d_cf_w_0_300_s_9_000=2.75e-11
+  mcm3d_ca_w_2_400_s_0_300=1.23e-05 mcm3d_cc_w_2_400_s_0_300=1.20e-10 mcm3d_cf_w_2_400_s_0_300=2.06e-12
+  mcm3d_ca_w_2_400_s_0_360=1.23e-05 mcm3d_cc_w_2_400_s_0_360=1.13e-10 mcm3d_cf_w_2_400_s_0_360=2.42e-12
+  mcm3d_ca_w_2_400_s_0_450=1.23e-05 mcm3d_cc_w_2_400_s_0_450=1.04e-10 mcm3d_cf_w_2_400_s_0_450=2.95e-12
+  mcm3d_ca_w_2_400_s_0_600=1.23e-05 mcm3d_cc_w_2_400_s_0_600=9.09e-11 mcm3d_cf_w_2_400_s_0_600=3.82e-12
+  mcm3d_ca_w_2_400_s_0_800=1.23e-05 mcm3d_cc_w_2_400_s_0_800=7.81e-11 mcm3d_cf_w_2_400_s_0_800=4.96e-12
+  mcm3d_ca_w_2_400_s_1_000=1.23e-05 mcm3d_cc_w_2_400_s_1_000=6.84e-11 mcm3d_cf_w_2_400_s_1_000=6.07e-12
+  mcm3d_ca_w_2_400_s_1_200=1.23e-05 mcm3d_cc_w_2_400_s_1_200=6.10e-11 mcm3d_cf_w_2_400_s_1_200=7.16e-12
+  mcm3d_ca_w_2_400_s_2_100=1.23e-05 mcm3d_cc_w_2_400_s_2_100=4.20e-11 mcm3d_cf_w_2_400_s_2_100=1.17e-11
+  mcm3d_ca_w_2_400_s_3_300=1.23e-05 mcm3d_cc_w_2_400_s_3_300=2.98e-11 mcm3d_cf_w_2_400_s_3_300=1.67e-11
+  mcm3d_ca_w_2_400_s_9_000=1.23e-05 mcm3d_cc_w_2_400_s_9_000=1.02e-11 mcm3d_cf_w_2_400_s_9_000=3.04e-11
+  mcm3p1_ca_w_0_300_s_0_300=1.35e-05 mcm3p1_cc_w_0_300_s_0_300=9.49e-11 mcm3p1_cf_w_0_300_s_0_300=2.21e-12
+  mcm3p1_ca_w_0_300_s_0_360=1.35e-05 mcm3p1_cc_w_0_300_s_0_360=8.92e-11 mcm3p1_cf_w_0_300_s_0_360=2.60e-12
+  mcm3p1_ca_w_0_300_s_0_450=1.35e-05 mcm3p1_cc_w_0_300_s_0_450=8.12e-11 mcm3p1_cf_w_0_300_s_0_450=3.20e-12
+  mcm3p1_ca_w_0_300_s_0_600=1.35e-05 mcm3p1_cc_w_0_300_s_0_600=7.04e-11 mcm3p1_cf_w_0_300_s_0_600=4.18e-12
+  mcm3p1_ca_w_0_300_s_0_800=1.35e-05 mcm3p1_cc_w_0_300_s_0_800=6.01e-11 mcm3p1_cf_w_0_300_s_0_800=5.34e-12
+  mcm3p1_ca_w_0_300_s_1_000=1.35e-05 mcm3p1_cc_w_0_300_s_1_000=5.20e-11 mcm3p1_cf_w_0_300_s_1_000=6.53e-12
+  mcm3p1_ca_w_0_300_s_1_200=1.35e-05 mcm3p1_cc_w_0_300_s_1_200=4.59e-11 mcm3p1_cf_w_0_300_s_1_200=7.68e-12
+  mcm3p1_ca_w_0_300_s_2_100=1.35e-05 mcm3p1_cc_w_0_300_s_2_100=3.02e-11 mcm3p1_cf_w_0_300_s_2_100=1.27e-11
+  mcm3p1_ca_w_0_300_s_3_300=1.35e-05 mcm3p1_cc_w_0_300_s_3_300=2.08e-11 mcm3p1_cf_w_0_300_s_3_300=1.74e-11
+  mcm3p1_ca_w_0_300_s_9_000=1.35e-05 mcm3p1_cc_w_0_300_s_9_000=6.03e-12 mcm3p1_cf_w_0_300_s_9_000=2.88e-11
+  mcm3p1_ca_w_2_400_s_0_300=1.35e-05 mcm3p1_cc_w_2_400_s_0_300=1.20e-10 mcm3p1_cf_w_2_400_s_0_300=2.27e-12
+  mcm3p1_ca_w_2_400_s_0_360=1.35e-05 mcm3p1_cc_w_2_400_s_0_360=1.12e-10 mcm3p1_cf_w_2_400_s_0_360=2.66e-12
+  mcm3p1_ca_w_2_400_s_0_450=1.35e-05 mcm3p1_cc_w_2_400_s_0_450=1.03e-10 mcm3p1_cf_w_2_400_s_0_450=3.24e-12
+  mcm3p1_ca_w_2_400_s_0_600=1.35e-05 mcm3p1_cc_w_2_400_s_0_600=9.00e-11 mcm3p1_cf_w_2_400_s_0_600=4.18e-12
+  mcm3p1_ca_w_2_400_s_0_800=1.35e-05 mcm3p1_cc_w_2_400_s_0_800=7.72e-11 mcm3p1_cf_w_2_400_s_0_800=5.42e-12
+  mcm3p1_ca_w_2_400_s_1_000=1.35e-05 mcm3p1_cc_w_2_400_s_1_000=6.75e-11 mcm3p1_cf_w_2_400_s_1_000=6.62e-12
+  mcm3p1_ca_w_2_400_s_1_200=1.35e-05 mcm3p1_cc_w_2_400_s_1_200=6.01e-11 mcm3p1_cf_w_2_400_s_1_200=7.80e-12
+  mcm3p1_ca_w_2_400_s_2_100=1.35e-05 mcm3p1_cc_w_2_400_s_2_100=4.11e-11 mcm3p1_cf_w_2_400_s_2_100=1.26e-11
+  mcm3p1_ca_w_2_400_s_3_300=1.35e-05 mcm3p1_cc_w_2_400_s_3_300=2.89e-11 mcm3p1_cf_w_2_400_s_3_300=1.80e-11
+  mcm3p1_ca_w_2_400_s_9_000=1.35e-05 mcm3p1_cc_w_2_400_s_9_000=9.69e-12 mcm3p1_cf_w_2_400_s_9_000=3.18e-11
+  mcm3l1_ca_w_0_300_s_0_300=1.74e-05 mcm3l1_cc_w_0_300_s_0_300=9.40e-11 mcm3l1_cf_w_0_300_s_0_300=2.83e-12
+  mcm3l1_ca_w_0_300_s_0_360=1.74e-05 mcm3l1_cc_w_0_300_s_0_360=8.82e-11 mcm3l1_cf_w_0_300_s_0_360=3.32e-12
+  mcm3l1_ca_w_0_300_s_0_450=1.74e-05 mcm3l1_cc_w_0_300_s_0_450=8.00e-11 mcm3l1_cf_w_0_300_s_0_450=4.08e-12
+  mcm3l1_ca_w_0_300_s_0_600=1.74e-05 mcm3l1_cc_w_0_300_s_0_600=6.92e-11 mcm3l1_cf_w_0_300_s_0_600=5.30e-12
+  mcm3l1_ca_w_0_300_s_0_800=1.74e-05 mcm3l1_cc_w_0_300_s_0_800=5.86e-11 mcm3l1_cf_w_0_300_s_0_800=6.76e-12
+  mcm3l1_ca_w_0_300_s_1_000=1.74e-05 mcm3l1_cc_w_0_300_s_1_000=5.04e-11 mcm3l1_cf_w_0_300_s_1_000=8.24e-12
+  mcm3l1_ca_w_0_300_s_1_200=1.74e-05 mcm3l1_cc_w_0_300_s_1_200=4.42e-11 mcm3l1_cf_w_0_300_s_1_200=9.65e-12
+  mcm3l1_ca_w_0_300_s_2_100=1.74e-05 mcm3l1_cc_w_0_300_s_2_100=2.80e-11 mcm3l1_cf_w_0_300_s_2_100=1.56e-11
+  mcm3l1_ca_w_0_300_s_3_300=1.74e-05 mcm3l1_cc_w_0_300_s_3_300=1.87e-11 mcm3l1_cf_w_0_300_s_3_300=2.09e-11
+  mcm3l1_ca_w_0_300_s_9_000=1.74e-05 mcm3l1_cc_w_0_300_s_9_000=4.94e-12 mcm3l1_cf_w_0_300_s_9_000=3.22e-11
+  mcm3l1_ca_w_2_400_s_0_300=1.74e-05 mcm3l1_cc_w_2_400_s_0_300=1.17e-10 mcm3l1_cf_w_2_400_s_0_300=2.86e-12
+  mcm3l1_ca_w_2_400_s_0_360=1.74e-05 mcm3l1_cc_w_2_400_s_0_360=1.10e-10 mcm3l1_cf_w_2_400_s_0_360=3.35e-12
+  mcm3l1_ca_w_2_400_s_0_450=1.74e-05 mcm3l1_cc_w_2_400_s_0_450=1.00e-10 mcm3l1_cf_w_2_400_s_0_450=4.09e-12
+  mcm3l1_ca_w_2_400_s_0_600=1.74e-05 mcm3l1_cc_w_2_400_s_0_600=8.74e-11 mcm3l1_cf_w_2_400_s_0_600=5.28e-12
+  mcm3l1_ca_w_2_400_s_0_800=1.74e-05 mcm3l1_cc_w_2_400_s_0_800=7.46e-11 mcm3l1_cf_w_2_400_s_0_800=6.83e-12
+  mcm3l1_ca_w_2_400_s_1_000=1.74e-05 mcm3l1_cc_w_2_400_s_1_000=6.48e-11 mcm3l1_cf_w_2_400_s_1_000=8.33e-12
+  mcm3l1_ca_w_2_400_s_1_200=1.74e-05 mcm3l1_cc_w_2_400_s_1_200=5.74e-11 mcm3l1_cf_w_2_400_s_1_200=9.76e-12
+  mcm3l1_ca_w_2_400_s_2_100=1.74e-05 mcm3l1_cc_w_2_400_s_2_100=3.84e-11 mcm3l1_cf_w_2_400_s_2_100=1.56e-11
+  mcm3l1_ca_w_2_400_s_3_300=1.74e-05 mcm3l1_cc_w_2_400_s_3_300=2.64e-11 mcm3l1_cf_w_2_400_s_3_300=2.17e-11
+  mcm3l1_ca_w_2_400_s_9_000=1.74e-05 mcm3l1_cc_w_2_400_s_9_000=8.25e-12 mcm3l1_cf_w_2_400_s_9_000=3.58e-11
+  mcm3m1_ca_w_0_300_s_0_300=2.75e-05 mcm3m1_cc_w_0_300_s_0_300=9.16e-11 mcm3m1_cf_w_0_300_s_0_300=4.41e-12
+  mcm3m1_ca_w_0_300_s_0_360=2.75e-05 mcm3m1_cc_w_0_300_s_0_360=8.54e-11 mcm3m1_cf_w_0_300_s_0_360=5.16e-12
+  mcm3m1_ca_w_0_300_s_0_450=2.75e-05 mcm3m1_cc_w_0_300_s_0_450=7.73e-11 mcm3m1_cf_w_0_300_s_0_450=6.30e-12
+  mcm3m1_ca_w_0_300_s_0_600=2.75e-05 mcm3m1_cc_w_0_300_s_0_600=6.62e-11 mcm3m1_cf_w_0_300_s_0_600=8.11e-12
+  mcm3m1_ca_w_0_300_s_0_800=2.75e-05 mcm3m1_cc_w_0_300_s_0_800=5.52e-11 mcm3m1_cf_w_0_300_s_0_800=1.03e-11
+  mcm3m1_ca_w_0_300_s_1_000=2.75e-05 mcm3m1_cc_w_0_300_s_1_000=4.69e-11 mcm3m1_cf_w_0_300_s_1_000=1.24e-11
+  mcm3m1_ca_w_0_300_s_1_200=2.75e-05 mcm3m1_cc_w_0_300_s_1_200=4.05e-11 mcm3m1_cf_w_0_300_s_1_200=1.44e-11
+  mcm3m1_ca_w_0_300_s_2_100=2.75e-05 mcm3m1_cc_w_0_300_s_2_100=2.41e-11 mcm3m1_cf_w_0_300_s_2_100=2.23e-11
+  mcm3m1_ca_w_0_300_s_3_300=2.75e-05 mcm3m1_cc_w_0_300_s_3_300=1.51e-11 mcm3m1_cf_w_0_300_s_3_300=2.84e-11
+  mcm3m1_ca_w_0_300_s_9_000=2.75e-05 mcm3m1_cc_w_0_300_s_9_000=3.43e-12 mcm3m1_cf_w_0_300_s_9_000=3.87e-11
+  mcm3m1_ca_w_2_400_s_0_300=2.75e-05 mcm3m1_cc_w_2_400_s_0_300=1.12e-10 mcm3m1_cf_w_2_400_s_0_300=4.42e-12
+  mcm3m1_ca_w_2_400_s_0_360=2.75e-05 mcm3m1_cc_w_2_400_s_0_360=1.05e-10 mcm3m1_cf_w_2_400_s_0_360=5.18e-12
+  mcm3m1_ca_w_2_400_s_0_450=2.75e-05 mcm3m1_cc_w_2_400_s_0_450=9.54e-11 mcm3m1_cf_w_2_400_s_0_450=6.30e-12
+  mcm3m1_ca_w_2_400_s_0_600=2.75e-05 mcm3m1_cc_w_2_400_s_0_600=8.25e-11 mcm3m1_cf_w_2_400_s_0_600=8.09e-12
+  mcm3m1_ca_w_2_400_s_0_800=2.75e-05 mcm3m1_cc_w_2_400_s_0_800=6.98e-11 mcm3m1_cf_w_2_400_s_0_800=1.04e-11
+  mcm3m1_ca_w_2_400_s_1_000=2.75e-05 mcm3m1_cc_w_2_400_s_1_000=6.01e-11 mcm3m1_cf_w_2_400_s_1_000=1.25e-11
+  mcm3m1_ca_w_2_400_s_1_200=2.75e-05 mcm3m1_cc_w_2_400_s_1_200=5.27e-11 mcm3m1_cf_w_2_400_s_1_200=1.45e-11
+  mcm3m1_ca_w_2_400_s_2_100=2.75e-05 mcm3m1_cc_w_2_400_s_2_100=3.40e-11 mcm3m1_cf_w_2_400_s_2_100=2.22e-11
+  mcm3m1_ca_w_2_400_s_3_300=2.75e-05 mcm3m1_cc_w_2_400_s_3_300=2.23e-11 mcm3m1_cf_w_2_400_s_3_300=2.95e-11
+  mcm3m1_ca_w_2_400_s_9_000=2.75e-05 mcm3m1_cc_w_2_400_s_9_000=6.30e-12 mcm3m1_cf_w_2_400_s_9_000=4.32e-11
+  mcm3m2_ca_w_0_300_s_0_300=6.49e-05 mcm3m2_cc_w_0_300_s_0_300=8.47e-11 mcm3m2_cf_w_0_300_s_0_300=9.82e-12
+  mcm3m2_ca_w_0_300_s_0_360=6.49e-05 mcm3m2_cc_w_0_300_s_0_360=7.86e-11 mcm3m2_cf_w_0_300_s_0_360=1.14e-11
+  mcm3m2_ca_w_0_300_s_0_450=6.49e-05 mcm3m2_cc_w_0_300_s_0_450=7.02e-11 mcm3m2_cf_w_0_300_s_0_450=1.36e-11
+  mcm3m2_ca_w_0_300_s_0_600=6.49e-05 mcm3m2_cc_w_0_300_s_0_600=5.87e-11 mcm3m2_cf_w_0_300_s_0_600=1.72e-11
+  mcm3m2_ca_w_0_300_s_0_800=6.49e-05 mcm3m2_cc_w_0_300_s_0_800=4.78e-11 mcm3m2_cf_w_0_300_s_0_800=2.11e-11
+  mcm3m2_ca_w_0_300_s_1_000=6.49e-05 mcm3m2_cc_w_0_300_s_1_000=3.94e-11 mcm3m2_cf_w_0_300_s_1_000=2.47e-11
+  mcm3m2_ca_w_0_300_s_1_200=6.49e-05 mcm3m2_cc_w_0_300_s_1_200=3.31e-11 mcm3m2_cf_w_0_300_s_1_200=2.78e-11
+  mcm3m2_ca_w_0_300_s_2_100=6.49e-05 mcm3m2_cc_w_0_300_s_2_100=1.74e-11 mcm3m2_cf_w_0_300_s_2_100=3.82e-11
+  mcm3m2_ca_w_0_300_s_3_300=6.49e-05 mcm3m2_cc_w_0_300_s_3_300=9.90e-12 mcm3m2_cf_w_0_300_s_3_300=4.44e-11
+  mcm3m2_ca_w_0_300_s_9_000=6.49e-05 mcm3m2_cc_w_0_300_s_9_000=2.00e-12 mcm3m2_cf_w_0_300_s_9_000=5.20e-11
+  mcm3m2_ca_w_2_400_s_0_300=6.49e-05 mcm3m2_cc_w_2_400_s_0_300=1.02e-10 mcm3m2_cf_w_2_400_s_0_300=9.84e-12
+  mcm3m2_ca_w_2_400_s_0_360=6.49e-05 mcm3m2_cc_w_2_400_s_0_360=9.55e-11 mcm3m2_cf_w_2_400_s_0_360=1.14e-11
+  mcm3m2_ca_w_2_400_s_0_450=6.49e-05 mcm3m2_cc_w_2_400_s_0_450=8.62e-11 mcm3m2_cf_w_2_400_s_0_450=1.37e-11
+  mcm3m2_ca_w_2_400_s_0_600=6.49e-05 mcm3m2_cc_w_2_400_s_0_600=7.35e-11 mcm3m2_cf_w_2_400_s_0_600=1.71e-11
+  mcm3m2_ca_w_2_400_s_0_800=6.49e-05 mcm3m2_cc_w_2_400_s_0_800=6.10e-11 mcm3m2_cf_w_2_400_s_0_800=2.12e-11
+  mcm3m2_ca_w_2_400_s_1_000=6.49e-05 mcm3m2_cc_w_2_400_s_1_000=5.16e-11 mcm3m2_cf_w_2_400_s_1_000=2.47e-11
+  mcm3m2_ca_w_2_400_s_1_200=6.49e-05 mcm3m2_cc_w_2_400_s_1_200=4.46e-11 mcm3m2_cf_w_2_400_s_1_200=2.79e-11
+  mcm3m2_ca_w_2_400_s_2_100=6.49e-05 mcm3m2_cc_w_2_400_s_2_100=2.71e-11 mcm3m2_cf_w_2_400_s_2_100=3.82e-11
+  mcm3m2_ca_w_2_400_s_3_300=6.49e-05 mcm3m2_cc_w_2_400_s_3_300=1.69e-11 mcm3m2_cf_w_2_400_s_3_300=4.61e-11
+  mcm3m2_ca_w_2_400_s_9_000=6.49e-05 mcm3m2_cc_w_2_400_s_9_000=4.30e-12 mcm3m2_cf_w_2_400_s_9_000=5.78e-11
+  mcm4f_ca_w_0_300_s_0_300=7.66e-06 mcm4f_cc_w_0_300_s_0_300=9.68e-11 mcm4f_cf_w_0_300_s_0_300=1.26e-12
+  mcm4f_ca_w_0_300_s_0_360=7.66e-06 mcm4f_cc_w_0_300_s_0_360=9.10e-11 mcm4f_cf_w_0_300_s_0_360=1.49e-12
+  mcm4f_ca_w_0_300_s_0_450=7.66e-06 mcm4f_cc_w_0_300_s_0_450=8.31e-11 mcm4f_cf_w_0_300_s_0_450=1.84e-12
+  mcm4f_ca_w_0_300_s_0_600=7.66e-06 mcm4f_cc_w_0_300_s_0_600=7.29e-11 mcm4f_cf_w_0_300_s_0_600=2.42e-12
+  mcm4f_ca_w_0_300_s_0_800=7.66e-06 mcm4f_cc_w_0_300_s_0_800=6.29e-11 mcm4f_cf_w_0_300_s_0_800=3.09e-12
+  mcm4f_ca_w_0_300_s_1_000=7.66e-06 mcm4f_cc_w_0_300_s_1_000=5.52e-11 mcm4f_cf_w_0_300_s_1_000=3.79e-12
+  mcm4f_ca_w_0_300_s_1_200=7.66e-06 mcm4f_cc_w_0_300_s_1_200=4.93e-11 mcm4f_cf_w_0_300_s_1_200=4.49e-12
+  mcm4f_ca_w_0_300_s_2_100=7.66e-06 mcm4f_cc_w_0_300_s_2_100=3.45e-11 mcm4f_cf_w_0_300_s_2_100=7.71e-12
+  mcm4f_ca_w_0_300_s_3_300=7.66e-06 mcm4f_cc_w_0_300_s_3_300=2.53e-11 mcm4f_cf_w_0_300_s_3_300=1.09e-11
+  mcm4f_ca_w_0_300_s_9_000=7.66e-06 mcm4f_cc_w_0_300_s_9_000=9.24e-12 mcm4f_cf_w_0_300_s_9_000=2.12e-11
+  mcm4f_ca_w_2_400_s_0_300=7.66e-06 mcm4f_cc_w_2_400_s_0_300=1.25e-10 mcm4f_cf_w_2_400_s_0_300=1.28e-12
+  mcm4f_ca_w_2_400_s_0_360=7.66e-06 mcm4f_cc_w_2_400_s_0_360=1.18e-10 mcm4f_cf_w_2_400_s_0_360=1.50e-12
+  mcm4f_ca_w_2_400_s_0_450=7.66e-06 mcm4f_cc_w_2_400_s_0_450=1.09e-10 mcm4f_cf_w_2_400_s_0_450=1.84e-12
+  mcm4f_ca_w_2_400_s_0_600=7.66e-06 mcm4f_cc_w_2_400_s_0_600=9.60e-11 mcm4f_cf_w_2_400_s_0_600=2.39e-12
+  mcm4f_ca_w_2_400_s_0_800=7.66e-06 mcm4f_cc_w_2_400_s_0_800=8.30e-11 mcm4f_cf_w_2_400_s_0_800=3.12e-12
+  mcm4f_ca_w_2_400_s_1_000=7.66e-06 mcm4f_cc_w_2_400_s_1_000=7.34e-11 mcm4f_cf_w_2_400_s_1_000=3.84e-12
+  mcm4f_ca_w_2_400_s_1_200=7.66e-06 mcm4f_cc_w_2_400_s_1_200=6.60e-11 mcm4f_cf_w_2_400_s_1_200=4.54e-12
+  mcm4f_ca_w_2_400_s_2_100=7.66e-06 mcm4f_cc_w_2_400_s_2_100=4.67e-11 mcm4f_cf_w_2_400_s_2_100=7.57e-12
+  mcm4f_ca_w_2_400_s_3_300=7.66e-06 mcm4f_cc_w_2_400_s_3_300=3.43e-11 mcm4f_cf_w_2_400_s_3_300=1.12e-11
+  mcm4f_ca_w_2_400_s_9_000=7.66e-06 mcm4f_cc_w_2_400_s_9_000=1.35e-11 mcm4f_cf_w_2_400_s_9_000=2.31e-11
+  mcm4d_ca_w_0_300_s_0_300=8.37e-06 mcm4d_cc_w_0_300_s_0_300=9.66e-11 mcm4d_cf_w_0_300_s_0_300=1.38e-12
+  mcm4d_ca_w_0_300_s_0_360=8.37e-06 mcm4d_cc_w_0_300_s_0_360=9.08e-11 mcm4d_cf_w_0_300_s_0_360=1.63e-12
+  mcm4d_ca_w_0_300_s_0_450=8.37e-06 mcm4d_cc_w_0_300_s_0_450=8.29e-11 mcm4d_cf_w_0_300_s_0_450=2.01e-12
+  mcm4d_ca_w_0_300_s_0_600=8.37e-06 mcm4d_cc_w_0_300_s_0_600=7.26e-11 mcm4d_cf_w_0_300_s_0_600=2.64e-12
+  mcm4d_ca_w_0_300_s_0_800=8.37e-06 mcm4d_cc_w_0_300_s_0_800=6.26e-11 mcm4d_cf_w_0_300_s_0_800=3.37e-12
+  mcm4d_ca_w_0_300_s_1_000=8.37e-06 mcm4d_cc_w_0_300_s_1_000=5.48e-11 mcm4d_cf_w_0_300_s_1_000=4.13e-12
+  mcm4d_ca_w_0_300_s_1_200=8.37e-06 mcm4d_cc_w_0_300_s_1_200=4.89e-11 mcm4d_cf_w_0_300_s_1_200=4.89e-12
+  mcm4d_ca_w_0_300_s_2_100=8.37e-06 mcm4d_cc_w_0_300_s_2_100=3.40e-11 mcm4d_cf_w_0_300_s_2_100=8.33e-12
+  mcm4d_ca_w_0_300_s_3_300=8.37e-06 mcm4d_cc_w_0_300_s_3_300=2.47e-11 mcm4d_cf_w_0_300_s_3_300=1.18e-11
+  mcm4d_ca_w_0_300_s_9_000=8.37e-06 mcm4d_cc_w_0_300_s_9_000=8.66e-12 mcm4d_cf_w_0_300_s_9_000=2.23e-11
+  mcm4d_ca_w_2_400_s_0_300=8.37e-06 mcm4d_cc_w_2_400_s_0_300=1.24e-10 mcm4d_cf_w_2_400_s_0_300=1.40e-12
+  mcm4d_ca_w_2_400_s_0_360=8.37e-06 mcm4d_cc_w_2_400_s_0_360=1.17e-10 mcm4d_cf_w_2_400_s_0_360=1.64e-12
+  mcm4d_ca_w_2_400_s_0_450=8.37e-06 mcm4d_cc_w_2_400_s_0_450=1.08e-10 mcm4d_cf_w_2_400_s_0_450=2.01e-12
+  mcm4d_ca_w_2_400_s_0_600=8.37e-06 mcm4d_cc_w_2_400_s_0_600=9.53e-11 mcm4d_cf_w_2_400_s_0_600=2.61e-12
+  mcm4d_ca_w_2_400_s_0_800=8.37e-06 mcm4d_cc_w_2_400_s_0_800=8.23e-11 mcm4d_cf_w_2_400_s_0_800=3.41e-12
+  mcm4d_ca_w_2_400_s_1_000=8.37e-06 mcm4d_cc_w_2_400_s_1_000=7.27e-11 mcm4d_cf_w_2_400_s_1_000=4.18e-12
+  mcm4d_ca_w_2_400_s_1_200=8.37e-06 mcm4d_cc_w_2_400_s_1_200=6.52e-11 mcm4d_cf_w_2_400_s_1_200=4.94e-12
+  mcm4d_ca_w_2_400_s_2_100=8.37e-06 mcm4d_cc_w_2_400_s_2_100=4.59e-11 mcm4d_cf_w_2_400_s_2_100=8.21e-12
+  mcm4d_ca_w_2_400_s_3_300=8.37e-06 mcm4d_cc_w_2_400_s_3_300=3.34e-11 mcm4d_cf_w_2_400_s_3_300=1.21e-11
+  mcm4d_ca_w_2_400_s_9_000=8.37e-06 mcm4d_cc_w_2_400_s_9_000=1.27e-11 mcm4d_cf_w_2_400_s_9_000=2.44e-11
+  mcm4p1_ca_w_0_300_s_0_300=8.88e-06 mcm4p1_cc_w_0_300_s_0_300=9.63e-11 mcm4p1_cf_w_0_300_s_0_300=1.46e-12
+  mcm4p1_ca_w_0_300_s_0_360=8.88e-06 mcm4p1_cc_w_0_300_s_0_360=9.07e-11 mcm4p1_cf_w_0_300_s_0_360=1.73e-12
+  mcm4p1_ca_w_0_300_s_0_450=8.88e-06 mcm4p1_cc_w_0_300_s_0_450=8.28e-11 mcm4p1_cf_w_0_300_s_0_450=2.13e-12
+  mcm4p1_ca_w_0_300_s_0_600=8.88e-06 mcm4p1_cc_w_0_300_s_0_600=7.25e-11 mcm4p1_cf_w_0_300_s_0_600=2.80e-12
+  mcm4p1_ca_w_0_300_s_0_800=8.88e-06 mcm4p1_cc_w_0_300_s_0_800=6.24e-11 mcm4p1_cf_w_0_300_s_0_800=3.58e-12
+  mcm4p1_ca_w_0_300_s_1_000=8.88e-06 mcm4p1_cc_w_0_300_s_1_000=5.45e-11 mcm4p1_cf_w_0_300_s_1_000=4.38e-12
+  mcm4p1_ca_w_0_300_s_1_200=8.88e-06 mcm4p1_cc_w_0_300_s_1_200=4.86e-11 mcm4p1_cf_w_0_300_s_1_200=5.18e-12
+  mcm4p1_ca_w_0_300_s_2_100=8.88e-06 mcm4p1_cc_w_0_300_s_2_100=3.36e-11 mcm4p1_cf_w_0_300_s_2_100=8.79e-12
+  mcm4p1_ca_w_0_300_s_3_300=8.88e-06 mcm4p1_cc_w_0_300_s_3_300=2.42e-11 mcm4p1_cf_w_0_300_s_3_300=1.24e-11
+  mcm4p1_ca_w_0_300_s_9_000=8.88e-06 mcm4p1_cc_w_0_300_s_9_000=8.28e-12 mcm4p1_cf_w_0_300_s_9_000=2.31e-11
+  mcm4p1_ca_w_2_400_s_0_300=8.88e-06 mcm4p1_cc_w_2_400_s_0_300=1.24e-10 mcm4p1_cf_w_2_400_s_0_300=1.50e-12
+  mcm4p1_ca_w_2_400_s_0_360=8.88e-06 mcm4p1_cc_w_2_400_s_0_360=1.17e-10 mcm4p1_cf_w_2_400_s_0_360=1.76e-12
+  mcm4p1_ca_w_2_400_s_0_450=8.88e-06 mcm4p1_cc_w_2_400_s_0_450=1.07e-10 mcm4p1_cf_w_2_400_s_0_450=2.14e-12
+  mcm4p1_ca_w_2_400_s_0_600=8.88e-06 mcm4p1_cc_w_2_400_s_0_600=9.47e-11 mcm4p1_cf_w_2_400_s_0_600=2.78e-12
+  mcm4p1_ca_w_2_400_s_0_800=8.88e-06 mcm4p1_cc_w_2_400_s_0_800=8.18e-11 mcm4p1_cf_w_2_400_s_0_800=3.62e-12
+  mcm4p1_ca_w_2_400_s_1_000=8.88e-06 mcm4p1_cc_w_2_400_s_1_000=7.21e-11 mcm4p1_cf_w_2_400_s_1_000=4.44e-12
+  mcm4p1_ca_w_2_400_s_1_200=8.88e-06 mcm4p1_cc_w_2_400_s_1_200=6.46e-11 mcm4p1_cf_w_2_400_s_1_200=5.25e-12
+  mcm4p1_ca_w_2_400_s_2_100=8.88e-06 mcm4p1_cc_w_2_400_s_2_100=4.53e-11 mcm4p1_cf_w_2_400_s_2_100=8.69e-12
+  mcm4p1_ca_w_2_400_s_3_300=8.88e-06 mcm4p1_cc_w_2_400_s_3_300=3.28e-11 mcm4p1_cf_w_2_400_s_3_300=1.28e-11
+  mcm4p1_ca_w_2_400_s_9_000=8.88e-06 mcm4p1_cc_w_2_400_s_9_000=1.22e-11 mcm4p1_cf_w_2_400_s_9_000=2.53e-11
+  mcm4l1_ca_w_0_300_s_0_300=1.04e-05 mcm4l1_cc_w_0_300_s_0_300=9.60e-11 mcm4l1_cf_w_0_300_s_0_300=1.71e-12
+  mcm4l1_ca_w_0_300_s_0_360=1.04e-05 mcm4l1_cc_w_0_300_s_0_360=9.02e-11 mcm4l1_cf_w_0_300_s_0_360=2.01e-12
+  mcm4l1_ca_w_0_300_s_0_450=1.04e-05 mcm4l1_cc_w_0_300_s_0_450=8.23e-11 mcm4l1_cf_w_0_300_s_0_450=2.49e-12
+  mcm4l1_ca_w_0_300_s_0_600=1.04e-05 mcm4l1_cc_w_0_300_s_0_600=7.19e-11 mcm4l1_cf_w_0_300_s_0_600=3.26e-12
+  mcm4l1_ca_w_0_300_s_0_800=1.04e-05 mcm4l1_cc_w_0_300_s_0_800=6.18e-11 mcm4l1_cf_w_0_300_s_0_800=4.16e-12
+  mcm4l1_ca_w_0_300_s_1_000=1.04e-05 mcm4l1_cc_w_0_300_s_1_000=5.38e-11 mcm4l1_cf_w_0_300_s_1_000=5.09e-12
+  mcm4l1_ca_w_0_300_s_1_200=1.04e-05 mcm4l1_cc_w_0_300_s_1_200=4.79e-11 mcm4l1_cf_w_0_300_s_1_200=6.01e-12
+  mcm4l1_ca_w_0_300_s_2_100=1.04e-05 mcm4l1_cc_w_0_300_s_2_100=3.25e-11 mcm4l1_cf_w_0_300_s_2_100=1.01e-11
+  mcm4l1_ca_w_0_300_s_3_300=1.04e-05 mcm4l1_cc_w_0_300_s_3_300=2.30e-11 mcm4l1_cf_w_0_300_s_3_300=1.41e-11
+  mcm4l1_ca_w_0_300_s_9_000=1.04e-05 mcm4l1_cc_w_0_300_s_9_000=7.31e-12 mcm4l1_cf_w_0_300_s_9_000=2.53e-11
+  mcm4l1_ca_w_2_400_s_0_300=1.04e-05 mcm4l1_cc_w_2_400_s_0_300=1.23e-10 mcm4l1_cf_w_2_400_s_0_300=1.73e-12
+  mcm4l1_ca_w_2_400_s_0_360=1.04e-05 mcm4l1_cc_w_2_400_s_0_360=1.16e-10 mcm4l1_cf_w_2_400_s_0_360=2.03e-12
+  mcm4l1_ca_w_2_400_s_0_450=1.04e-05 mcm4l1_cc_w_2_400_s_0_450=1.06e-10 mcm4l1_cf_w_2_400_s_0_450=2.48e-12
+  mcm4l1_ca_w_2_400_s_0_600=1.04e-05 mcm4l1_cc_w_2_400_s_0_600=9.33e-11 mcm4l1_cf_w_2_400_s_0_600=3.22e-12
+  mcm4l1_ca_w_2_400_s_0_800=1.04e-05 mcm4l1_cc_w_2_400_s_0_800=8.04e-11 mcm4l1_cf_w_2_400_s_0_800=4.20e-12
+  mcm4l1_ca_w_2_400_s_1_000=1.04e-05 mcm4l1_cc_w_2_400_s_1_000=7.06e-11 mcm4l1_cf_w_2_400_s_1_000=5.15e-12
+  mcm4l1_ca_w_2_400_s_1_200=1.04e-05 mcm4l1_cc_w_2_400_s_1_200=6.31e-11 mcm4l1_cf_w_2_400_s_1_200=6.08e-12
+  mcm4l1_ca_w_2_400_s_2_100=1.04e-05 mcm4l1_cc_w_2_400_s_2_100=4.38e-11 mcm4l1_cf_w_2_400_s_2_100=1.00e-11
+  mcm4l1_ca_w_2_400_s_3_300=1.04e-05 mcm4l1_cc_w_2_400_s_3_300=3.12e-11 mcm4l1_cf_w_2_400_s_3_300=1.46e-11
+  mcm4l1_ca_w_2_400_s_9_000=1.04e-05 mcm4l1_cc_w_2_400_s_9_000=1.10e-11 mcm4l1_cf_w_2_400_s_9_000=2.78e-11
+  mcm4m1_ca_w_0_300_s_0_300=1.34e-05 mcm4m1_cc_w_0_300_s_0_300=9.52e-11 mcm4m1_cf_w_0_300_s_0_300=2.18e-12
+  mcm4m1_ca_w_0_300_s_0_360=1.34e-05 mcm4m1_cc_w_0_300_s_0_360=8.93e-11 mcm4m1_cf_w_0_300_s_0_360=2.57e-12
+  mcm4m1_ca_w_0_300_s_0_450=1.34e-05 mcm4m1_cc_w_0_300_s_0_450=8.14e-11 mcm4m1_cf_w_0_300_s_0_450=3.17e-12
+  mcm4m1_ca_w_0_300_s_0_600=1.34e-05 mcm4m1_cc_w_0_300_s_0_600=7.09e-11 mcm4m1_cf_w_0_300_s_0_600=4.14e-12
+  mcm4m1_ca_w_0_300_s_0_800=1.34e-05 mcm4m1_cc_w_0_300_s_0_800=6.05e-11 mcm4m1_cf_w_0_300_s_0_800=5.28e-12
+  mcm4m1_ca_w_0_300_s_1_000=1.34e-05 mcm4m1_cc_w_0_300_s_1_000=5.25e-11 mcm4m1_cf_w_0_300_s_1_000=6.44e-12
+  mcm4m1_ca_w_0_300_s_1_200=1.34e-05 mcm4m1_cc_w_0_300_s_1_200=4.64e-11 mcm4m1_cf_w_0_300_s_1_200=7.57e-12
+  mcm4m1_ca_w_0_300_s_2_100=1.34e-05 mcm4m1_cc_w_0_300_s_2_100=3.06e-11 mcm4m1_cf_w_0_300_s_2_100=1.25e-11
+  mcm4m1_ca_w_0_300_s_3_300=1.34e-05 mcm4m1_cc_w_0_300_s_3_300=2.10e-11 mcm4m1_cf_w_0_300_s_3_300=1.72e-11
+  mcm4m1_ca_w_0_300_s_9_000=1.34e-05 mcm4m1_cc_w_0_300_s_9_000=5.93e-12 mcm4m1_cf_w_0_300_s_9_000=2.87e-11
+  mcm4m1_ca_w_2_400_s_0_300=1.34e-05 mcm4m1_cc_w_2_400_s_0_300=1.20e-10 mcm4m1_cf_w_2_400_s_0_300=2.19e-12
+  mcm4m1_ca_w_2_400_s_0_360=1.34e-05 mcm4m1_cc_w_2_400_s_0_360=1.13e-10 mcm4m1_cf_w_2_400_s_0_360=2.58e-12
+  mcm4m1_ca_w_2_400_s_0_450=1.34e-05 mcm4m1_cc_w_2_400_s_0_450=1.04e-10 mcm4m1_cf_w_2_400_s_0_450=3.16e-12
+  mcm4m1_ca_w_2_400_s_0_600=1.34e-05 mcm4m1_cc_w_2_400_s_0_600=9.09e-11 mcm4m1_cf_w_2_400_s_0_600=4.09e-12
+  mcm4m1_ca_w_2_400_s_0_800=1.34e-05 mcm4m1_cc_w_2_400_s_0_800=7.80e-11 mcm4m1_cf_w_2_400_s_0_800=5.32e-12
+  mcm4m1_ca_w_2_400_s_1_000=1.34e-05 mcm4m1_cc_w_2_400_s_1_000=6.82e-11 mcm4m1_cf_w_2_400_s_1_000=6.51e-12
+  mcm4m1_ca_w_2_400_s_1_200=1.34e-05 mcm4m1_cc_w_2_400_s_1_200=6.07e-11 mcm4m1_cf_w_2_400_s_1_200=7.66e-12
+  mcm4m1_ca_w_2_400_s_2_100=1.34e-05 mcm4m1_cc_w_2_400_s_2_100=4.13e-11 mcm4m1_cf_w_2_400_s_2_100=1.24e-11
+  mcm4m1_ca_w_2_400_s_3_300=1.34e-05 mcm4m1_cc_w_2_400_s_3_300=2.88e-11 mcm4m1_cf_w_2_400_s_3_300=1.78e-11
+  mcm4m1_ca_w_2_400_s_9_000=1.34e-05 mcm4m1_cc_w_2_400_s_9_000=9.34e-12 mcm4m1_cf_w_2_400_s_9_000=3.17e-11
+  mcm4m2_ca_w_0_300_s_0_300=1.86e-05 mcm4m2_cc_w_0_300_s_0_300=9.39e-11 mcm4m2_cf_w_0_300_s_0_300=3.01e-12
+  mcm4m2_ca_w_0_300_s_0_360=1.86e-05 mcm4m2_cc_w_0_300_s_0_360=8.80e-11 mcm4m2_cf_w_0_300_s_0_360=3.54e-12
+  mcm4m2_ca_w_0_300_s_0_450=1.86e-05 mcm4m2_cc_w_0_300_s_0_450=8.00e-11 mcm4m2_cf_w_0_300_s_0_450=4.34e-12
+  mcm4m2_ca_w_0_300_s_0_600=1.86e-05 mcm4m2_cc_w_0_300_s_0_600=6.92e-11 mcm4m2_cf_w_0_300_s_0_600=5.64e-12
+  mcm4m2_ca_w_0_300_s_0_800=1.86e-05 mcm4m2_cc_w_0_300_s_0_800=5.86e-11 mcm4m2_cf_w_0_300_s_0_800=7.19e-12
+  mcm4m2_ca_w_0_300_s_1_000=1.86e-05 mcm4m2_cc_w_0_300_s_1_000=5.04e-11 mcm4m2_cf_w_0_300_s_1_000=8.72e-12
+  mcm4m2_ca_w_0_300_s_1_200=1.86e-05 mcm4m2_cc_w_0_300_s_1_200=4.41e-11 mcm4m2_cf_w_0_300_s_1_200=1.02e-11
+  mcm4m2_ca_w_0_300_s_2_100=1.86e-05 mcm4m2_cc_w_0_300_s_2_100=2.79e-11 mcm4m2_cf_w_0_300_s_2_100=1.64e-11
+  mcm4m2_ca_w_0_300_s_3_300=1.86e-05 mcm4m2_cc_w_0_300_s_3_300=1.83e-11 mcm4m2_cf_w_0_300_s_3_300=2.19e-11
+  mcm4m2_ca_w_0_300_s_9_000=1.86e-05 mcm4m2_cc_w_0_300_s_9_000=4.55e-12 mcm4m2_cf_w_0_300_s_9_000=3.32e-11
+  mcm4m2_ca_w_2_400_s_0_300=1.86e-05 mcm4m2_cc_w_2_400_s_0_300=1.17e-10 mcm4m2_cf_w_2_400_s_0_300=3.02e-12
+  mcm4m2_ca_w_2_400_s_0_360=1.86e-05 mcm4m2_cc_w_2_400_s_0_360=1.10e-10 mcm4m2_cf_w_2_400_s_0_360=3.55e-12
+  mcm4m2_ca_w_2_400_s_0_450=1.86e-05 mcm4m2_cc_w_2_400_s_0_450=1.01e-10 mcm4m2_cf_w_2_400_s_0_450=4.33e-12
+  mcm4m2_ca_w_2_400_s_0_600=1.86e-05 mcm4m2_cc_w_2_400_s_0_600=8.76e-11 mcm4m2_cf_w_2_400_s_0_600=5.60e-12
+  mcm4m2_ca_w_2_400_s_0_800=1.86e-05 mcm4m2_cc_w_2_400_s_0_800=7.46e-11 mcm4m2_cf_w_2_400_s_0_800=7.24e-12
+  mcm4m2_ca_w_2_400_s_1_000=1.86e-05 mcm4m2_cc_w_2_400_s_1_000=6.48e-11 mcm4m2_cf_w_2_400_s_1_000=8.82e-12
+  mcm4m2_ca_w_2_400_s_1_200=1.86e-05 mcm4m2_cc_w_2_400_s_1_200=5.73e-11 mcm4m2_cf_w_2_400_s_1_200=1.03e-11
+  mcm4m2_ca_w_2_400_s_2_100=1.86e-05 mcm4m2_cc_w_2_400_s_2_100=3.80e-11 mcm4m2_cf_w_2_400_s_2_100=1.64e-11
+  mcm4m2_ca_w_2_400_s_3_300=1.86e-05 mcm4m2_cc_w_2_400_s_3_300=2.57e-11 mcm4m2_cf_w_2_400_s_3_300=2.27e-11
+  mcm4m2_ca_w_2_400_s_9_000=1.86e-05 mcm4m2_cc_w_2_400_s_9_000=7.55e-12 mcm4m2_cf_w_2_400_s_9_000=3.69e-11
+  mcm4m3_ca_w_0_300_s_0_300=6.43e-05 mcm4m3_cc_w_0_300_s_0_300=8.52e-11 mcm4m3_cf_w_0_300_s_0_300=9.76e-12
+  mcm4m3_ca_w_0_300_s_0_360=6.43e-05 mcm4m3_cc_w_0_300_s_0_360=7.90e-11 mcm4m3_cf_w_0_300_s_0_360=1.13e-11
+  mcm4m3_ca_w_0_300_s_0_450=6.43e-05 mcm4m3_cc_w_0_300_s_0_450=7.05e-11 mcm4m3_cf_w_0_300_s_0_450=1.36e-11
+  mcm4m3_ca_w_0_300_s_0_600=6.43e-05 mcm4m3_cc_w_0_300_s_0_600=5.91e-11 mcm4m3_cf_w_0_300_s_0_600=1.70e-11
+  mcm4m3_ca_w_0_300_s_0_800=6.43e-05 mcm4m3_cc_w_0_300_s_0_800=4.82e-11 mcm4m3_cf_w_0_300_s_0_800=2.10e-11
+  mcm4m3_ca_w_0_300_s_1_000=6.43e-05 mcm4m3_cc_w_0_300_s_1_000=3.99e-11 mcm4m3_cf_w_0_300_s_1_000=2.45e-11
+  mcm4m3_ca_w_0_300_s_1_200=6.43e-05 mcm4m3_cc_w_0_300_s_1_200=3.36e-11 mcm4m3_cf_w_0_300_s_1_200=2.76e-11
+  mcm4m3_ca_w_0_300_s_2_100=6.43e-05 mcm4m3_cc_w_0_300_s_2_100=1.79e-11 mcm4m3_cf_w_0_300_s_2_100=3.79e-11
+  mcm4m3_ca_w_0_300_s_3_300=6.43e-05 mcm4m3_cc_w_0_300_s_3_300=1.01e-11 mcm4m3_cf_w_0_300_s_3_300=4.43e-11
+  mcm4m3_ca_w_0_300_s_9_000=6.43e-05 mcm4m3_cc_w_0_300_s_9_000=1.95e-12 mcm4m3_cf_w_0_300_s_9_000=5.21e-11
+  mcm4m3_ca_w_2_400_s_0_300=6.43e-05 mcm4m3_cc_w_2_400_s_0_300=1.04e-10 mcm4m3_cf_w_2_400_s_0_300=9.78e-12
+  mcm4m3_ca_w_2_400_s_0_360=6.43e-05 mcm4m3_cc_w_2_400_s_0_360=9.66e-11 mcm4m3_cf_w_2_400_s_0_360=1.13e-11
+  mcm4m3_ca_w_2_400_s_0_450=6.43e-05 mcm4m3_cc_w_2_400_s_0_450=8.71e-11 mcm4m3_cf_w_2_400_s_0_450=1.36e-11
+  mcm4m3_ca_w_2_400_s_0_600=6.43e-05 mcm4m3_cc_w_2_400_s_0_600=7.44e-11 mcm4m3_cf_w_2_400_s_0_600=1.70e-11
+  mcm4m3_ca_w_2_400_s_0_800=6.43e-05 mcm4m3_cc_w_2_400_s_0_800=6.17e-11 mcm4m3_cf_w_2_400_s_0_800=2.11e-11
+  mcm4m3_ca_w_2_400_s_1_000=6.43e-05 mcm4m3_cc_w_2_400_s_1_000=5.23e-11 mcm4m3_cf_w_2_400_s_1_000=2.46e-11
+  mcm4m3_ca_w_2_400_s_1_200=6.43e-05 mcm4m3_cc_w_2_400_s_1_200=4.51e-11 mcm4m3_cf_w_2_400_s_1_200=2.78e-11
+  mcm4m3_ca_w_2_400_s_2_100=6.43e-05 mcm4m3_cc_w_2_400_s_2_100=2.74e-11 mcm4m3_cf_w_2_400_s_2_100=3.80e-11
+  mcm4m3_ca_w_2_400_s_3_300=6.43e-05 mcm4m3_cc_w_2_400_s_3_300=1.68e-11 mcm4m3_cf_w_2_400_s_3_300=4.62e-11
+  mcm4m3_ca_w_2_400_s_9_000=6.43e-05 mcm4m3_cc_w_2_400_s_9_000=4.10e-12 mcm4m3_cf_w_2_400_s_9_000=5.80e-11
+  mcm5f_ca_w_1_600_s_1_600=5.81e-06 mcm5f_cc_w_1_600_s_1_600=6.73e-11 mcm5f_cf_w_1_600_s_1_600=4.71e-12
+  mcm5f_ca_w_1_600_s_1_700=5.81e-06 mcm5f_cc_w_1_600_s_1_700=6.42e-11 mcm5f_cf_w_1_600_s_1_700=4.98e-12
+  mcm5f_ca_w_1_600_s_1_900=5.81e-06 mcm5f_cc_w_1_600_s_1_900=5.91e-11 mcm5f_cf_w_1_600_s_1_900=5.51e-12
+  mcm5f_ca_w_1_600_s_2_000=5.81e-06 mcm5f_cc_w_1_600_s_2_000=5.69e-11 mcm5f_cf_w_1_600_s_2_000=5.77e-12
+  mcm5f_ca_w_1_600_s_2_400=5.81e-06 mcm5f_cc_w_1_600_s_2_400=4.97e-11 mcm5f_cf_w_1_600_s_2_400=6.81e-12
+  mcm5f_ca_w_1_600_s_2_800=5.81e-06 mcm5f_cc_w_1_600_s_2_800=4.43e-11 mcm5f_cf_w_1_600_s_2_800=7.81e-12
+  mcm5f_ca_w_1_600_s_3_200=5.81e-06 mcm5f_cc_w_1_600_s_3_200=4.00e-11 mcm5f_cf_w_1_600_s_3_200=8.79e-12
+  mcm5f_ca_w_1_600_s_4_800=5.81e-06 mcm5f_cc_w_1_600_s_4_800=2.90e-11 mcm5f_cf_w_1_600_s_4_800=1.24e-11
+  mcm5f_ca_w_1_600_s_10_000=5.81e-06 mcm5f_cc_w_1_600_s_10_000=1.42e-11 mcm5f_cf_w_1_600_s_10_000=2.09e-11
+  mcm5f_ca_w_1_600_s_12_000=5.81e-06 mcm5f_cc_w_1_600_s_12_000=1.14e-11 mcm5f_cf_w_1_600_s_12_000=2.31e-11
+  mcm5f_ca_w_4_000_s_1_600=5.81e-06 mcm5f_cc_w_4_000_s_1_600=7.46e-11 mcm5f_cf_w_4_000_s_1_600=4.71e-12
+  mcm5f_ca_w_4_000_s_1_700=5.81e-06 mcm5f_cc_w_4_000_s_1_700=7.13e-11 mcm5f_cf_w_4_000_s_1_700=4.98e-12
+  mcm5f_ca_w_4_000_s_1_900=5.81e-06 mcm5f_cc_w_4_000_s_1_900=6.58e-11 mcm5f_cf_w_4_000_s_1_900=5.51e-12
+  mcm5f_ca_w_4_000_s_2_000=5.81e-06 mcm5f_cc_w_4_000_s_2_000=6.35e-11 mcm5f_cf_w_4_000_s_2_000=5.78e-12
+  mcm5f_ca_w_4_000_s_2_400=5.81e-06 mcm5f_cc_w_4_000_s_2_400=5.58e-11 mcm5f_cf_w_4_000_s_2_400=6.82e-12
+  mcm5f_ca_w_4_000_s_2_800=5.81e-06 mcm5f_cc_w_4_000_s_2_800=4.99e-11 mcm5f_cf_w_4_000_s_2_800=7.83e-12
+  mcm5f_ca_w_4_000_s_3_200=5.81e-06 mcm5f_cc_w_4_000_s_3_200=4.52e-11 mcm5f_cf_w_4_000_s_3_200=8.82e-12
+  mcm5f_ca_w_4_000_s_4_800=5.81e-06 mcm5f_cc_w_4_000_s_4_800=3.32e-11 mcm5f_cf_w_4_000_s_4_800=1.25e-11
+  mcm5f_ca_w_4_000_s_10_000=5.81e-06 mcm5f_cc_w_4_000_s_10_000=1.69e-11 mcm5f_cf_w_4_000_s_10_000=2.13e-11
+  mcm5f_ca_w_4_000_s_12_000=5.81e-06 mcm5f_cc_w_4_000_s_12_000=1.38e-11 mcm5f_cf_w_4_000_s_12_000=2.37e-11
+  mcm5d_ca_w_1_600_s_1_600=6.21e-06 mcm5d_cc_w_1_600_s_1_600=6.68e-11 mcm5d_cf_w_1_600_s_1_600=5.02e-12
+  mcm5d_ca_w_1_600_s_1_700=6.21e-06 mcm5d_cc_w_1_600_s_1_700=6.38e-11 mcm5d_cf_w_1_600_s_1_700=5.31e-12
+  mcm5d_ca_w_1_600_s_1_900=6.21e-06 mcm5d_cc_w_1_600_s_1_900=5.86e-11 mcm5d_cf_w_1_600_s_1_900=5.87e-12
+  mcm5d_ca_w_1_600_s_2_000=6.21e-06 mcm5d_cc_w_1_600_s_2_000=5.64e-11 mcm5d_cf_w_1_600_s_2_000=6.15e-12
+  mcm5d_ca_w_1_600_s_2_400=6.21e-06 mcm5d_cc_w_1_600_s_2_400=4.92e-11 mcm5d_cf_w_1_600_s_2_400=7.25e-12
+  mcm5d_ca_w_1_600_s_2_800=6.21e-06 mcm5d_cc_w_1_600_s_2_800=4.38e-11 mcm5d_cf_w_1_600_s_2_800=8.31e-12
+  mcm5d_ca_w_1_600_s_3_200=6.21e-06 mcm5d_cc_w_1_600_s_3_200=3.95e-11 mcm5d_cf_w_1_600_s_3_200=9.34e-12
+  mcm5d_ca_w_1_600_s_4_800=6.21e-06 mcm5d_cc_w_1_600_s_4_800=2.84e-11 mcm5d_cf_w_1_600_s_4_800=1.31e-11
+  mcm5d_ca_w_1_600_s_10_000=6.21e-06 mcm5d_cc_w_1_600_s_10_000=1.36e-11 mcm5d_cf_w_1_600_s_10_000=2.19e-11
+  mcm5d_ca_w_1_600_s_12_000=6.21e-06 mcm5d_cc_w_1_600_s_12_000=1.09e-11 mcm5d_cf_w_1_600_s_12_000=2.41e-11
+  mcm5d_ca_w_4_000_s_1_600=6.21e-06 mcm5d_cc_w_4_000_s_1_600=7.41e-11 mcm5d_cf_w_4_000_s_1_600=5.03e-12
+  mcm5d_ca_w_4_000_s_1_700=6.21e-06 mcm5d_cc_w_4_000_s_1_700=7.07e-11 mcm5d_cf_w_4_000_s_1_700=5.31e-12
+  mcm5d_ca_w_4_000_s_1_900=6.21e-06 mcm5d_cc_w_4_000_s_1_900=6.51e-11 mcm5d_cf_w_4_000_s_1_900=5.88e-12
+  mcm5d_ca_w_4_000_s_2_000=6.21e-06 mcm5d_cc_w_4_000_s_2_000=6.28e-11 mcm5d_cf_w_4_000_s_2_000=6.16e-12
+  mcm5d_ca_w_4_000_s_2_400=6.21e-06 mcm5d_cc_w_4_000_s_2_400=5.51e-11 mcm5d_cf_w_4_000_s_2_400=7.26e-12
+  mcm5d_ca_w_4_000_s_2_800=6.21e-06 mcm5d_cc_w_4_000_s_2_800=4.93e-11 mcm5d_cf_w_4_000_s_2_800=8.34e-12
+  mcm5d_ca_w_4_000_s_3_200=6.21e-06 mcm5d_cc_w_4_000_s_3_200=4.46e-11 mcm5d_cf_w_4_000_s_3_200=9.37e-12
+  mcm5d_ca_w_4_000_s_4_800=6.21e-06 mcm5d_cc_w_4_000_s_4_800=3.26e-11 mcm5d_cf_w_4_000_s_4_800=1.32e-11
+  mcm5d_ca_w_4_000_s_10_000=6.21e-06 mcm5d_cc_w_4_000_s_10_000=1.63e-11 mcm5d_cf_w_4_000_s_10_000=2.23e-11
+  mcm5d_ca_w_4_000_s_12_000=6.21e-06 mcm5d_cc_w_4_000_s_12_000=1.33e-11 mcm5d_cf_w_4_000_s_12_000=2.47e-11
+  mcm5p1_ca_w_1_600_s_1_600=6.49e-06 mcm5p1_cc_w_1_600_s_1_600=6.65e-11 mcm5p1_cf_w_1_600_s_1_600=5.25e-12
+  mcm5p1_ca_w_1_600_s_1_700=6.49e-06 mcm5p1_cc_w_1_600_s_1_700=6.35e-11 mcm5p1_cf_w_1_600_s_1_700=5.54e-12
+  mcm5p1_ca_w_1_600_s_1_900=6.49e-06 mcm5p1_cc_w_1_600_s_1_900=5.82e-11 mcm5p1_cf_w_1_600_s_1_900=6.13e-12
+  mcm5p1_ca_w_1_600_s_2_000=6.49e-06 mcm5p1_cc_w_1_600_s_2_000=5.61e-11 mcm5p1_cf_w_1_600_s_2_000=6.42e-12
+  mcm5p1_ca_w_1_600_s_2_400=6.49e-06 mcm5p1_cc_w_1_600_s_2_400=4.88e-11 mcm5p1_cf_w_1_600_s_2_400=7.56e-12
+  mcm5p1_ca_w_1_600_s_2_800=6.49e-06 mcm5p1_cc_w_1_600_s_2_800=4.34e-11 mcm5p1_cf_w_1_600_s_2_800=8.67e-12
+  mcm5p1_ca_w_1_600_s_3_200=6.49e-06 mcm5p1_cc_w_1_600_s_3_200=3.91e-11 mcm5p1_cf_w_1_600_s_3_200=9.73e-12
+  mcm5p1_ca_w_1_600_s_4_800=6.49e-06 mcm5p1_cc_w_1_600_s_4_800=2.80e-11 mcm5p1_cf_w_1_600_s_4_800=1.36e-11
+  mcm5p1_ca_w_1_600_s_10_000=6.49e-06 mcm5p1_cc_w_1_600_s_10_000=1.33e-11 mcm5p1_cf_w_1_600_s_10_000=2.25e-11
+  mcm5p1_ca_w_1_600_s_12_000=6.49e-06 mcm5p1_cc_w_1_600_s_12_000=1.05e-11 mcm5p1_cf_w_1_600_s_12_000=2.47e-11
+  mcm5p1_ca_w_4_000_s_1_600=6.49e-06 mcm5p1_cc_w_4_000_s_1_600=7.37e-11 mcm5p1_cf_w_4_000_s_1_600=5.25e-12
+  mcm5p1_ca_w_4_000_s_1_700=6.49e-06 mcm5p1_cc_w_4_000_s_1_700=7.03e-11 mcm5p1_cf_w_4_000_s_1_700=5.55e-12
+  mcm5p1_ca_w_4_000_s_1_900=6.49e-06 mcm5p1_cc_w_4_000_s_1_900=6.47e-11 mcm5p1_cf_w_4_000_s_1_900=6.14e-12
+  mcm5p1_ca_w_4_000_s_2_000=6.49e-06 mcm5p1_cc_w_4_000_s_2_000=6.24e-11 mcm5p1_cf_w_4_000_s_2_000=6.43e-12
+  mcm5p1_ca_w_4_000_s_2_400=6.49e-06 mcm5p1_cc_w_4_000_s_2_400=5.46e-11 mcm5p1_cf_w_4_000_s_2_400=7.58e-12
+  mcm5p1_ca_w_4_000_s_2_800=6.49e-06 mcm5p1_cc_w_4_000_s_2_800=4.88e-11 mcm5p1_cf_w_4_000_s_2_800=8.69e-12
+  mcm5p1_ca_w_4_000_s_3_200=6.49e-06 mcm5p1_cc_w_4_000_s_3_200=4.42e-11 mcm5p1_cf_w_4_000_s_3_200=9.77e-12
+  mcm5p1_ca_w_4_000_s_4_800=6.49e-06 mcm5p1_cc_w_4_000_s_4_800=3.21e-11 mcm5p1_cf_w_4_000_s_4_800=1.37e-11
+  mcm5p1_ca_w_4_000_s_10_000=6.49e-06 mcm5p1_cc_w_4_000_s_10_000=1.59e-11 mcm5p1_cf_w_4_000_s_10_000=2.30e-11
+  mcm5p1_ca_w_4_000_s_12_000=6.49e-06 mcm5p1_cc_w_4_000_s_12_000=1.29e-11 mcm5p1_cf_w_4_000_s_12_000=2.54e-11
+  mcm5l1_ca_w_1_600_s_1_600=7.27e-06 mcm5l1_cc_w_1_600_s_1_600=6.57e-11 mcm5l1_cf_w_1_600_s_1_600=5.84e-12
+  mcm5l1_ca_w_1_600_s_1_700=7.27e-06 mcm5l1_cc_w_1_600_s_1_700=6.27e-11 mcm5l1_cf_w_1_600_s_1_700=6.17e-12
+  mcm5l1_ca_w_1_600_s_1_900=7.27e-06 mcm5l1_cc_w_1_600_s_1_900=5.74e-11 mcm5l1_cf_w_1_600_s_1_900=6.81e-12
+  mcm5l1_ca_w_1_600_s_2_000=7.27e-06 mcm5l1_cc_w_1_600_s_2_000=5.52e-11 mcm5l1_cf_w_1_600_s_2_000=7.14e-12
+  mcm5l1_ca_w_1_600_s_2_400=7.27e-06 mcm5l1_cc_w_1_600_s_2_400=4.79e-11 mcm5l1_cf_w_1_600_s_2_400=8.40e-12
+  mcm5l1_ca_w_1_600_s_2_800=7.27e-06 mcm5l1_cc_w_1_600_s_2_800=4.24e-11 mcm5l1_cf_w_1_600_s_2_800=9.61e-12
+  mcm5l1_ca_w_1_600_s_3_200=7.27e-06 mcm5l1_cc_w_1_600_s_3_200=3.81e-11 mcm5l1_cf_w_1_600_s_3_200=1.08e-11
+  mcm5l1_ca_w_1_600_s_4_800=7.27e-06 mcm5l1_cc_w_1_600_s_4_800=2.70e-11 mcm5l1_cf_w_1_600_s_4_800=1.50e-11
+  mcm5l1_ca_w_1_600_s_10_000=7.27e-06 mcm5l1_cc_w_1_600_s_10_000=1.24e-11 mcm5l1_cf_w_1_600_s_10_000=2.43e-11
+  mcm5l1_ca_w_1_600_s_12_000=7.27e-06 mcm5l1_cc_w_1_600_s_12_000=9.73e-12 mcm5l1_cf_w_1_600_s_12_000=2.65e-11
+  mcm5l1_ca_w_4_000_s_1_600=7.27e-06 mcm5l1_cc_w_4_000_s_1_600=7.25e-11 mcm5l1_cf_w_4_000_s_1_600=5.84e-12
+  mcm5l1_ca_w_4_000_s_1_700=7.27e-06 mcm5l1_cc_w_4_000_s_1_700=6.92e-11 mcm5l1_cf_w_4_000_s_1_700=6.18e-12
+  mcm5l1_ca_w_4_000_s_1_900=7.27e-06 mcm5l1_cc_w_4_000_s_1_900=6.36e-11 mcm5l1_cf_w_4_000_s_1_900=6.82e-12
+  mcm5l1_ca_w_4_000_s_2_000=7.27e-06 mcm5l1_cc_w_4_000_s_2_000=6.13e-11 mcm5l1_cf_w_4_000_s_2_000=7.14e-12
+  mcm5l1_ca_w_4_000_s_2_400=7.27e-06 mcm5l1_cc_w_4_000_s_2_400=5.35e-11 mcm5l1_cf_w_4_000_s_2_400=8.41e-12
+  mcm5l1_ca_w_4_000_s_2_800=7.27e-06 mcm5l1_cc_w_4_000_s_2_800=4.76e-11 mcm5l1_cf_w_4_000_s_2_800=9.63e-12
+  mcm5l1_ca_w_4_000_s_3_200=7.27e-06 mcm5l1_cc_w_4_000_s_3_200=4.30e-11 mcm5l1_cf_w_4_000_s_3_200=1.08e-11
+  mcm5l1_ca_w_4_000_s_4_800=7.27e-06 mcm5l1_cc_w_4_000_s_4_800=3.10e-11 mcm5l1_cf_w_4_000_s_4_800=1.51e-11
+  mcm5l1_ca_w_4_000_s_10_000=7.27e-06 mcm5l1_cc_w_4_000_s_10_000=1.50e-11 mcm5l1_cf_w_4_000_s_10_000=2.48e-11
+  mcm5l1_ca_w_4_000_s_12_000=7.27e-06 mcm5l1_cc_w_4_000_s_12_000=1.20e-11 mcm5l1_cf_w_4_000_s_12_000=2.72e-11
+  mcm5m1_ca_w_1_600_s_1_600=8.59e-06 mcm5m1_cc_w_1_600_s_1_600=6.44e-11 mcm5m1_cf_w_1_600_s_1_600=6.85e-12
+  mcm5m1_ca_w_1_600_s_1_700=8.59e-06 mcm5m1_cc_w_1_600_s_1_700=6.13e-11 mcm5m1_cf_w_1_600_s_1_700=7.22e-12
+  mcm5m1_ca_w_1_600_s_1_900=8.59e-06 mcm5m1_cc_w_1_600_s_1_900=5.60e-11 mcm5m1_cf_w_1_600_s_1_900=7.97e-12
+  mcm5m1_ca_w_1_600_s_2_000=8.59e-06 mcm5m1_cc_w_1_600_s_2_000=5.39e-11 mcm5m1_cf_w_1_600_s_2_000=8.35e-12
+  mcm5m1_ca_w_1_600_s_2_400=8.59e-06 mcm5m1_cc_w_1_600_s_2_400=4.65e-11 mcm5m1_cf_w_1_600_s_2_400=9.80e-12
+  mcm5m1_ca_w_1_600_s_2_800=8.59e-06 mcm5m1_cc_w_1_600_s_2_800=4.10e-11 mcm5m1_cf_w_1_600_s_2_800=1.12e-11
+  mcm5m1_ca_w_1_600_s_3_200=8.59e-06 mcm5m1_cc_w_1_600_s_3_200=3.66e-11 mcm5m1_cf_w_1_600_s_3_200=1.25e-11
+  mcm5m1_ca_w_1_600_s_4_800=8.59e-06 mcm5m1_cc_w_1_600_s_4_800=2.55e-11 mcm5m1_cf_w_1_600_s_4_800=1.72e-11
+  mcm5m1_ca_w_1_600_s_10_000=8.59e-06 mcm5m1_cc_w_1_600_s_10_000=1.11e-11 mcm5m1_cf_w_1_600_s_10_000=2.70e-11
+  mcm5m1_ca_w_1_600_s_12_000=8.59e-06 mcm5m1_cc_w_1_600_s_12_000=8.62e-12 mcm5m1_cf_w_1_600_s_12_000=2.91e-11
+  mcm5m1_ca_w_4_000_s_1_600=8.59e-06 mcm5m1_cc_w_4_000_s_1_600=7.08e-11 mcm5m1_cf_w_4_000_s_1_600=6.85e-12
+  mcm5m1_ca_w_4_000_s_1_700=8.59e-06 mcm5m1_cc_w_4_000_s_1_700=6.75e-11 mcm5m1_cf_w_4_000_s_1_700=7.23e-12
+  mcm5m1_ca_w_4_000_s_1_900=8.59e-06 mcm5m1_cc_w_4_000_s_1_900=6.20e-11 mcm5m1_cf_w_4_000_s_1_900=7.99e-12
+  mcm5m1_ca_w_4_000_s_2_000=8.59e-06 mcm5m1_cc_w_4_000_s_2_000=5.96e-11 mcm5m1_cf_w_4_000_s_2_000=8.36e-12
+  mcm5m1_ca_w_4_000_s_2_400=8.59e-06 mcm5m1_cc_w_4_000_s_2_400=5.18e-11 mcm5m1_cf_w_4_000_s_2_400=9.82e-12
+  mcm5m1_ca_w_4_000_s_2_800=8.59e-06 mcm5m1_cc_w_4_000_s_2_800=4.59e-11 mcm5m1_cf_w_4_000_s_2_800=1.12e-11
+  mcm5m1_ca_w_4_000_s_3_200=8.59e-06 mcm5m1_cc_w_4_000_s_3_200=4.13e-11 mcm5m1_cf_w_4_000_s_3_200=1.26e-11
+  mcm5m1_ca_w_4_000_s_4_800=8.59e-06 mcm5m1_cc_w_4_000_s_4_800=2.93e-11 mcm5m1_cf_w_4_000_s_4_800=1.73e-11
+  mcm5m1_ca_w_4_000_s_10_000=8.59e-06 mcm5m1_cc_w_4_000_s_10_000=1.36e-11 mcm5m1_cf_w_4_000_s_10_000=2.76e-11
+  mcm5m1_ca_w_4_000_s_12_000=8.59e-06 mcm5m1_cc_w_4_000_s_12_000=1.08e-11 mcm5m1_cf_w_4_000_s_12_000=2.99e-11
+  mcm5m2_ca_w_1_600_s_1_600=1.05e-05 mcm5m2_cc_w_1_600_s_1_600=6.26e-11 mcm5m2_cf_w_1_600_s_1_600=8.24e-12
+  mcm5m2_ca_w_1_600_s_1_700=1.05e-05 mcm5m2_cc_w_1_600_s_1_700=5.96e-11 mcm5m2_cf_w_1_600_s_1_700=8.70e-12
+  mcm5m2_ca_w_1_600_s_1_900=1.05e-05 mcm5m2_cc_w_1_600_s_1_900=5.43e-11 mcm5m2_cf_w_1_600_s_1_900=9.59e-12
+  mcm5m2_ca_w_1_600_s_2_000=1.05e-05 mcm5m2_cc_w_1_600_s_2_000=5.21e-11 mcm5m2_cf_w_1_600_s_2_000=1.00e-11
+  mcm5m2_ca_w_1_600_s_2_400=1.05e-05 mcm5m2_cc_w_1_600_s_2_400=4.47e-11 mcm5m2_cf_w_1_600_s_2_400=1.17e-11
+  mcm5m2_ca_w_1_600_s_2_800=1.05e-05 mcm5m2_cc_w_1_600_s_2_800=3.91e-11 mcm5m2_cf_w_1_600_s_2_800=1.33e-11
+  mcm5m2_ca_w_1_600_s_3_200=1.05e-05 mcm5m2_cc_w_1_600_s_3_200=3.48e-11 mcm5m2_cf_w_1_600_s_3_200=1.49e-11
+  mcm5m2_ca_w_1_600_s_4_800=1.05e-05 mcm5m2_cc_w_1_600_s_4_800=2.36e-11 mcm5m2_cf_w_1_600_s_4_800=2.02e-11
+  mcm5m2_ca_w_1_600_s_10_000=1.05e-05 mcm5m2_cc_w_1_600_s_10_000=9.73e-12 mcm5m2_cf_w_1_600_s_10_000=3.02e-11
+  mcm5m2_ca_w_1_600_s_12_000=1.05e-05 mcm5m2_cc_w_1_600_s_12_000=7.46e-12 mcm5m2_cf_w_1_600_s_12_000=3.23e-11
+  mcm5m2_ca_w_4_000_s_1_600=1.05e-05 mcm5m2_cc_w_4_000_s_1_600=6.88e-11 mcm5m2_cf_w_4_000_s_1_600=8.25e-12
+  mcm5m2_ca_w_4_000_s_1_700=1.05e-05 mcm5m2_cc_w_4_000_s_1_700=6.55e-11 mcm5m2_cf_w_4_000_s_1_700=8.71e-12
+  mcm5m2_ca_w_4_000_s_1_900=1.05e-05 mcm5m2_cc_w_4_000_s_1_900=5.99e-11 mcm5m2_cf_w_4_000_s_1_900=9.60e-12
+  mcm5m2_ca_w_4_000_s_2_000=1.05e-05 mcm5m2_cc_w_4_000_s_2_000=5.75e-11 mcm5m2_cf_w_4_000_s_2_000=1.00e-11
+  mcm5m2_ca_w_4_000_s_2_400=1.05e-05 mcm5m2_cc_w_4_000_s_2_400=4.97e-11 mcm5m2_cf_w_4_000_s_2_400=1.17e-11
+  mcm5m2_ca_w_4_000_s_2_800=1.05e-05 mcm5m2_cc_w_4_000_s_2_800=4.39e-11 mcm5m2_cf_w_4_000_s_2_800=1.34e-11
+  mcm5m2_ca_w_4_000_s_3_200=1.05e-05 mcm5m2_cc_w_4_000_s_3_200=3.92e-11 mcm5m2_cf_w_4_000_s_3_200=1.49e-11
+  mcm5m2_ca_w_4_000_s_4_800=1.05e-05 mcm5m2_cc_w_4_000_s_4_800=2.73e-11 mcm5m2_cf_w_4_000_s_4_800=2.03e-11
+  mcm5m2_ca_w_4_000_s_10_000=1.05e-05 mcm5m2_cc_w_4_000_s_10_000=1.22e-11 mcm5m2_cf_w_4_000_s_10_000=3.09e-11
+  mcm5m2_ca_w_4_000_s_12_000=1.05e-05 mcm5m2_cc_w_4_000_s_12_000=9.55e-12 mcm5m2_cf_w_4_000_s_12_000=3.32e-11
+  mcm5m3_ca_w_1_600_s_1_600=1.75e-05 mcm5m3_cc_w_1_600_s_1_600=5.77e-11 mcm5m3_cf_w_1_600_s_1_600=1.32e-11
+  mcm5m3_ca_w_1_600_s_1_700=1.75e-05 mcm5m3_cc_w_1_600_s_1_700=5.45e-11 mcm5m3_cf_w_1_600_s_1_700=1.39e-11
+  mcm5m3_ca_w_1_600_s_1_900=1.75e-05 mcm5m3_cc_w_1_600_s_1_900=4.93e-11 mcm5m3_cf_w_1_600_s_1_900=1.52e-11
+  mcm5m3_ca_w_1_600_s_2_000=1.75e-05 mcm5m3_cc_w_1_600_s_2_000=4.71e-11 mcm5m3_cf_w_1_600_s_2_000=1.58e-11
+  mcm5m3_ca_w_1_600_s_2_400=1.75e-05 mcm5m3_cc_w_1_600_s_2_400=3.96e-11 mcm5m3_cf_w_1_600_s_2_400=1.83e-11
+  mcm5m3_ca_w_1_600_s_2_800=1.75e-05 mcm5m3_cc_w_1_600_s_2_800=3.41e-11 mcm5m3_cf_w_1_600_s_2_800=2.06e-11
+  mcm5m3_ca_w_1_600_s_3_200=1.75e-05 mcm5m3_cc_w_1_600_s_3_200=2.99e-11 mcm5m3_cf_w_1_600_s_3_200=2.26e-11
+  mcm5m3_ca_w_1_600_s_4_800=1.75e-05 mcm5m3_cc_w_1_600_s_4_800=1.90e-11 mcm5m3_cf_w_1_600_s_4_800=2.92e-11
+  mcm5m3_ca_w_1_600_s_10_000=1.75e-05 mcm5m3_cc_w_1_600_s_10_000=6.90e-12 mcm5m3_cf_w_1_600_s_10_000=3.93e-11
+  mcm5m3_ca_w_1_600_s_12_000=1.75e-05 mcm5m3_cc_w_1_600_s_12_000=5.25e-12 mcm5m3_cf_w_1_600_s_12_000=4.09e-11
+  mcm5m3_ca_w_4_000_s_1_600=1.75e-05 mcm5m3_cc_w_4_000_s_1_600=6.32e-11 mcm5m3_cf_w_4_000_s_1_600=1.32e-11
+  mcm5m3_ca_w_4_000_s_1_700=1.75e-05 mcm5m3_cc_w_4_000_s_1_700=6.00e-11 mcm5m3_cf_w_4_000_s_1_700=1.39e-11
+  mcm5m3_ca_w_4_000_s_1_900=1.75e-05 mcm5m3_cc_w_4_000_s_1_900=5.44e-11 mcm5m3_cf_w_4_000_s_1_900=1.52e-11
+  mcm5m3_ca_w_4_000_s_2_000=1.75e-05 mcm5m3_cc_w_4_000_s_2_000=5.21e-11 mcm5m3_cf_w_4_000_s_2_000=1.58e-11
+  mcm5m3_ca_w_4_000_s_2_400=1.75e-05 mcm5m3_cc_w_4_000_s_2_400=4.43e-11 mcm5m3_cf_w_4_000_s_2_400=1.83e-11
+  mcm5m3_ca_w_4_000_s_2_800=1.75e-05 mcm5m3_cc_w_4_000_s_2_800=3.85e-11 mcm5m3_cf_w_4_000_s_2_800=2.06e-11
+  mcm5m3_ca_w_4_000_s_3_200=1.75e-05 mcm5m3_cc_w_4_000_s_3_200=3.40e-11 mcm5m3_cf_w_4_000_s_3_200=2.27e-11
+  mcm5m3_ca_w_4_000_s_4_800=1.75e-05 mcm5m3_cc_w_4_000_s_4_800=2.26e-11 mcm5m3_cf_w_4_000_s_4_800=2.94e-11
+  mcm5m3_ca_w_4_000_s_10_000=1.75e-05 mcm5m3_cc_w_4_000_s_10_000=9.25e-12 mcm5m3_cf_w_4_000_s_10_000=4.02e-11
+  mcm5m3_ca_w_4_000_s_12_000=1.75e-05 mcm5m3_cc_w_4_000_s_12_000=7.15e-12 mcm5m3_cf_w_4_000_s_12_000=4.21e-11
+  mcm5m4_ca_w_1_600_s_1_600=5.30e-05 mcm5m4_cc_w_1_600_s_1_600=4.63e-11 mcm5m4_cf_w_1_600_s_1_600=3.26e-11
+  mcm5m4_ca_w_1_600_s_1_700=5.30e-05 mcm5m4_cc_w_1_600_s_1_700=4.32e-11 mcm5m4_cf_w_1_600_s_1_700=3.38e-11
+  mcm5m4_ca_w_1_600_s_1_900=5.30e-05 mcm5m4_cc_w_1_600_s_1_900=3.82e-11 mcm5m4_cf_w_1_600_s_1_900=3.62e-11
+  mcm5m4_ca_w_1_600_s_2_000=5.30e-05 mcm5m4_cc_w_1_600_s_2_000=3.61e-11 mcm5m4_cf_w_1_600_s_2_000=3.73e-11
+  mcm5m4_ca_w_1_600_s_2_400=5.30e-05 mcm5m4_cc_w_1_600_s_2_400=2.92e-11 mcm5m4_cf_w_1_600_s_2_400=4.12e-11
+  mcm5m4_ca_w_1_600_s_2_800=5.30e-05 mcm5m4_cc_w_1_600_s_2_800=2.42e-11 mcm5m4_cf_w_1_600_s_2_800=4.45e-11
+  mcm5m4_ca_w_1_600_s_3_200=5.30e-05 mcm5m4_cc_w_1_600_s_3_200=2.05e-11 mcm5m4_cf_w_1_600_s_3_200=4.71e-11
+  mcm5m4_ca_w_1_600_s_4_800=5.30e-05 mcm5m4_cc_w_1_600_s_4_800=1.20e-11 mcm5m4_cf_w_1_600_s_4_800=5.41e-11
+  mcm5m4_ca_w_1_600_s_10_000=5.30e-05 mcm5m4_cc_w_1_600_s_10_000=4.00e-12 mcm5m4_cf_w_1_600_s_10_000=6.16e-11
+  mcm5m4_ca_w_1_600_s_12_000=5.30e-05 mcm5m4_cc_w_1_600_s_12_000=3.00e-12 mcm5m4_cf_w_1_600_s_12_000=6.26e-11
+  mcm5m4_ca_w_4_000_s_1_600=5.30e-05 mcm5m4_cc_w_4_000_s_1_600=5.16e-11 mcm5m4_cf_w_4_000_s_1_600=3.26e-11
+  mcm5m4_ca_w_4_000_s_1_700=5.30e-05 mcm5m4_cc_w_4_000_s_1_700=4.85e-11 mcm5m4_cf_w_4_000_s_1_700=3.38e-11
+  mcm5m4_ca_w_4_000_s_1_900=5.30e-05 mcm5m4_cc_w_4_000_s_1_900=4.33e-11 mcm5m4_cf_w_4_000_s_1_900=3.63e-11
+  mcm5m4_ca_w_4_000_s_2_000=5.30e-05 mcm5m4_cc_w_4_000_s_2_000=4.11e-11 mcm5m4_cf_w_4_000_s_2_000=3.73e-11
+  mcm5m4_ca_w_4_000_s_2_400=5.30e-05 mcm5m4_cc_w_4_000_s_2_400=3.39e-11 mcm5m4_cf_w_4_000_s_2_400=4.13e-11
+  mcm5m4_ca_w_4_000_s_2_800=5.30e-05 mcm5m4_cc_w_4_000_s_2_800=2.88e-11 mcm5m4_cf_w_4_000_s_2_800=4.45e-11
+  mcm5m4_ca_w_4_000_s_3_200=5.30e-05 mcm5m4_cc_w_4_000_s_3_200=2.48e-11 mcm5m4_cf_w_4_000_s_3_200=4.72e-11
+  mcm5m4_ca_w_4_000_s_4_800=5.30e-05 mcm5m4_cc_w_4_000_s_4_800=1.56e-11 mcm5m4_cf_w_4_000_s_4_800=5.45e-11
+  mcm5m4_ca_w_4_000_s_10_000=5.30e-05 mcm5m4_cc_w_4_000_s_10_000=6.05e-12 mcm5m4_cf_w_4_000_s_10_000=6.33e-11
+  mcm5m4_ca_w_4_000_s_12_000=5.30e-05 mcm5m4_cc_w_4_000_s_12_000=4.65e-12 mcm5m4_cf_w_4_000_s_12_000=6.47e-11
+  mcrdlf_ca_w_10_000_s_5_000=2.26e-06 mcrdlf_cc_w_10_000_s_5_000=4.39e-11 mcrdlf_cf_w_10_000_s_5_000=5.98e-12
+  mcrdlf_ca_w_10_000_s_8_000=2.26e-06 mcrdlf_cc_w_10_000_s_8_000=3.32e-11 mcrdlf_cf_w_10_000_s_8_000=8.69e-12
+  mcrdlf_ca_w_10_000_s_10_000=2.26e-06 mcrdlf_cc_w_10_000_s_10_000=2.88e-11 mcrdlf_cf_w_10_000_s_10_000=1.03e-11
+  mcrdlf_ca_w_10_000_s_12_000=2.26e-06 mcrdlf_cc_w_10_000_s_12_000=2.54e-11 mcrdlf_cf_w_10_000_s_12_000=1.18e-11
+  mcrdlf_ca_w_10_000_s_30_000=2.26e-06 mcrdlf_cc_w_10_000_s_30_000=1.15e-11 mcrdlf_cf_w_10_000_s_30_000=2.11e-11
+  mcrdlf_ca_w_40_000_s_5_000=2.26e-06 mcrdlf_cc_w_40_000_s_5_000=5.53e-11 mcrdlf_cf_w_40_000_s_5_000=6.06e-12
+  mcrdlf_ca_w_40_000_s_8_000=2.26e-06 mcrdlf_cc_w_40_000_s_8_000=4.36e-11 mcrdlf_cf_w_40_000_s_8_000=8.77e-12
+  mcrdlf_ca_w_40_000_s_10_000=2.26e-06 mcrdlf_cc_w_40_000_s_10_000=3.86e-11 mcrdlf_cf_w_40_000_s_10_000=1.04e-11
+  mcrdlf_ca_w_40_000_s_12_000=2.26e-06 mcrdlf_cc_w_40_000_s_12_000=3.48e-11 mcrdlf_cf_w_40_000_s_12_000=1.20e-11
+  mcrdlf_ca_w_40_000_s_30_000=2.26e-06 mcrdlf_cc_w_40_000_s_30_000=1.87e-11 mcrdlf_cf_w_40_000_s_30_000=2.19e-11
+  mcrdld_ca_w_10_000_s_5_000=2.32e-06 mcrdld_cc_w_10_000_s_5_000=4.37e-11 mcrdld_cf_w_10_000_s_5_000=6.12e-12
+  mcrdld_ca_w_10_000_s_8_000=2.32e-06 mcrdld_cc_w_10_000_s_8_000=3.30e-11 mcrdld_cf_w_10_000_s_8_000=8.88e-12
+  mcrdld_ca_w_10_000_s_10_000=2.32e-06 mcrdld_cc_w_10_000_s_10_000=2.85e-11 mcrdld_cf_w_10_000_s_10_000=1.06e-11
+  mcrdld_ca_w_10_000_s_12_000=2.32e-06 mcrdld_cc_w_10_000_s_12_000=2.52e-11 mcrdld_cf_w_10_000_s_12_000=1.21e-11
+  mcrdld_ca_w_10_000_s_30_000=2.32e-06 mcrdld_cc_w_10_000_s_30_000=1.14e-11 mcrdld_cf_w_10_000_s_30_000=2.14e-11
+  mcrdld_ca_w_40_000_s_5_000=2.32e-06 mcrdld_cc_w_40_000_s_5_000=5.50e-11 mcrdld_cf_w_40_000_s_5_000=6.21e-12
+  mcrdld_ca_w_40_000_s_8_000=2.32e-06 mcrdld_cc_w_40_000_s_8_000=4.34e-11 mcrdld_cf_w_40_000_s_8_000=8.98e-12
+  mcrdld_ca_w_40_000_s_10_000=2.32e-06 mcrdld_cc_w_40_000_s_10_000=3.84e-11 mcrdld_cf_w_40_000_s_10_000=1.07e-11
+  mcrdld_ca_w_40_000_s_12_000=2.32e-06 mcrdld_cc_w_40_000_s_12_000=3.47e-11 mcrdld_cf_w_40_000_s_12_000=1.22e-11
+  mcrdld_ca_w_40_000_s_30_000=2.32e-06 mcrdld_cc_w_40_000_s_30_000=1.86e-11 mcrdld_cf_w_40_000_s_30_000=2.22e-11
+  mcrdlp1_ca_w_10_000_s_5_000=2.36e-06 mcrdlp1_cc_w_10_000_s_5_000=4.36e-11 mcrdlp1_cf_w_10_000_s_5_000=6.21e-12
+  mcrdlp1_ca_w_10_000_s_8_000=2.36e-06 mcrdlp1_cc_w_10_000_s_8_000=3.28e-11 mcrdlp1_cf_w_10_000_s_8_000=9.00e-12
+  mcrdlp1_ca_w_10_000_s_10_000=2.36e-06 mcrdlp1_cc_w_10_000_s_10_000=2.84e-11 mcrdlp1_cf_w_10_000_s_10_000=1.07e-11
+  mcrdlp1_ca_w_10_000_s_12_000=2.36e-06 mcrdlp1_cc_w_10_000_s_12_000=2.51e-11 mcrdlp1_cf_w_10_000_s_12_000=1.22e-11
+  mcrdlp1_ca_w_10_000_s_30_000=2.36e-06 mcrdlp1_cc_w_10_000_s_30_000=1.13e-11 mcrdlp1_cf_w_10_000_s_30_000=2.16e-11
+  mcrdlp1_ca_w_40_000_s_5_000=2.36e-06 mcrdlp1_cc_w_40_000_s_5_000=5.49e-11 mcrdlp1_cf_w_40_000_s_5_000=6.31e-12
+  mcrdlp1_ca_w_40_000_s_8_000=2.36e-06 mcrdlp1_cc_w_40_000_s_8_000=4.33e-11 mcrdlp1_cf_w_40_000_s_8_000=9.12e-12
+  mcrdlp1_ca_w_40_000_s_10_000=2.36e-06 mcrdlp1_cc_w_40_000_s_10_000=3.83e-11 mcrdlp1_cf_w_40_000_s_10_000=1.08e-11
+  mcrdlp1_ca_w_40_000_s_12_000=2.36e-06 mcrdlp1_cc_w_40_000_s_12_000=3.45e-11 mcrdlp1_cf_w_40_000_s_12_000=1.24e-11
+  mcrdlp1_ca_w_40_000_s_30_000=2.36e-06 mcrdlp1_cc_w_40_000_s_30_000=1.84e-11 mcrdlp1_cf_w_40_000_s_30_000=2.24e-11
+  mcrdll1_ca_w_10_000_s_5_000=2.45e-06 mcrdll1_cc_w_10_000_s_5_000=4.32e-11 mcrdll1_cf_w_10_000_s_5_000=6.43e-12
+  mcrdll1_ca_w_10_000_s_8_000=2.45e-06 mcrdll1_cc_w_10_000_s_8_000=3.25e-11 mcrdll1_cf_w_10_000_s_8_000=9.31e-12
+  mcrdll1_ca_w_10_000_s_10_000=2.45e-06 mcrdll1_cc_w_10_000_s_10_000=2.81e-11 mcrdll1_cf_w_10_000_s_10_000=1.10e-11
+  mcrdll1_ca_w_10_000_s_12_000=2.45e-06 mcrdll1_cc_w_10_000_s_12_000=2.47e-11 mcrdll1_cf_w_10_000_s_12_000=1.26e-11
+  mcrdll1_ca_w_10_000_s_30_000=2.45e-06 mcrdll1_cc_w_10_000_s_30_000=1.10e-11 mcrdll1_cf_w_10_000_s_30_000=2.20e-11
+  mcrdll1_ca_w_40_000_s_5_000=2.45e-06 mcrdll1_cc_w_40_000_s_5_000=5.45e-11 mcrdll1_cf_w_40_000_s_5_000=6.53e-12
+  mcrdll1_ca_w_40_000_s_8_000=2.45e-06 mcrdll1_cc_w_40_000_s_8_000=4.28e-11 mcrdll1_cf_w_40_000_s_8_000=9.41e-12
+  mcrdll1_ca_w_40_000_s_10_000=2.45e-06 mcrdll1_cc_w_40_000_s_10_000=3.79e-11 mcrdll1_cf_w_40_000_s_10_000=1.12e-11
+  mcrdll1_ca_w_40_000_s_12_000=2.45e-06 mcrdll1_cc_w_40_000_s_12_000=3.42e-11 mcrdll1_cf_w_40_000_s_12_000=1.28e-11
+  mcrdll1_ca_w_40_000_s_30_000=2.45e-06 mcrdll1_cc_w_40_000_s_30_000=1.82e-11 mcrdll1_cf_w_40_000_s_30_000=2.29e-11
+  mcrdlm1_ca_w_10_000_s_5_000=2.58e-06 mcrdlm1_cc_w_10_000_s_5_000=4.28e-11 mcrdlm1_cf_w_10_000_s_5_000=6.75e-12
+  mcrdlm1_ca_w_10_000_s_8_000=2.58e-06 mcrdlm1_cc_w_10_000_s_8_000=3.21e-11 mcrdlm1_cf_w_10_000_s_8_000=9.74e-12
+  mcrdlm1_ca_w_10_000_s_10_000=2.58e-06 mcrdlm1_cc_w_10_000_s_10_000=2.77e-11 mcrdlm1_cf_w_10_000_s_10_000=1.15e-11
+  mcrdlm1_ca_w_10_000_s_12_000=2.58e-06 mcrdlm1_cc_w_10_000_s_12_000=2.43e-11 mcrdlm1_cf_w_10_000_s_12_000=1.32e-11
+  mcrdlm1_ca_w_10_000_s_30_000=2.58e-06 mcrdlm1_cc_w_10_000_s_30_000=1.07e-11 mcrdlm1_cf_w_10_000_s_30_000=2.27e-11
+  mcrdlm1_ca_w_40_000_s_5_000=2.58e-06 mcrdlm1_cc_w_40_000_s_5_000=5.40e-11 mcrdlm1_cf_w_40_000_s_5_000=6.83e-12
+  mcrdlm1_ca_w_40_000_s_8_000=2.58e-06 mcrdlm1_cc_w_40_000_s_8_000=4.24e-11 mcrdlm1_cf_w_40_000_s_8_000=9.84e-12
+  mcrdlm1_ca_w_40_000_s_10_000=2.58e-06 mcrdlm1_cc_w_40_000_s_10_000=3.74e-11 mcrdlm1_cf_w_40_000_s_10_000=1.16e-11
+  mcrdlm1_ca_w_40_000_s_12_000=2.58e-06 mcrdlm1_cc_w_40_000_s_12_000=3.37e-11 mcrdlm1_cf_w_40_000_s_12_000=1.33e-11
+  mcrdlm1_ca_w_40_000_s_30_000=2.58e-06 mcrdlm1_cc_w_40_000_s_30_000=1.78e-11 mcrdlm1_cf_w_40_000_s_30_000=2.36e-11
+  mcrdlm2_ca_w_10_000_s_5_000=2.73e-06 mcrdlm2_cc_w_10_000_s_5_000=4.24e-11 mcrdlm2_cf_w_10_000_s_5_000=7.09e-12
+  mcrdlm2_ca_w_10_000_s_8_000=2.73e-06 mcrdlm2_cc_w_10_000_s_8_000=3.16e-11 mcrdlm2_cf_w_10_000_s_8_000=1.02e-11
+  mcrdlm2_ca_w_10_000_s_10_000=2.73e-06 mcrdlm2_cc_w_10_000_s_10_000=2.72e-11 mcrdlm2_cf_w_10_000_s_10_000=1.21e-11
+  mcrdlm2_ca_w_10_000_s_12_000=2.73e-06 mcrdlm2_cc_w_10_000_s_12_000=2.38e-11 mcrdlm2_cf_w_10_000_s_12_000=1.37e-11
+  mcrdlm2_ca_w_10_000_s_30_000=2.73e-06 mcrdlm2_cc_w_10_000_s_30_000=1.04e-11 mcrdlm2_cf_w_10_000_s_30_000=2.34e-11
+  mcrdlm2_ca_w_40_000_s_5_000=2.73e-06 mcrdlm2_cc_w_40_000_s_5_000=5.35e-11 mcrdlm2_cf_w_40_000_s_5_000=7.18e-12
+  mcrdlm2_ca_w_40_000_s_8_000=2.73e-06 mcrdlm2_cc_w_40_000_s_8_000=4.19e-11 mcrdlm2_cf_w_40_000_s_8_000=1.03e-11
+  mcrdlm2_ca_w_40_000_s_10_000=2.73e-06 mcrdlm2_cc_w_40_000_s_10_000=3.70e-11 mcrdlm2_cf_w_40_000_s_10_000=1.22e-11
+  mcrdlm2_ca_w_40_000_s_12_000=2.73e-06 mcrdlm2_cc_w_40_000_s_12_000=3.33e-11 mcrdlm2_cf_w_40_000_s_12_000=1.39e-11
+  mcrdlm2_ca_w_40_000_s_30_000=2.73e-06 mcrdlm2_cc_w_40_000_s_30_000=1.75e-11 mcrdlm2_cf_w_40_000_s_30_000=2.43e-11
+  mcrdlm3_ca_w_10_000_s_5_000=3.06e-06 mcrdlm3_cc_w_10_000_s_5_000=4.14e-11 mcrdlm3_cf_w_10_000_s_5_000=7.78e-12
+  mcrdlm3_ca_w_10_000_s_8_000=3.06e-06 mcrdlm3_cc_w_10_000_s_8_000=3.07e-11 mcrdlm3_cf_w_10_000_s_8_000=1.11e-11
+  mcrdlm3_ca_w_10_000_s_10_000=3.06e-06 mcrdlm3_cc_w_10_000_s_10_000=2.63e-11 mcrdlm3_cf_w_10_000_s_10_000=1.31e-11
+  mcrdlm3_ca_w_10_000_s_12_000=3.06e-06 mcrdlm3_cc_w_10_000_s_12_000=2.30e-11 mcrdlm3_cf_w_10_000_s_12_000=1.49e-11
+  mcrdlm3_ca_w_10_000_s_30_000=3.06e-06 mcrdlm3_cc_w_10_000_s_30_000=9.75e-12 mcrdlm3_cf_w_10_000_s_30_000=2.47e-11
+  mcrdlm3_ca_w_40_000_s_5_000=3.06e-06 mcrdlm3_cc_w_40_000_s_5_000=5.26e-11 mcrdlm3_cf_w_40_000_s_5_000=7.72e-12
+  mcrdlm3_ca_w_40_000_s_8_000=3.06e-06 mcrdlm3_cc_w_40_000_s_8_000=4.10e-11 mcrdlm3_cf_w_40_000_s_8_000=1.11e-11
+  mcrdlm3_ca_w_40_000_s_10_000=3.06e-06 mcrdlm3_cc_w_40_000_s_10_000=3.61e-11 mcrdlm3_cf_w_40_000_s_10_000=1.31e-11
+  mcrdlm3_ca_w_40_000_s_12_000=3.06e-06 mcrdlm3_cc_w_40_000_s_12_000=3.24e-11 mcrdlm3_cf_w_40_000_s_12_000=1.49e-11
+  mcrdlm3_ca_w_40_000_s_30_000=3.06e-06 mcrdlm3_cc_w_40_000_s_30_000=1.69e-11 mcrdlm3_cf_w_40_000_s_30_000=2.56e-11
+  mcrdlm4_ca_w_10_000_s_5_000=3.47e-06 mcrdlm4_cc_w_10_000_s_5_000=4.04e-11 mcrdlm4_cf_w_10_000_s_5_000=8.67e-12
+  mcrdlm4_ca_w_10_000_s_8_000=3.47e-06 mcrdlm4_cc_w_10_000_s_8_000=2.98e-11 mcrdlm4_cf_w_10_000_s_8_000=1.23e-11
+  mcrdlm4_ca_w_10_000_s_10_000=3.47e-06 mcrdlm4_cc_w_10_000_s_10_000=2.53e-11 mcrdlm4_cf_w_10_000_s_10_000=1.44e-11
+  mcrdlm4_ca_w_10_000_s_12_000=3.47e-06 mcrdlm4_cc_w_10_000_s_12_000=2.21e-11 mcrdlm4_cf_w_10_000_s_12_000=1.63e-11
+  mcrdlm4_ca_w_10_000_s_30_000=3.47e-06 mcrdlm4_cc_w_10_000_s_30_000=9.11e-12 mcrdlm4_cf_w_10_000_s_30_000=2.62e-11
+  mcrdlm4_ca_w_40_000_s_5_000=3.47e-06 mcrdlm4_cc_w_40_000_s_5_000=5.15e-11 mcrdlm4_cf_w_40_000_s_5_000=8.56e-12
+  mcrdlm4_ca_w_40_000_s_8_000=3.47e-06 mcrdlm4_cc_w_40_000_s_8_000=4.00e-11 mcrdlm4_cf_w_40_000_s_8_000=1.22e-11
+  mcrdlm4_ca_w_40_000_s_10_000=3.47e-06 mcrdlm4_cc_w_40_000_s_10_000=3.52e-11 mcrdlm4_cf_w_40_000_s_10_000=1.44e-11
+  mcrdlm4_ca_w_40_000_s_12_000=3.47e-06 mcrdlm4_cc_w_40_000_s_12_000=3.14e-11 mcrdlm4_cf_w_40_000_s_12_000=1.63e-11
+  mcrdlm4_ca_w_40_000_s_30_000=3.47e-06 mcrdlm4_cc_w_40_000_s_30_000=1.62e-11 mcrdlm4_cf_w_40_000_s_30_000=2.72e-11
+  mcrdlm5_ca_w_10_000_s_5_000=4.58e-06 mcrdlm5_cc_w_10_000_s_5_000=3.83e-11 mcrdlm5_cf_w_10_000_s_5_000=1.10e-11
+  mcrdlm5_ca_w_10_000_s_8_000=4.58e-06 mcrdlm5_cc_w_10_000_s_8_000=2.77e-11 mcrdlm5_cf_w_10_000_s_8_000=1.53e-11
+  mcrdlm5_ca_w_10_000_s_10_000=4.58e-06 mcrdlm5_cc_w_10_000_s_10_000=2.34e-11 mcrdlm5_cf_w_10_000_s_10_000=1.77e-11
+  mcrdlm5_ca_w_10_000_s_12_000=4.58e-06 mcrdlm5_cc_w_10_000_s_12_000=2.02e-11 mcrdlm5_cf_w_10_000_s_12_000=1.98e-11
+  mcrdlm5_ca_w_10_000_s_30_000=4.58e-06 mcrdlm5_cc_w_10_000_s_30_000=8.00e-12 mcrdlm5_cf_w_10_000_s_30_000=2.97e-11
+  mcrdlm5_ca_w_40_000_s_5_000=4.58e-06 mcrdlm5_cc_w_40_000_s_5_000=4.94e-11 mcrdlm5_cf_w_40_000_s_5_000=1.09e-11
+  mcrdlm5_ca_w_40_000_s_8_000=4.58e-06 mcrdlm5_cc_w_40_000_s_8_000=3.80e-11 mcrdlm5_cf_w_40_000_s_8_000=1.52e-11
+  mcrdlm5_ca_w_40_000_s_10_000=4.58e-06 mcrdlm5_cc_w_40_000_s_10_000=3.32e-11 mcrdlm5_cf_w_40_000_s_10_000=1.77e-11
+  mcrdlm5_ca_w_40_000_s_12_000=4.58e-06 mcrdlm5_cc_w_40_000_s_12_000=2.96e-11 mcrdlm5_cf_w_40_000_s_12_000=1.98e-11
+  mcrdlm5_ca_w_40_000_s_30_000=4.58e-06 mcrdlm5_cc_w_40_000_s_30_000=1.50e-11 mcrdlm5_cf_w_40_000_s_30_000=3.11e-11
+  mcl1p1f_ca_w_0_150_s_0_210=1.58e-04 mcl1p1f_cc_w_0_150_s_0_210=5.88e-11 mcl1p1f_cf_w_0_150_s_0_210=1.62e-11
+  mcl1p1f_ca_w_0_150_s_0_263=1.58e-04 mcl1p1f_cc_w_0_150_s_0_263=4.66e-11 mcl1p1f_cf_w_0_150_s_0_263=1.95e-11
+  mcl1p1f_ca_w_0_150_s_0_315=1.58e-04 mcl1p1f_cc_w_0_150_s_0_315=3.78e-11 mcl1p1f_cf_w_0_150_s_0_315=2.26e-11
+  mcl1p1f_ca_w_0_150_s_0_420=1.58e-04 mcl1p1f_cc_w_0_150_s_0_420=2.64e-11 mcl1p1f_cf_w_0_150_s_0_420=2.80e-11
+  mcl1p1f_ca_w_0_150_s_0_525=1.58e-04 mcl1p1f_cc_w_0_150_s_0_525=1.89e-11 mcl1p1f_cf_w_0_150_s_0_525=3.24e-11
+  mcl1p1f_ca_w_0_150_s_0_630=1.58e-04 mcl1p1f_cc_w_0_150_s_0_630=1.37e-11 mcl1p1f_cf_w_0_150_s_0_630=3.59e-11
+  mcl1p1f_ca_w_0_150_s_0_840=1.58e-04 mcl1p1f_cc_w_0_150_s_0_840=7.42e-12 mcl1p1f_cf_w_0_150_s_0_840=4.10e-11
+  mcl1p1f_ca_w_0_150_s_1_260=1.58e-04 mcl1p1f_cc_w_0_150_s_1_260=2.26e-12 mcl1p1f_cf_w_0_150_s_1_260=4.57e-11
+  mcl1p1f_ca_w_0_150_s_2_310=1.58e-04 mcl1p1f_cc_w_0_150_s_2_310=1.80e-13 mcl1p1f_cf_w_0_150_s_2_310=4.76e-11
+  mcl1p1f_ca_w_0_150_s_5_250=1.58e-04 mcl1p1f_cc_w_0_150_s_5_250=0.00e+00 mcl1p1f_cf_w_0_150_s_5_250=4.78e-11
+  mcl1p1f_ca_w_1_200_s_0_210=1.58e-04 mcl1p1f_cc_w_1_200_s_0_210=6.23e-11 mcl1p1f_cf_w_1_200_s_0_210=1.62e-11
+  mcl1p1f_ca_w_1_200_s_0_263=1.58e-04 mcl1p1f_cc_w_1_200_s_0_263=4.94e-11 mcl1p1f_cf_w_1_200_s_0_263=1.95e-11
+  mcl1p1f_ca_w_1_200_s_0_315=1.58e-04 mcl1p1f_cc_w_1_200_s_0_315=4.04e-11 mcl1p1f_cf_w_1_200_s_0_315=2.26e-11
+  mcl1p1f_ca_w_1_200_s_0_420=1.58e-04 mcl1p1f_cc_w_1_200_s_0_420=2.81e-11 mcl1p1f_cf_w_1_200_s_0_420=2.81e-11
+  mcl1p1f_ca_w_1_200_s_0_525=1.58e-04 mcl1p1f_cc_w_1_200_s_0_525=2.01e-11 mcl1p1f_cf_w_1_200_s_0_525=3.27e-11
+  mcl1p1f_ca_w_1_200_s_0_630=1.58e-04 mcl1p1f_cc_w_1_200_s_0_630=1.48e-11 mcl1p1f_cf_w_1_200_s_0_630=3.64e-11
+  mcl1p1f_ca_w_1_200_s_0_840=1.58e-04 mcl1p1f_cc_w_1_200_s_0_840=8.05e-12 mcl1p1f_cf_w_1_200_s_0_840=4.17e-11
+  mcl1p1f_ca_w_1_200_s_1_260=1.58e-04 mcl1p1f_cc_w_1_200_s_1_260=2.50e-12 mcl1p1f_cf_w_1_200_s_1_260=4.67e-11
+  mcl1p1f_ca_w_1_200_s_2_310=1.58e-04 mcl1p1f_cc_w_1_200_s_2_310=2.00e-13 mcl1p1f_cf_w_1_200_s_2_310=4.89e-11
+  mcl1p1f_ca_w_1_200_s_5_250=1.58e-04 mcl1p1f_cc_w_1_200_s_5_250=0.00e+00 mcl1p1f_cf_w_1_200_s_5_250=4.91e-11
+  mcm1p1f_ca_w_0_150_s_0_210=1.22e-04 mcm1p1f_cc_w_0_150_s_0_210=6.32e-11 mcm1p1f_cf_w_0_150_s_0_210=1.29e-11
+  mcm1p1f_ca_w_0_150_s_0_263=1.22e-04 mcm1p1f_cc_w_0_150_s_0_263=5.12e-11 mcm1p1f_cf_w_0_150_s_0_263=1.55e-11
+  mcm1p1f_ca_w_0_150_s_0_315=1.22e-04 mcm1p1f_cc_w_0_150_s_0_315=4.27e-11 mcm1p1f_cf_w_0_150_s_0_315=1.79e-11
+  mcm1p1f_ca_w_0_150_s_0_420=1.22e-04 mcm1p1f_cc_w_0_150_s_0_420=3.14e-11 mcm1p1f_cf_w_0_150_s_0_420=2.25e-11
+  mcm1p1f_ca_w_0_150_s_0_525=1.22e-04 mcm1p1f_cc_w_0_150_s_0_525=2.39e-11 mcm1p1f_cf_w_0_150_s_0_525=2.64e-11
+  mcm1p1f_ca_w_0_150_s_0_630=1.22e-04 mcm1p1f_cc_w_0_150_s_0_630=1.85e-11 mcm1p1f_cf_w_0_150_s_0_630=2.97e-11
+  mcm1p1f_ca_w_0_150_s_0_840=1.22e-04 mcm1p1f_cc_w_0_150_s_0_840=1.15e-11 mcm1p1f_cf_w_0_150_s_0_840=3.47e-11
+  mcm1p1f_ca_w_0_150_s_1_260=1.22e-04 mcm1p1f_cc_w_0_150_s_1_260=4.81e-12 mcm1p1f_cf_w_0_150_s_1_260=4.04e-11
+  mcm1p1f_ca_w_0_150_s_2_310=1.22e-04 mcm1p1f_cc_w_0_150_s_2_310=6.35e-13 mcm1p1f_cf_w_0_150_s_2_310=4.42e-11
+  mcm1p1f_ca_w_0_150_s_5_250=1.22e-04 mcm1p1f_cc_w_0_150_s_5_250=2.50e-14 mcm1p1f_cf_w_0_150_s_5_250=4.49e-11
+  mcm1p1f_ca_w_1_200_s_0_210=1.22e-04 mcm1p1f_cc_w_1_200_s_0_210=7.01e-11 mcm1p1f_cf_w_1_200_s_0_210=1.28e-11
+  mcm1p1f_ca_w_1_200_s_0_263=1.22e-04 mcm1p1f_cc_w_1_200_s_0_263=5.70e-11 mcm1p1f_cf_w_1_200_s_0_263=1.55e-11
+  mcm1p1f_ca_w_1_200_s_0_315=1.22e-04 mcm1p1f_cc_w_1_200_s_0_315=4.78e-11 mcm1p1f_cf_w_1_200_s_0_315=1.80e-11
+  mcm1p1f_ca_w_1_200_s_0_420=1.22e-04 mcm1p1f_cc_w_1_200_s_0_420=3.54e-11 mcm1p1f_cf_w_1_200_s_0_420=2.26e-11
+  mcm1p1f_ca_w_1_200_s_0_525=1.22e-04 mcm1p1f_cc_w_1_200_s_0_525=2.72e-11 mcm1p1f_cf_w_1_200_s_0_525=2.67e-11
+  mcm1p1f_ca_w_1_200_s_0_630=1.22e-04 mcm1p1f_cc_w_1_200_s_0_630=2.13e-11 mcm1p1f_cf_w_1_200_s_0_630=3.01e-11
+  mcm1p1f_ca_w_1_200_s_0_840=1.22e-04 mcm1p1f_cc_w_1_200_s_0_840=1.35e-11 mcm1p1f_cf_w_1_200_s_0_840=3.55e-11
+  mcm1p1f_ca_w_1_200_s_1_260=1.22e-04 mcm1p1f_cc_w_1_200_s_1_260=5.80e-12 mcm1p1f_cf_w_1_200_s_1_260=4.19e-11
+  mcm1p1f_ca_w_1_200_s_2_310=1.22e-04 mcm1p1f_cc_w_1_200_s_2_310=8.40e-13 mcm1p1f_cf_w_1_200_s_2_310=4.66e-11
+  mcm1p1f_ca_w_1_200_s_5_250=1.22e-04 mcm1p1f_cc_w_1_200_s_5_250=2.00e-14 mcm1p1f_cf_w_1_200_s_5_250=4.74e-11
+  mcm2p1f_ca_w_0_150_s_0_210=1.07e-04 mcm2p1f_cc_w_0_150_s_0_210=6.54e-11 mcm2p1f_cf_w_0_150_s_0_210=1.13e-11
+  mcm2p1f_ca_w_0_150_s_0_263=1.07e-04 mcm2p1f_cc_w_0_150_s_0_263=5.35e-11 mcm2p1f_cf_w_0_150_s_0_263=1.36e-11
+  mcm2p1f_ca_w_0_150_s_0_315=1.07e-04 mcm2p1f_cc_w_0_150_s_0_315=4.54e-11 mcm2p1f_cf_w_0_150_s_0_315=1.58e-11
+  mcm2p1f_ca_w_0_150_s_0_420=1.07e-04 mcm2p1f_cc_w_0_150_s_0_420=3.42e-11 mcm2p1f_cf_w_0_150_s_0_420=1.99e-11
+  mcm2p1f_ca_w_0_150_s_0_525=1.07e-04 mcm2p1f_cc_w_0_150_s_0_525=2.69e-11 mcm2p1f_cf_w_0_150_s_0_525=2.34e-11
+  mcm2p1f_ca_w_0_150_s_0_630=1.07e-04 mcm2p1f_cc_w_0_150_s_0_630=2.16e-11 mcm2p1f_cf_w_0_150_s_0_630=2.64e-11
+  mcm2p1f_ca_w_0_150_s_0_840=1.07e-04 mcm2p1f_cc_w_0_150_s_0_840=1.45e-11 mcm2p1f_cf_w_0_150_s_0_840=3.13e-11
+  mcm2p1f_ca_w_0_150_s_1_260=1.07e-04 mcm2p1f_cc_w_0_150_s_1_260=7.08e-12 mcm2p1f_cf_w_0_150_s_1_260=3.73e-11
+  mcm2p1f_ca_w_0_150_s_2_310=1.07e-04 mcm2p1f_cc_w_0_150_s_2_310=1.56e-12 mcm2p1f_cf_w_0_150_s_2_310=4.23e-11
+  mcm2p1f_ca_w_0_150_s_5_250=1.07e-04 mcm2p1f_cc_w_0_150_s_5_250=4.50e-14 mcm2p1f_cf_w_0_150_s_5_250=4.38e-11
+  mcm2p1f_ca_w_1_200_s_0_210=1.07e-04 mcm2p1f_cc_w_1_200_s_0_210=7.57e-11 mcm2p1f_cf_w_1_200_s_0_210=1.12e-11
+  mcm2p1f_ca_w_1_200_s_0_263=1.07e-04 mcm2p1f_cc_w_1_200_s_0_263=6.26e-11 mcm2p1f_cf_w_1_200_s_0_263=1.36e-11
+  mcm2p1f_ca_w_1_200_s_0_315=1.07e-04 mcm2p1f_cc_w_1_200_s_0_315=5.35e-11 mcm2p1f_cf_w_1_200_s_0_315=1.58e-11
+  mcm2p1f_ca_w_1_200_s_0_420=1.07e-04 mcm2p1f_cc_w_1_200_s_0_420=4.11e-11 mcm2p1f_cf_w_1_200_s_0_420=1.99e-11
+  mcm2p1f_ca_w_1_200_s_0_525=1.07e-04 mcm2p1f_cc_w_1_200_s_0_525=3.28e-11 mcm2p1f_cf_w_1_200_s_0_525=2.36e-11
+  mcm2p1f_ca_w_1_200_s_0_630=1.07e-04 mcm2p1f_cc_w_1_200_s_0_630=2.67e-11 mcm2p1f_cf_w_1_200_s_0_630=2.68e-11
+  mcm2p1f_ca_w_1_200_s_0_840=1.07e-04 mcm2p1f_cc_w_1_200_s_0_840=1.86e-11 mcm2p1f_cf_w_1_200_s_0_840=3.20e-11
+  mcm2p1f_ca_w_1_200_s_1_260=1.07e-04 mcm2p1f_cc_w_1_200_s_1_260=9.69e-12 mcm2p1f_cf_w_1_200_s_1_260=3.89e-11
+  mcm2p1f_ca_w_1_200_s_2_310=1.07e-04 mcm2p1f_cc_w_1_200_s_2_310=2.27e-12 mcm2p1f_cf_w_1_200_s_2_310=4.56e-11
+  mcm2p1f_ca_w_1_200_s_5_250=1.07e-04 mcm2p1f_cc_w_1_200_s_5_250=9.00e-14 mcm2p1f_cf_w_1_200_s_5_250=4.77e-11
+  mcm3p1f_ca_w_0_150_s_0_210=1.00e-04 mcm3p1f_cc_w_0_150_s_0_210=6.64e-11 mcm3p1f_cf_w_0_150_s_0_210=1.06e-11
+  mcm3p1f_ca_w_0_150_s_0_263=1.00e-04 mcm3p1f_cc_w_0_150_s_0_263=5.47e-11 mcm3p1f_cf_w_0_150_s_0_263=1.27e-11
+  mcm3p1f_ca_w_0_150_s_0_315=1.00e-04 mcm3p1f_cc_w_0_150_s_0_315=4.67e-11 mcm3p1f_cf_w_0_150_s_0_315=1.47e-11
+  mcm3p1f_ca_w_0_150_s_0_420=1.00e-04 mcm3p1f_cc_w_0_150_s_0_420=3.57e-11 mcm3p1f_cf_w_0_150_s_0_420=1.86e-11
+  mcm3p1f_ca_w_0_150_s_0_525=1.00e-04 mcm3p1f_cc_w_0_150_s_0_525=2.85e-11 mcm3p1f_cf_w_0_150_s_0_525=2.19e-11
+  mcm3p1f_ca_w_0_150_s_0_630=1.00e-04 mcm3p1f_cc_w_0_150_s_0_630=2.33e-11 mcm3p1f_cf_w_0_150_s_0_630=2.48e-11
+  mcm3p1f_ca_w_0_150_s_0_840=1.00e-04 mcm3p1f_cc_w_0_150_s_0_840=1.63e-11 mcm3p1f_cf_w_0_150_s_0_840=2.95e-11
+  mcm3p1f_ca_w_0_150_s_1_260=1.00e-04 mcm3p1f_cc_w_0_150_s_1_260=8.50e-12 mcm3p1f_cf_w_0_150_s_1_260=3.57e-11
+  mcm3p1f_ca_w_0_150_s_2_310=1.00e-04 mcm3p1f_cc_w_0_150_s_2_310=2.36e-12 mcm3p1f_cf_w_0_150_s_2_310=4.12e-11
+  mcm3p1f_ca_w_0_150_s_5_250=1.00e-04 mcm3p1f_cc_w_0_150_s_5_250=1.70e-13 mcm3p1f_cf_w_0_150_s_5_250=4.34e-11
+  mcm3p1f_ca_w_1_200_s_0_210=1.00e-04 mcm3p1f_cc_w_1_200_s_0_210=7.91e-11 mcm3p1f_cf_w_1_200_s_0_210=1.05e-11
+  mcm3p1f_ca_w_1_200_s_0_263=1.00e-04 mcm3p1f_cc_w_1_200_s_0_263=6.60e-11 mcm3p1f_cf_w_1_200_s_0_263=1.27e-11
+  mcm3p1f_ca_w_1_200_s_0_315=1.00e-04 mcm3p1f_cc_w_1_200_s_0_315=5.70e-11 mcm3p1f_cf_w_1_200_s_0_315=1.48e-11
+  mcm3p1f_ca_w_1_200_s_0_420=1.00e-04 mcm3p1f_cc_w_1_200_s_0_420=4.45e-11 mcm3p1f_cf_w_1_200_s_0_420=1.86e-11
+  mcm3p1f_ca_w_1_200_s_0_525=1.00e-04 mcm3p1f_cc_w_1_200_s_0_525=3.63e-11 mcm3p1f_cf_w_1_200_s_0_525=2.21e-11
+  mcm3p1f_ca_w_1_200_s_0_630=1.00e-04 mcm3p1f_cc_w_1_200_s_0_630=3.02e-11 mcm3p1f_cf_w_1_200_s_0_630=2.52e-11
+  mcm3p1f_ca_w_1_200_s_0_840=1.00e-04 mcm3p1f_cc_w_1_200_s_0_840=2.19e-11 mcm3p1f_cf_w_1_200_s_0_840=3.03e-11
+  mcm3p1f_ca_w_1_200_s_1_260=1.00e-04 mcm3p1f_cc_w_1_200_s_1_260=1.25e-11 mcm3p1f_cf_w_1_200_s_1_260=3.72e-11
+  mcm3p1f_ca_w_1_200_s_2_310=1.00e-04 mcm3p1f_cc_w_1_200_s_2_310=3.86e-12 mcm3p1f_cf_w_1_200_s_2_310=4.48e-11
+  mcm3p1f_ca_w_1_200_s_5_250=1.00e-04 mcm3p1f_cc_w_1_200_s_5_250=2.75e-13 mcm3p1f_cf_w_1_200_s_5_250=4.84e-11
+  mcm4p1f_ca_w_0_150_s_0_210=9.56e-05 mcm4p1f_cc_w_0_150_s_0_210=6.71e-11 mcm4p1f_cf_w_0_150_s_0_210=1.01e-11
+  mcm4p1f_ca_w_0_150_s_0_263=9.56e-05 mcm4p1f_cc_w_0_150_s_0_263=5.54e-11 mcm4p1f_cf_w_0_150_s_0_263=1.21e-11
+  mcm4p1f_ca_w_0_150_s_0_315=9.56e-05 mcm4p1f_cc_w_0_150_s_0_315=4.75e-11 mcm4p1f_cf_w_0_150_s_0_315=1.40e-11
+  mcm4p1f_ca_w_0_150_s_0_420=9.56e-05 mcm4p1f_cc_w_0_150_s_0_420=3.66e-11 mcm4p1f_cf_w_0_150_s_0_420=1.77e-11
+  mcm4p1f_ca_w_0_150_s_0_525=9.56e-05 mcm4p1f_cc_w_0_150_s_0_525=2.96e-11 mcm4p1f_cf_w_0_150_s_0_525=2.09e-11
+  mcm4p1f_ca_w_0_150_s_0_630=9.56e-05 mcm4p1f_cc_w_0_150_s_0_630=2.45e-11 mcm4p1f_cf_w_0_150_s_0_630=2.37e-11
+  mcm4p1f_ca_w_0_150_s_0_840=9.56e-05 mcm4p1f_cc_w_0_150_s_0_840=1.75e-11 mcm4p1f_cf_w_0_150_s_0_840=2.83e-11
+  mcm4p1f_ca_w_0_150_s_1_260=9.56e-05 mcm4p1f_cc_w_0_150_s_1_260=9.60e-12 mcm4p1f_cf_w_0_150_s_1_260=3.46e-11
+  mcm4p1f_ca_w_0_150_s_2_310=9.56e-05 mcm4p1f_cc_w_0_150_s_2_310=3.12e-12 mcm4p1f_cf_w_0_150_s_2_310=4.03e-11
+  mcm4p1f_ca_w_0_150_s_5_250=9.56e-05 mcm4p1f_cc_w_0_150_s_5_250=3.35e-13 mcm4p1f_cf_w_0_150_s_5_250=4.31e-11
+  mcm4p1f_ca_w_1_200_s_0_210=9.56e-05 mcm4p1f_cc_w_1_200_s_0_210=8.15e-11 mcm4p1f_cf_w_1_200_s_0_210=1.00e-11
+  mcm4p1f_ca_w_1_200_s_0_263=9.56e-05 mcm4p1f_cc_w_1_200_s_0_263=6.86e-11 mcm4p1f_cf_w_1_200_s_0_263=1.21e-11
+  mcm4p1f_ca_w_1_200_s_0_315=9.56e-05 mcm4p1f_cc_w_1_200_s_0_315=5.96e-11 mcm4p1f_cf_w_1_200_s_0_315=1.41e-11
+  mcm4p1f_ca_w_1_200_s_0_420=9.56e-05 mcm4p1f_cc_w_1_200_s_0_420=4.72e-11 mcm4p1f_cf_w_1_200_s_0_420=1.78e-11
+  mcm4p1f_ca_w_1_200_s_0_525=9.56e-05 mcm4p1f_cc_w_1_200_s_0_525=3.89e-11 mcm4p1f_cf_w_1_200_s_0_525=2.11e-11
+  mcm4p1f_ca_w_1_200_s_0_630=9.56e-05 mcm4p1f_cc_w_1_200_s_0_630=3.29e-11 mcm4p1f_cf_w_1_200_s_0_630=2.40e-11
+  mcm4p1f_ca_w_1_200_s_0_840=9.56e-05 mcm4p1f_cc_w_1_200_s_0_840=2.46e-11 mcm4p1f_cf_w_1_200_s_0_840=2.90e-11
+  mcm4p1f_ca_w_1_200_s_1_260=9.56e-05 mcm4p1f_cc_w_1_200_s_1_260=1.51e-11 mcm4p1f_cf_w_1_200_s_1_260=3.59e-11
+  mcm4p1f_ca_w_1_200_s_2_310=9.56e-05 mcm4p1f_cc_w_1_200_s_2_310=5.65e-12 mcm4p1f_cf_w_1_200_s_2_310=4.41e-11
+  mcm4p1f_ca_w_1_200_s_5_250=9.56e-05 mcm4p1f_cc_w_1_200_s_5_250=5.85e-13 mcm4p1f_cf_w_1_200_s_5_250=4.89e-11
+  mcm5p1f_ca_w_0_150_s_0_210=9.32e-05 mcm5p1f_cc_w_0_150_s_0_210=6.74e-11 mcm5p1f_cf_w_0_150_s_0_210=9.81e-12
+  mcm5p1f_ca_w_0_150_s_0_263=9.32e-05 mcm5p1f_cc_w_0_150_s_0_263=5.58e-11 mcm5p1f_cf_w_0_150_s_0_263=1.18e-11
+  mcm5p1f_ca_w_0_150_s_0_315=9.32e-05 mcm5p1f_cc_w_0_150_s_0_315=4.80e-11 mcm5p1f_cf_w_0_150_s_0_315=1.37e-11
+  mcm5p1f_ca_w_0_150_s_0_420=9.32e-05 mcm5p1f_cc_w_0_150_s_0_420=3.71e-11 mcm5p1f_cf_w_0_150_s_0_420=1.73e-11
+  mcm5p1f_ca_w_0_150_s_0_525=9.32e-05 mcm5p1f_cc_w_0_150_s_0_525=3.02e-11 mcm5p1f_cf_w_0_150_s_0_525=2.04e-11
+  mcm5p1f_ca_w_0_150_s_0_630=9.32e-05 mcm5p1f_cc_w_0_150_s_0_630=2.52e-11 mcm5p1f_cf_w_0_150_s_0_630=2.31e-11
+  mcm5p1f_ca_w_0_150_s_0_840=9.32e-05 mcm5p1f_cc_w_0_150_s_0_840=1.82e-11 mcm5p1f_cf_w_0_150_s_0_840=2.76e-11
+  mcm5p1f_ca_w_0_150_s_1_260=9.32e-05 mcm5p1f_cc_w_0_150_s_1_260=1.02e-11 mcm5p1f_cf_w_0_150_s_1_260=3.40e-11
+  mcm5p1f_ca_w_0_150_s_2_310=9.32e-05 mcm5p1f_cc_w_0_150_s_2_310=3.63e-12 mcm5p1f_cf_w_0_150_s_2_310=3.98e-11
+  mcm5p1f_ca_w_0_150_s_5_250=9.32e-05 mcm5p1f_cc_w_0_150_s_5_250=4.92e-13 mcm5p1f_cf_w_0_150_s_5_250=4.29e-11
+  mcm5p1f_ca_w_1_200_s_0_210=9.32e-05 mcm5p1f_cc_w_1_200_s_0_210=8.29e-11 mcm5p1f_cf_w_1_200_s_0_210=9.74e-12
+  mcm5p1f_ca_w_1_200_s_0_263=9.32e-05 mcm5p1f_cc_w_1_200_s_0_263=7.00e-11 mcm5p1f_cf_w_1_200_s_0_263=1.18e-11
+  mcm5p1f_ca_w_1_200_s_0_315=9.32e-05 mcm5p1f_cc_w_1_200_s_0_315=6.10e-11 mcm5p1f_cf_w_1_200_s_0_315=1.37e-11
+  mcm5p1f_ca_w_1_200_s_0_420=9.32e-05 mcm5p1f_cc_w_1_200_s_0_420=4.88e-11 mcm5p1f_cf_w_1_200_s_0_420=1.73e-11
+  mcm5p1f_ca_w_1_200_s_0_525=9.32e-05 mcm5p1f_cc_w_1_200_s_0_525=4.06e-11 mcm5p1f_cf_w_1_200_s_0_525=2.05e-11
+  mcm5p1f_ca_w_1_200_s_0_630=9.32e-05 mcm5p1f_cc_w_1_200_s_0_630=3.46e-11 mcm5p1f_cf_w_1_200_s_0_630=2.34e-11
+  mcm5p1f_ca_w_1_200_s_0_840=9.32e-05 mcm5p1f_cc_w_1_200_s_0_840=2.62e-11 mcm5p1f_cf_w_1_200_s_0_840=2.83e-11
+  mcm5p1f_ca_w_1_200_s_1_260=9.32e-05 mcm5p1f_cc_w_1_200_s_1_260=1.66e-11 mcm5p1f_cf_w_1_200_s_1_260=3.52e-11
+  mcm5p1f_ca_w_1_200_s_2_310=9.32e-05 mcm5p1f_cc_w_1_200_s_2_310=6.78e-12 mcm5p1f_cf_w_1_200_s_2_310=4.37e-11
+  mcm5p1f_ca_w_1_200_s_5_250=9.32e-05 mcm5p1f_cc_w_1_200_s_5_250=1.05e-12 mcm5p1f_cf_w_1_200_s_5_250=4.92e-11
+  mcrdlp1f_ca_w_0_150_s_0_210=8.90e-05 mcrdlp1f_cc_w_0_150_s_0_210=6.80e-11 mcrdlp1f_cf_w_0_150_s_0_210=9.34e-12
+  mcrdlp1f_ca_w_0_150_s_0_263=8.90e-05 mcrdlp1f_cc_w_0_150_s_0_263=5.64e-11 mcrdlp1f_cf_w_0_150_s_0_263=1.12e-11
+  mcrdlp1f_ca_w_0_150_s_0_315=8.90e-05 mcrdlp1f_cc_w_0_150_s_0_315=4.88e-11 mcrdlp1f_cf_w_0_150_s_0_315=1.30e-11
+  mcrdlp1f_ca_w_0_150_s_0_420=8.90e-05 mcrdlp1f_cc_w_0_150_s_0_420=3.79e-11 mcrdlp1f_cf_w_0_150_s_0_420=1.65e-11
+  mcrdlp1f_ca_w_0_150_s_0_525=8.90e-05 mcrdlp1f_cc_w_0_150_s_0_525=3.12e-11 mcrdlp1f_cf_w_0_150_s_0_525=1.94e-11
+  mcrdlp1f_ca_w_0_150_s_0_630=8.90e-05 mcrdlp1f_cc_w_0_150_s_0_630=2.63e-11 mcrdlp1f_cf_w_0_150_s_0_630=2.20e-11
+  mcrdlp1f_ca_w_0_150_s_0_840=8.90e-05 mcrdlp1f_cc_w_0_150_s_0_840=1.94e-11 mcrdlp1f_cf_w_0_150_s_0_840=2.65e-11
+  mcrdlp1f_ca_w_0_150_s_1_260=8.90e-05 mcrdlp1f_cc_w_0_150_s_1_260=1.14e-11 mcrdlp1f_cf_w_0_150_s_1_260=3.28e-11
+  mcrdlp1f_ca_w_0_150_s_2_310=8.90e-05 mcrdlp1f_cc_w_0_150_s_2_310=4.65e-12 mcrdlp1f_cf_w_0_150_s_2_310=3.89e-11
+  mcrdlp1f_ca_w_0_150_s_5_250=8.90e-05 mcrdlp1f_cc_w_0_150_s_5_250=9.24e-13 mcrdlp1f_cf_w_0_150_s_5_250=4.25e-11
+  mcrdlp1f_ca_w_1_200_s_0_210=8.90e-05 mcrdlp1f_cc_w_1_200_s_0_210=8.53e-11 mcrdlp1f_cf_w_1_200_s_0_210=9.27e-12
+  mcrdlp1f_ca_w_1_200_s_0_263=8.90e-05 mcrdlp1f_cc_w_1_200_s_0_263=7.25e-11 mcrdlp1f_cf_w_1_200_s_0_263=1.12e-11
+  mcrdlp1f_ca_w_1_200_s_0_315=8.90e-05 mcrdlp1f_cc_w_1_200_s_0_315=6.36e-11 mcrdlp1f_cf_w_1_200_s_0_315=1.31e-11
+  mcrdlp1f_ca_w_1_200_s_0_420=8.90e-05 mcrdlp1f_cc_w_1_200_s_0_420=5.14e-11 mcrdlp1f_cf_w_1_200_s_0_420=1.65e-11
+  mcrdlp1f_ca_w_1_200_s_0_525=8.90e-05 mcrdlp1f_cc_w_1_200_s_0_525=4.34e-11 mcrdlp1f_cf_w_1_200_s_0_525=1.96e-11
+  mcrdlp1f_ca_w_1_200_s_0_630=8.90e-05 mcrdlp1f_cc_w_1_200_s_0_630=3.75e-11 mcrdlp1f_cf_w_1_200_s_0_630=2.23e-11
+  mcrdlp1f_ca_w_1_200_s_0_840=8.90e-05 mcrdlp1f_cc_w_1_200_s_0_840=2.92e-11 mcrdlp1f_cf_w_1_200_s_0_840=2.71e-11
+  mcrdlp1f_ca_w_1_200_s_1_260=8.90e-05 mcrdlp1f_cc_w_1_200_s_1_260=1.97e-11 mcrdlp1f_cf_w_1_200_s_1_260=3.39e-11
+  mcrdlp1f_ca_w_1_200_s_2_310=8.90e-05 mcrdlp1f_cc_w_1_200_s_2_310=9.36e-12 mcrdlp1f_cf_w_1_200_s_2_310=4.28e-11
+  mcrdlp1f_ca_w_1_200_s_5_250=8.90e-05 mcrdlp1f_cc_w_1_200_s_5_250=2.40e-12 mcrdlp1f_cf_w_1_200_s_5_250=4.95e-11
+  mcm1l1f_ca_w_0_170_s_0_180=1.19e-04 mcm1l1f_cc_w_0_170_s_0_180=5.82e-11 mcm1l1f_cf_w_0_170_s_0_180=1.12e-11
+  mcm1l1f_ca_w_0_170_s_0_225=1.19e-04 mcm1l1f_cc_w_0_170_s_0_225=4.89e-11 mcm1l1f_cf_w_0_170_s_0_225=1.35e-11
+  mcm1l1f_ca_w_0_170_s_0_270=1.19e-04 mcm1l1f_cc_w_0_170_s_0_270=4.19e-11 mcm1l1f_cf_w_0_170_s_0_270=1.55e-11
+  mcm1l1f_ca_w_0_170_s_0_360=1.19e-04 mcm1l1f_cc_w_0_170_s_0_360=3.19e-11 mcm1l1f_cf_w_0_170_s_0_360=1.95e-11
+  mcm1l1f_ca_w_0_170_s_0_450=1.19e-04 mcm1l1f_cc_w_0_170_s_0_450=2.52e-11 mcm1l1f_cf_w_0_170_s_0_450=2.28e-11
+  mcm1l1f_ca_w_0_170_s_0_540=1.19e-04 mcm1l1f_cc_w_0_170_s_0_540=2.02e-11 mcm1l1f_cf_w_0_170_s_0_540=2.58e-11
+  mcm1l1f_ca_w_0_170_s_0_720=1.19e-04 mcm1l1f_cc_w_0_170_s_0_720=1.34e-11 mcm1l1f_cf_w_0_170_s_0_720=3.05e-11
+  mcm1l1f_ca_w_0_170_s_1_080=1.19e-04 mcm1l1f_cc_w_0_170_s_1_080=6.23e-12 mcm1l1f_cf_w_0_170_s_1_080=3.63e-11
+  mcm1l1f_ca_w_0_170_s_1_980=1.19e-04 mcm1l1f_cc_w_0_170_s_1_980=1.05e-12 mcm1l1f_cf_w_0_170_s_1_980=4.10e-11
+  mcm1l1f_ca_w_0_170_s_4_500=1.19e-04 mcm1l1f_cc_w_0_170_s_4_500=5.00e-14 mcm1l1f_cf_w_0_170_s_4_500=4.20e-11
+  mcm1l1f_ca_w_1_360_s_0_180=1.19e-04 mcm1l1f_cc_w_1_360_s_0_180=6.54e-11 mcm1l1f_cf_w_1_360_s_0_180=1.12e-11
+  mcm1l1f_ca_w_1_360_s_0_225=1.19e-04 mcm1l1f_cc_w_1_360_s_0_225=5.51e-11 mcm1l1f_cf_w_1_360_s_0_225=1.34e-11
+  mcm1l1f_ca_w_1_360_s_0_270=1.19e-04 mcm1l1f_cc_w_1_360_s_0_270=4.76e-11 mcm1l1f_cf_w_1_360_s_0_270=1.56e-11
+  mcm1l1f_ca_w_1_360_s_0_360=1.19e-04 mcm1l1f_cc_w_1_360_s_0_360=3.66e-11 mcm1l1f_cf_w_1_360_s_0_360=1.95e-11
+  mcm1l1f_ca_w_1_360_s_0_450=1.19e-04 mcm1l1f_cc_w_1_360_s_0_450=2.91e-11 mcm1l1f_cf_w_1_360_s_0_450=2.30e-11
+  mcm1l1f_ca_w_1_360_s_0_540=1.19e-04 mcm1l1f_cc_w_1_360_s_0_540=2.35e-11 mcm1l1f_cf_w_1_360_s_0_540=2.61e-11
+  mcm1l1f_ca_w_1_360_s_0_720=1.19e-04 mcm1l1f_cc_w_1_360_s_0_720=1.59e-11 mcm1l1f_cf_w_1_360_s_0_720=3.12e-11
+  mcm1l1f_ca_w_1_360_s_1_080=1.19e-04 mcm1l1f_cc_w_1_360_s_1_080=7.61e-12 mcm1l1f_cf_w_1_360_s_1_080=3.77e-11
+  mcm1l1f_ca_w_1_360_s_1_980=1.19e-04 mcm1l1f_cc_w_1_360_s_1_980=1.40e-12 mcm1l1f_cf_w_1_360_s_1_980=4.34e-11
+  mcm1l1f_ca_w_1_360_s_4_500=1.19e-04 mcm1l1f_cc_w_1_360_s_4_500=1.50e-14 mcm1l1f_cf_w_1_360_s_4_500=4.47e-11
+  mcm1l1d_ca_w_0_170_s_0_180=1.35e-04 mcm1l1d_cc_w_0_170_s_0_180=5.61e-11 mcm1l1d_cf_w_0_170_s_0_180=1.28e-11
+  mcm1l1d_ca_w_0_170_s_0_225=1.35e-04 mcm1l1d_cc_w_0_170_s_0_225=4.66e-11 mcm1l1d_cf_w_0_170_s_0_225=1.53e-11
+  mcm1l1d_ca_w_0_170_s_0_270=1.35e-04 mcm1l1d_cc_w_0_170_s_0_270=3.94e-11 mcm1l1d_cf_w_0_170_s_0_270=1.76e-11
+  mcm1l1d_ca_w_0_170_s_0_360=1.35e-04 mcm1l1d_cc_w_0_170_s_0_360=2.93e-11 mcm1l1d_cf_w_0_170_s_0_360=2.19e-11
+  mcm1l1d_ca_w_0_170_s_0_450=1.35e-04 mcm1l1d_cc_w_0_170_s_0_450=2.25e-11 mcm1l1d_cf_w_0_170_s_0_450=2.56e-11
+  mcm1l1d_ca_w_0_170_s_0_540=1.35e-04 mcm1l1d_cc_w_0_170_s_0_540=1.75e-11 mcm1l1d_cf_w_0_170_s_0_540=2.87e-11
+  mcm1l1d_ca_w_0_170_s_0_720=1.35e-04 mcm1l1d_cc_w_0_170_s_0_720=1.09e-11 mcm1l1d_cf_w_0_170_s_0_720=3.35e-11
+  mcm1l1d_ca_w_0_170_s_1_080=1.35e-04 mcm1l1d_cc_w_0_170_s_1_080=4.41e-12 mcm1l1d_cf_w_0_170_s_1_080=3.90e-11
+  mcm1l1d_ca_w_0_170_s_1_980=1.35e-04 mcm1l1d_cc_w_0_170_s_1_980=5.05e-13 mcm1l1d_cf_w_0_170_s_1_980=4.27e-11
+  mcm1l1d_ca_w_0_170_s_4_500=1.35e-04 mcm1l1d_cc_w_0_170_s_4_500=4.50e-14 mcm1l1d_cf_w_0_170_s_4_500=4.32e-11
+  mcm1l1d_ca_w_1_360_s_0_180=1.35e-04 mcm1l1d_cc_w_1_360_s_0_180=6.12e-11 mcm1l1d_cf_w_1_360_s_0_180=1.27e-11
+  mcm1l1d_ca_w_1_360_s_0_225=1.35e-04 mcm1l1d_cc_w_1_360_s_0_225=5.12e-11 mcm1l1d_cf_w_1_360_s_0_225=1.52e-11
+  mcm1l1d_ca_w_1_360_s_0_270=1.35e-04 mcm1l1d_cc_w_1_360_s_0_270=4.33e-11 mcm1l1d_cf_w_1_360_s_0_270=1.76e-11
+  mcm1l1d_ca_w_1_360_s_0_360=1.35e-04 mcm1l1d_cc_w_1_360_s_0_360=3.25e-11 mcm1l1d_cf_w_1_360_s_0_360=2.20e-11
+  mcm1l1d_ca_w_1_360_s_0_450=1.35e-04 mcm1l1d_cc_w_1_360_s_0_450=2.50e-11 mcm1l1d_cf_w_1_360_s_0_450=2.58e-11
+  mcm1l1d_ca_w_1_360_s_0_540=1.35e-04 mcm1l1d_cc_w_1_360_s_0_540=1.96e-11 mcm1l1d_cf_w_1_360_s_0_540=2.91e-11
+  mcm1l1d_ca_w_1_360_s_0_720=1.35e-04 mcm1l1d_cc_w_1_360_s_0_720=1.23e-11 mcm1l1d_cf_w_1_360_s_0_720=3.42e-11
+  mcm1l1d_ca_w_1_360_s_1_080=1.35e-04 mcm1l1d_cc_w_1_360_s_1_080=5.00e-12 mcm1l1d_cf_w_1_360_s_1_080=4.03e-11
+  mcm1l1d_ca_w_1_360_s_1_980=1.35e-04 mcm1l1d_cc_w_1_360_s_1_980=6.25e-13 mcm1l1d_cf_w_1_360_s_1_980=4.44e-11
+  mcm1l1d_ca_w_1_360_s_4_500=1.35e-04 mcm1l1d_cc_w_1_360_s_4_500=0.00e+00 mcm1l1d_cf_w_1_360_s_4_500=4.50e-11
+  mcm1l1p1_ca_w_0_170_s_0_180=1.59e-04 mcm1l1p1_cc_w_0_170_s_0_180=5.33e-11 mcm1l1p1_cf_w_0_170_s_0_180=1.49e-11
+  mcm1l1p1_ca_w_0_170_s_0_225=1.59e-04 mcm1l1p1_cc_w_0_170_s_0_225=4.37e-11 mcm1l1p1_cf_w_0_170_s_0_225=1.78e-11
+  mcm1l1p1_ca_w_0_170_s_0_270=1.59e-04 mcm1l1p1_cc_w_0_170_s_0_270=3.65e-11 mcm1l1p1_cf_w_0_170_s_0_270=2.04e-11
+  mcm1l1p1_ca_w_0_170_s_0_360=1.59e-04 mcm1l1p1_cc_w_0_170_s_0_360=2.64e-11 mcm1l1p1_cf_w_0_170_s_0_360=2.52e-11
+  mcm1l1p1_ca_w_0_170_s_0_450=1.59e-04 mcm1l1p1_cc_w_0_170_s_0_450=1.95e-11 mcm1l1p1_cf_w_0_170_s_0_450=2.91e-11
+  mcm1l1p1_ca_w_0_170_s_0_540=1.59e-04 mcm1l1p1_cc_w_0_170_s_0_540=1.48e-11 mcm1l1p1_cf_w_0_170_s_0_540=3.25e-11
+  mcm1l1p1_ca_w_0_170_s_0_720=1.59e-04 mcm1l1p1_cc_w_0_170_s_0_720=8.55e-12 mcm1l1p1_cf_w_0_170_s_0_720=3.73e-11
+  mcm1l1p1_ca_w_0_170_s_1_080=1.59e-04 mcm1l1p1_cc_w_0_170_s_1_080=2.95e-12 mcm1l1p1_cf_w_0_170_s_1_080=4.22e-11
+  mcm1l1p1_ca_w_0_170_s_1_980=1.59e-04 mcm1l1p1_cc_w_0_170_s_1_980=2.40e-13 mcm1l1p1_cf_w_0_170_s_1_980=4.48e-11
+  mcm1l1p1_ca_w_0_170_s_4_500=1.59e-04 mcm1l1p1_cc_w_0_170_s_4_500=5.00e-15 mcm1l1p1_cf_w_0_170_s_4_500=4.50e-11
+  mcm1l1p1_ca_w_1_360_s_0_180=1.59e-04 mcm1l1p1_cc_w_1_360_s_0_180=5.67e-11 mcm1l1p1_cf_w_1_360_s_0_180=1.48e-11
+  mcm1l1p1_ca_w_1_360_s_0_225=1.59e-04 mcm1l1p1_cc_w_1_360_s_0_225=4.67e-11 mcm1l1p1_cf_w_1_360_s_0_225=1.77e-11
+  mcm1l1p1_ca_w_1_360_s_0_270=1.59e-04 mcm1l1p1_cc_w_1_360_s_0_270=3.90e-11 mcm1l1p1_cf_w_1_360_s_0_270=2.04e-11
+  mcm1l1p1_ca_w_1_360_s_0_360=1.59e-04 mcm1l1p1_cc_w_1_360_s_0_360=2.82e-11 mcm1l1p1_cf_w_1_360_s_0_360=2.52e-11
+  mcm1l1p1_ca_w_1_360_s_0_450=1.59e-04 mcm1l1p1_cc_w_1_360_s_0_450=2.10e-11 mcm1l1p1_cf_w_1_360_s_0_450=2.94e-11
+  mcm1l1p1_ca_w_1_360_s_0_540=1.59e-04 mcm1l1p1_cc_w_1_360_s_0_540=1.59e-11 mcm1l1p1_cf_w_1_360_s_0_540=3.28e-11
+  mcm1l1p1_ca_w_1_360_s_0_720=1.59e-04 mcm1l1p1_cc_w_1_360_s_0_720=9.25e-12 mcm1l1p1_cf_w_1_360_s_0_720=3.79e-11
+  mcm1l1p1_ca_w_1_360_s_1_080=1.59e-04 mcm1l1p1_cc_w_1_360_s_1_080=3.25e-12 mcm1l1p1_cf_w_1_360_s_1_080=4.31e-11
+  mcm1l1p1_ca_w_1_360_s_1_980=1.59e-04 mcm1l1p1_cc_w_1_360_s_1_980=3.00e-13 mcm1l1p1_cf_w_1_360_s_1_980=4.60e-11
+  mcm1l1p1_ca_w_1_360_s_4_500=1.59e-04 mcm1l1p1_cc_w_1_360_s_4_500=1.29e-26 mcm1l1p1_cf_w_1_360_s_4_500=4.62e-11
+  mcm2l1f_ca_w_0_170_s_0_180=6.22e-05 mcm2l1f_cc_w_0_170_s_0_180=6.50e-11 mcm2l1f_cf_w_0_170_s_0_180=6.15e-12
+  mcm2l1f_ca_w_0_170_s_0_225=6.22e-05 mcm2l1f_cc_w_0_170_s_0_225=5.59e-11 mcm2l1f_cf_w_0_170_s_0_225=7.44e-12
+  mcm2l1f_ca_w_0_170_s_0_270=6.22e-05 mcm2l1f_cc_w_0_170_s_0_270=4.93e-11 mcm2l1f_cf_w_0_170_s_0_270=8.66e-12
+  mcm2l1f_ca_w_0_170_s_0_360=6.22e-05 mcm2l1f_cc_w_0_170_s_0_360=3.96e-11 mcm2l1f_cf_w_0_170_s_0_360=1.12e-11
+  mcm2l1f_ca_w_0_170_s_0_450=6.22e-05 mcm2l1f_cc_w_0_170_s_0_450=3.32e-11 mcm2l1f_cf_w_0_170_s_0_450=1.33e-11
+  mcm2l1f_ca_w_0_170_s_0_540=6.22e-05 mcm2l1f_cc_w_0_170_s_0_540=2.80e-11 mcm2l1f_cf_w_0_170_s_0_540=1.54e-11
+  mcm2l1f_ca_w_0_170_s_0_720=6.22e-05 mcm2l1f_cc_w_0_170_s_0_720=2.09e-11 mcm2l1f_cf_w_0_170_s_0_720=1.91e-11
+  mcm2l1f_ca_w_0_170_s_1_080=6.22e-05 mcm2l1f_cc_w_0_170_s_1_080=1.23e-11 mcm2l1f_cf_w_0_170_s_1_080=2.46e-11
+  mcm2l1f_ca_w_0_170_s_1_980=6.22e-05 mcm2l1f_cc_w_0_170_s_1_980=3.62e-12 mcm2l1f_cf_w_0_170_s_1_980=3.17e-11
+  mcm2l1f_ca_w_0_170_s_4_500=6.22e-05 mcm2l1f_cc_w_0_170_s_4_500=1.70e-13 mcm2l1f_cf_w_0_170_s_4_500=3.49e-11
+  mcm2l1f_ca_w_1_360_s_0_180=6.22e-05 mcm2l1f_cc_w_1_360_s_0_180=7.66e-11 mcm2l1f_cf_w_1_360_s_0_180=6.12e-12
+  mcm2l1f_ca_w_1_360_s_0_225=6.22e-05 mcm2l1f_cc_w_1_360_s_0_225=6.64e-11 mcm2l1f_cf_w_1_360_s_0_225=7.41e-12
+  mcm2l1f_ca_w_1_360_s_0_270=6.22e-05 mcm2l1f_cc_w_1_360_s_0_270=5.87e-11 mcm2l1f_cf_w_1_360_s_0_270=8.68e-12
+  mcm2l1f_ca_w_1_360_s_0_360=6.22e-05 mcm2l1f_cc_w_1_360_s_0_360=4.75e-11 mcm2l1f_cf_w_1_360_s_0_360=1.11e-11
+  mcm2l1f_ca_w_1_360_s_0_450=6.22e-05 mcm2l1f_cc_w_1_360_s_0_450=3.97e-11 mcm2l1f_cf_w_1_360_s_0_450=1.34e-11
+  mcm2l1f_ca_w_1_360_s_0_540=6.22e-05 mcm2l1f_cc_w_1_360_s_0_540=3.38e-11 mcm2l1f_cf_w_1_360_s_0_540=1.56e-11
+  mcm2l1f_ca_w_1_360_s_0_720=6.22e-05 mcm2l1f_cc_w_1_360_s_0_720=2.53e-11 mcm2l1f_cf_w_1_360_s_0_720=1.95e-11
+  mcm2l1f_ca_w_1_360_s_1_080=6.22e-05 mcm2l1f_cc_w_1_360_s_1_080=1.50e-11 mcm2l1f_cf_w_1_360_s_1_080=2.57e-11
+  mcm2l1f_ca_w_1_360_s_1_980=6.22e-05 mcm2l1f_cc_w_1_360_s_1_980=4.57e-12 mcm2l1f_cf_w_1_360_s_1_980=3.40e-11
+  mcm2l1f_ca_w_1_360_s_4_500=6.22e-05 mcm2l1f_cc_w_1_360_s_4_500=2.00e-13 mcm2l1f_cf_w_1_360_s_4_500=3.81e-11
+  mcm2l1d_ca_w_0_170_s_0_180=7.87e-05 mcm2l1d_cc_w_0_170_s_0_180=6.27e-11 mcm2l1d_cf_w_0_170_s_0_180=7.72e-12
+  mcm2l1d_ca_w_0_170_s_0_225=7.87e-05 mcm2l1d_cc_w_0_170_s_0_225=5.35e-11 mcm2l1d_cf_w_0_170_s_0_225=9.33e-12
+  mcm2l1d_ca_w_0_170_s_0_270=7.87e-05 mcm2l1d_cc_w_0_170_s_0_270=4.68e-11 mcm2l1d_cf_w_0_170_s_0_270=1.08e-11
+  mcm2l1d_ca_w_0_170_s_0_360=7.87e-05 mcm2l1d_cc_w_0_170_s_0_360=3.69e-11 mcm2l1d_cf_w_0_170_s_0_360=1.39e-11
+  mcm2l1d_ca_w_0_170_s_0_450=7.87e-05 mcm2l1d_cc_w_0_170_s_0_450=3.02e-11 mcm2l1d_cf_w_0_170_s_0_450=1.64e-11
+  mcm2l1d_ca_w_0_170_s_0_540=7.87e-05 mcm2l1d_cc_w_0_170_s_0_540=2.50e-11 mcm2l1d_cf_w_0_170_s_0_540=1.89e-11
+  mcm2l1d_ca_w_0_170_s_0_720=7.87e-05 mcm2l1d_cc_w_0_170_s_0_720=1.78e-11 mcm2l1d_cf_w_0_170_s_0_720=2.30e-11
+  mcm2l1d_ca_w_0_170_s_1_080=7.87e-05 mcm2l1d_cc_w_0_170_s_1_080=9.61e-12 mcm2l1d_cf_w_0_170_s_1_080=2.89e-11
+  mcm2l1d_ca_w_0_170_s_1_980=7.87e-05 mcm2l1d_cc_w_0_170_s_1_980=2.27e-12 mcm2l1d_cf_w_0_170_s_1_980=3.52e-11
+  mcm2l1d_ca_w_0_170_s_4_500=7.87e-05 mcm2l1d_cc_w_0_170_s_4_500=7.50e-14 mcm2l1d_cf_w_0_170_s_4_500=3.74e-11
+  mcm2l1d_ca_w_1_360_s_0_180=7.87e-05 mcm2l1d_cc_w_1_360_s_0_180=7.20e-11 mcm2l1d_cf_w_1_360_s_0_180=7.70e-12
+  mcm2l1d_ca_w_1_360_s_0_225=7.87e-05 mcm2l1d_cc_w_1_360_s_0_225=6.19e-11 mcm2l1d_cf_w_1_360_s_0_225=9.31e-12
+  mcm2l1d_ca_w_1_360_s_0_270=7.87e-05 mcm2l1d_cc_w_1_360_s_0_270=5.41e-11 mcm2l1d_cf_w_1_360_s_0_270=1.09e-11
+  mcm2l1d_ca_w_1_360_s_0_360=7.87e-05 mcm2l1d_cc_w_1_360_s_0_360=4.30e-11 mcm2l1d_cf_w_1_360_s_0_360=1.38e-11
+  mcm2l1d_ca_w_1_360_s_0_450=7.87e-05 mcm2l1d_cc_w_1_360_s_0_450=3.52e-11 mcm2l1d_cf_w_1_360_s_0_450=1.66e-11
+  mcm2l1d_ca_w_1_360_s_0_540=7.87e-05 mcm2l1d_cc_w_1_360_s_0_540=2.94e-11 mcm2l1d_cf_w_1_360_s_0_540=1.91e-11
+  mcm2l1d_ca_w_1_360_s_0_720=7.87e-05 mcm2l1d_cc_w_1_360_s_0_720=2.11e-11 mcm2l1d_cf_w_1_360_s_0_720=2.36e-11
+  mcm2l1d_ca_w_1_360_s_1_080=7.87e-05 mcm2l1d_cc_w_1_360_s_1_080=1.15e-11 mcm2l1d_cf_w_1_360_s_1_080=3.01e-11
+  mcm2l1d_ca_w_1_360_s_1_980=7.87e-05 mcm2l1d_cc_w_1_360_s_1_980=2.80e-12 mcm2l1d_cf_w_1_360_s_1_980=3.76e-11
+  mcm2l1d_ca_w_1_360_s_4_500=7.87e-05 mcm2l1d_cc_w_1_360_s_4_500=1.00e-13 mcm2l1d_cf_w_1_360_s_4_500=4.02e-11
+  mcm2l1p1_ca_w_0_170_s_0_180=1.02e-04 mcm2l1p1_cc_w_0_170_s_0_180=5.98e-11 mcm2l1p1_cf_w_0_170_s_0_180=9.88e-12
+  mcm2l1p1_ca_w_0_170_s_0_225=1.02e-04 mcm2l1p1_cc_w_0_170_s_0_225=5.06e-11 mcm2l1p1_cf_w_0_170_s_0_225=1.19e-11
+  mcm2l1p1_ca_w_0_170_s_0_270=1.02e-04 mcm2l1p1_cc_w_0_170_s_0_270=4.37e-11 mcm2l1p1_cf_w_0_170_s_0_270=1.38e-11
+  mcm2l1p1_ca_w_0_170_s_0_360=1.02e-04 mcm2l1p1_cc_w_0_170_s_0_360=3.37e-11 mcm2l1p1_cf_w_0_170_s_0_360=1.75e-11
+  mcm2l1p1_ca_w_0_170_s_0_450=1.02e-04 mcm2l1p1_cc_w_0_170_s_0_450=2.70e-11 mcm2l1p1_cf_w_0_170_s_0_450=2.05e-11
+  mcm2l1p1_ca_w_0_170_s_0_540=1.02e-04 mcm2l1p1_cc_w_0_170_s_0_540=2.18e-11 mcm2l1p1_cf_w_0_170_s_0_540=2.33e-11
+  mcm2l1p1_ca_w_0_170_s_0_720=1.02e-04 mcm2l1p1_cc_w_0_170_s_0_720=1.48e-11 mcm2l1p1_cf_w_0_170_s_0_720=2.79e-11
+  mcm2l1p1_ca_w_0_170_s_1_080=1.02e-04 mcm2l1p1_cc_w_0_170_s_1_080=7.22e-12 mcm2l1p1_cf_w_0_170_s_1_080=3.38e-11
+  mcm2l1p1_ca_w_0_170_s_1_980=1.02e-04 mcm2l1p1_cc_w_0_170_s_1_980=1.37e-12 mcm2l1p1_cf_w_0_170_s_1_980=3.91e-11
+  mcm2l1p1_ca_w_0_170_s_4_500=1.02e-04 mcm2l1p1_cc_w_0_170_s_4_500=4.00e-14 mcm2l1p1_cf_w_0_170_s_4_500=4.04e-11
+  mcm2l1p1_ca_w_1_360_s_0_180=1.02e-04 mcm2l1p1_cc_w_1_360_s_0_180=6.77e-11 mcm2l1p1_cf_w_1_360_s_0_180=9.85e-12
+  mcm2l1p1_ca_w_1_360_s_0_225=1.02e-04 mcm2l1p1_cc_w_1_360_s_0_225=5.75e-11 mcm2l1p1_cf_w_1_360_s_0_225=1.19e-11
+  mcm2l1p1_ca_w_1_360_s_0_270=1.02e-04 mcm2l1p1_cc_w_1_360_s_0_270=4.98e-11 mcm2l1p1_cf_w_1_360_s_0_270=1.38e-11
+  mcm2l1p1_ca_w_1_360_s_0_360=1.02e-04 mcm2l1p1_cc_w_1_360_s_0_360=3.88e-11 mcm2l1p1_cf_w_1_360_s_0_360=1.74e-11
+  mcm2l1p1_ca_w_1_360_s_0_450=1.02e-04 mcm2l1p1_cc_w_1_360_s_0_450=3.11e-11 mcm2l1p1_cf_w_1_360_s_0_450=2.07e-11
+  mcm2l1p1_ca_w_1_360_s_0_540=1.02e-04 mcm2l1p1_cc_w_1_360_s_0_540=2.54e-11 mcm2l1p1_cf_w_1_360_s_0_540=2.37e-11
+  mcm2l1p1_ca_w_1_360_s_0_720=1.02e-04 mcm2l1p1_cc_w_1_360_s_0_720=1.75e-11 mcm2l1p1_cf_w_1_360_s_0_720=2.86e-11
+  mcm2l1p1_ca_w_1_360_s_1_080=1.02e-04 mcm2l1p1_cc_w_1_360_s_1_080=8.81e-12 mcm2l1p1_cf_w_1_360_s_1_080=3.52e-11
+  mcm2l1p1_ca_w_1_360_s_1_980=1.02e-04 mcm2l1p1_cc_w_1_360_s_1_980=1.72e-12 mcm2l1p1_cf_w_1_360_s_1_980=4.16e-11
+  mcm2l1p1_ca_w_1_360_s_4_500=1.02e-04 mcm2l1p1_cc_w_1_360_s_4_500=5.00e-14 mcm2l1p1_cf_w_1_360_s_4_500=4.32e-11
+  mcm3l1f_ca_w_0_170_s_0_180=4.86e-05 mcm3l1f_cc_w_0_170_s_0_180=6.69e-11 mcm3l1f_cf_w_0_170_s_0_180=4.84e-12
+  mcm3l1f_ca_w_0_170_s_0_225=4.86e-05 mcm3l1f_cc_w_0_170_s_0_225=5.78e-11 mcm3l1f_cf_w_0_170_s_0_225=5.86e-12
+  mcm3l1f_ca_w_0_170_s_0_270=4.86e-05 mcm3l1f_cc_w_0_170_s_0_270=5.17e-11 mcm3l1f_cf_w_0_170_s_0_270=6.86e-12
+  mcm3l1f_ca_w_0_170_s_0_360=4.86e-05 mcm3l1f_cc_w_0_170_s_0_360=4.21e-11 mcm3l1f_cf_w_0_170_s_0_360=8.94e-12
+  mcm3l1f_ca_w_0_170_s_0_450=4.86e-05 mcm3l1f_cc_w_0_170_s_0_450=3.61e-11 mcm3l1f_cf_w_0_170_s_0_450=1.06e-11
+  mcm3l1f_ca_w_0_170_s_0_540=4.86e-05 mcm3l1f_cc_w_0_170_s_0_540=3.10e-11 mcm3l1f_cf_w_0_170_s_0_540=1.25e-11
+  mcm3l1f_ca_w_0_170_s_0_720=4.86e-05 mcm3l1f_cc_w_0_170_s_0_720=2.41e-11 mcm3l1f_cf_w_0_170_s_0_720=1.56e-11
+  mcm3l1f_ca_w_0_170_s_1_080=4.86e-05 mcm3l1f_cc_w_0_170_s_1_080=1.54e-11 mcm3l1f_cf_w_0_170_s_1_080=2.06e-11
+  mcm3l1f_ca_w_0_170_s_1_980=4.86e-05 mcm3l1f_cc_w_0_170_s_1_980=5.82e-12 mcm3l1f_cf_w_0_170_s_1_980=2.79e-11
+  mcm3l1f_ca_w_0_170_s_4_500=4.86e-05 mcm3l1f_cc_w_0_170_s_4_500=5.05e-13 mcm3l1f_cf_w_0_170_s_4_500=3.28e-11
+  mcm3l1f_ca_w_1_360_s_0_180=4.86e-05 mcm3l1f_cc_w_1_360_s_0_180=8.22e-11 mcm3l1f_cf_w_1_360_s_0_180=4.82e-12
+  mcm3l1f_ca_w_1_360_s_0_225=4.86e-05 mcm3l1f_cc_w_1_360_s_0_225=7.19e-11 mcm3l1f_cf_w_1_360_s_0_225=5.85e-12
+  mcm3l1f_ca_w_1_360_s_0_270=4.86e-05 mcm3l1f_cc_w_1_360_s_0_270=6.42e-11 mcm3l1f_cf_w_1_360_s_0_270=6.86e-12
+  mcm3l1f_ca_w_1_360_s_0_360=4.86e-05 mcm3l1f_cc_w_1_360_s_0_360=5.31e-11 mcm3l1f_cf_w_1_360_s_0_360=8.83e-12
+  mcm3l1f_ca_w_1_360_s_0_450=4.86e-05 mcm3l1f_cc_w_1_360_s_0_450=4.53e-11 mcm3l1f_cf_w_1_360_s_0_450=1.07e-11
+  mcm3l1f_ca_w_1_360_s_0_540=4.86e-05 mcm3l1f_cc_w_1_360_s_0_540=3.93e-11 mcm3l1f_cf_w_1_360_s_0_540=1.25e-11
+  mcm3l1f_ca_w_1_360_s_0_720=4.86e-05 mcm3l1f_cc_w_1_360_s_0_720=3.07e-11 mcm3l1f_cf_w_1_360_s_0_720=1.58e-11
+  mcm3l1f_ca_w_1_360_s_1_080=4.86e-05 mcm3l1f_cc_w_1_360_s_1_080=2.00e-11 mcm3l1f_cf_w_1_360_s_1_080=2.14e-11
+  mcm3l1f_ca_w_1_360_s_1_980=4.86e-05 mcm3l1f_cc_w_1_360_s_1_980=7.90e-12 mcm3l1f_cf_w_1_360_s_1_980=3.02e-11
+  mcm3l1f_ca_w_1_360_s_4_500=4.86e-05 mcm3l1f_cc_w_1_360_s_4_500=7.10e-13 mcm3l1f_cf_w_1_360_s_4_500=3.67e-11
+  mcm3l1d_ca_w_0_170_s_0_180=6.51e-05 mcm3l1d_cc_w_0_170_s_0_180=6.46e-11 mcm3l1d_cf_w_0_170_s_0_180=6.43e-12
+  mcm3l1d_ca_w_0_170_s_0_225=6.51e-05 mcm3l1d_cc_w_0_170_s_0_225=5.56e-11 mcm3l1d_cf_w_0_170_s_0_225=7.78e-12
+  mcm3l1d_ca_w_0_170_s_0_270=6.51e-05 mcm3l1d_cc_w_0_170_s_0_270=4.91e-11 mcm3l1d_cf_w_0_170_s_0_270=9.05e-12
+  mcm3l1d_ca_w_0_170_s_0_360=6.51e-05 mcm3l1d_cc_w_0_170_s_0_360=3.94e-11 mcm3l1d_cf_w_0_170_s_0_360=1.17e-11
+  mcm3l1d_ca_w_0_170_s_0_450=6.51e-05 mcm3l1d_cc_w_0_170_s_0_450=3.30e-11 mcm3l1d_cf_w_0_170_s_0_450=1.38e-11
+  mcm3l1d_ca_w_0_170_s_0_540=6.51e-05 mcm3l1d_cc_w_0_170_s_0_540=2.79e-11 mcm3l1d_cf_w_0_170_s_0_540=1.61e-11
+  mcm3l1d_ca_w_0_170_s_0_720=6.51e-05 mcm3l1d_cc_w_0_170_s_0_720=2.08e-11 mcm3l1d_cf_w_0_170_s_0_720=1.98e-11
+  mcm3l1d_ca_w_0_170_s_1_080=6.51e-05 mcm3l1d_cc_w_0_170_s_1_080=1.24e-11 mcm3l1d_cf_w_0_170_s_1_080=2.54e-11
+  mcm3l1d_ca_w_0_170_s_1_980=6.51e-05 mcm3l1d_cc_w_0_170_s_1_980=3.94e-12 mcm3l1d_cf_w_0_170_s_1_980=3.24e-11
+  mcm3l1d_ca_w_0_170_s_4_500=6.51e-05 mcm3l1d_cc_w_0_170_s_4_500=2.55e-13 mcm3l1d_cf_w_0_170_s_4_500=3.59e-11
+  mcm3l1d_ca_w_1_360_s_0_180=6.51e-05 mcm3l1d_cc_w_1_360_s_0_180=7.76e-11 mcm3l1d_cf_w_1_360_s_0_180=6.41e-12
+  mcm3l1d_ca_w_1_360_s_0_225=6.51e-05 mcm3l1d_cc_w_1_360_s_0_225=6.74e-11 mcm3l1d_cf_w_1_360_s_0_225=7.76e-12
+  mcm3l1d_ca_w_1_360_s_0_270=6.51e-05 mcm3l1d_cc_w_1_360_s_0_270=5.96e-11 mcm3l1d_cf_w_1_360_s_0_270=9.08e-12
+  mcm3l1d_ca_w_1_360_s_0_360=6.51e-05 mcm3l1d_cc_w_1_360_s_0_360=4.86e-11 mcm3l1d_cf_w_1_360_s_0_360=1.16e-11
+  mcm3l1d_ca_w_1_360_s_0_450=6.51e-05 mcm3l1d_cc_w_1_360_s_0_450=4.08e-11 mcm3l1d_cf_w_1_360_s_0_450=1.40e-11
+  mcm3l1d_ca_w_1_360_s_0_540=6.51e-05 mcm3l1d_cc_w_1_360_s_0_540=3.49e-11 mcm3l1d_cf_w_1_360_s_0_540=1.62e-11
+  mcm3l1d_ca_w_1_360_s_0_720=6.51e-05 mcm3l1d_cc_w_1_360_s_0_720=2.64e-11 mcm3l1d_cf_w_1_360_s_0_720=2.02e-11
+  mcm3l1d_ca_w_1_360_s_1_080=6.51e-05 mcm3l1d_cc_w_1_360_s_1_080=1.63e-11 mcm3l1d_cf_w_1_360_s_1_080=2.65e-11
+  mcm3l1d_ca_w_1_360_s_1_980=6.51e-05 mcm3l1d_cc_w_1_360_s_1_980=5.49e-12 mcm3l1d_cf_w_1_360_s_1_980=3.51e-11
+  mcm3l1d_ca_w_1_360_s_4_500=6.51e-05 mcm3l1d_cc_w_1_360_s_4_500=3.35e-13 mcm3l1d_cf_w_1_360_s_4_500=3.99e-11
+  mcm3l1p1_ca_w_0_170_s_0_180=8.83e-05 mcm3l1p1_cc_w_0_170_s_0_180=6.19e-11 mcm3l1p1_cf_w_0_170_s_0_180=8.62e-12
+  mcm3l1p1_ca_w_0_170_s_0_225=8.83e-05 mcm3l1p1_cc_w_0_170_s_0_225=5.26e-11 mcm3l1p1_cf_w_0_170_s_0_225=1.04e-11
+  mcm3l1p1_ca_w_0_170_s_0_270=8.83e-05 mcm3l1p1_cc_w_0_170_s_0_270=4.60e-11 mcm3l1p1_cf_w_0_170_s_0_270=1.20e-11
+  mcm3l1p1_ca_w_0_170_s_0_360=8.83e-05 mcm3l1p1_cc_w_0_170_s_0_360=3.61e-11 mcm3l1p1_cf_w_0_170_s_0_360=1.54e-11
+  mcm3l1p1_ca_w_0_170_s_0_450=8.83e-05 mcm3l1p1_cc_w_0_170_s_0_450=2.97e-11 mcm3l1p1_cf_w_0_170_s_0_450=1.81e-11
+  mcm3l1p1_ca_w_0_170_s_0_540=8.83e-05 mcm3l1p1_cc_w_0_170_s_0_540=2.44e-11 mcm3l1p1_cf_w_0_170_s_0_540=2.08e-11
+  mcm3l1p1_ca_w_0_170_s_0_720=8.83e-05 mcm3l1p1_cc_w_0_170_s_0_720=1.75e-11 mcm3l1p1_cf_w_0_170_s_0_720=2.51e-11
+  mcm3l1p1_ca_w_0_170_s_1_080=8.83e-05 mcm3l1p1_cc_w_0_170_s_1_080=9.59e-12 mcm3l1p1_cf_w_0_170_s_1_080=3.10e-11
+  mcm3l1p1_ca_w_0_170_s_1_980=8.83e-05 mcm3l1p1_cc_w_0_170_s_1_980=2.63e-12 mcm3l1p1_cf_w_0_170_s_1_980=3.71e-11
+  mcm3l1p1_ca_w_0_170_s_4_500=8.83e-05 mcm3l1p1_cc_w_0_170_s_4_500=1.45e-13 mcm3l1p1_cf_w_0_170_s_4_500=3.95e-11
+  mcm3l1p1_ca_w_1_360_s_0_180=8.83e-05 mcm3l1p1_cc_w_1_360_s_0_180=7.32e-11 mcm3l1p1_cf_w_1_360_s_0_180=8.62e-12
+  mcm3l1p1_ca_w_1_360_s_0_225=8.83e-05 mcm3l1p1_cc_w_1_360_s_0_225=6.31e-11 mcm3l1p1_cf_w_1_360_s_0_225=1.04e-11
+  mcm3l1p1_ca_w_1_360_s_0_270=8.83e-05 mcm3l1p1_cc_w_1_360_s_0_270=5.53e-11 mcm3l1p1_cf_w_1_360_s_0_270=1.21e-11
+  mcm3l1p1_ca_w_1_360_s_0_360=8.83e-05 mcm3l1p1_cc_w_1_360_s_0_360=4.42e-11 mcm3l1p1_cf_w_1_360_s_0_360=1.53e-11
+  mcm3l1p1_ca_w_1_360_s_0_450=8.83e-05 mcm3l1p1_cc_w_1_360_s_0_450=3.66e-11 mcm3l1p1_cf_w_1_360_s_0_450=1.83e-11
+  mcm3l1p1_ca_w_1_360_s_0_540=8.83e-05 mcm3l1p1_cc_w_1_360_s_0_540=3.08e-11 mcm3l1p1_cf_w_1_360_s_0_540=2.10e-11
+  mcm3l1p1_ca_w_1_360_s_0_720=8.83e-05 mcm3l1p1_cc_w_1_360_s_0_720=2.26e-11 mcm3l1p1_cf_w_1_360_s_0_720=2.56e-11
+  mcm3l1p1_ca_w_1_360_s_1_080=8.83e-05 mcm3l1p1_cc_w_1_360_s_1_080=1.31e-11 mcm3l1p1_cf_w_1_360_s_1_080=3.24e-11
+  mcm3l1p1_ca_w_1_360_s_1_980=8.83e-05 mcm3l1p1_cc_w_1_360_s_1_980=3.86e-12 mcm3l1p1_cf_w_1_360_s_1_980=4.03e-11
+  mcm3l1p1_ca_w_1_360_s_4_500=8.83e-05 mcm3l1p1_cc_w_1_360_s_4_500=2.55e-13 mcm3l1p1_cf_w_1_360_s_4_500=4.38e-11
+  mcm4l1f_ca_w_0_170_s_0_180=4.16e-05 mcm4l1f_cc_w_0_170_s_0_180=6.79e-11 mcm4l1f_cf_w_0_170_s_0_180=4.16e-12
+  mcm4l1f_ca_w_0_170_s_0_225=4.16e-05 mcm4l1f_cc_w_0_170_s_0_225=5.89e-11 mcm4l1f_cf_w_0_170_s_0_225=5.03e-12
+  mcm4l1f_ca_w_0_170_s_0_270=4.16e-05 mcm4l1f_cc_w_0_170_s_0_270=5.29e-11 mcm4l1f_cf_w_0_170_s_0_270=5.90e-12
+  mcm4l1f_ca_w_0_170_s_0_360=4.16e-05 mcm4l1f_cc_w_0_170_s_0_360=4.36e-11 mcm4l1f_cf_w_0_170_s_0_360=7.74e-12
+  mcm4l1f_ca_w_0_170_s_0_450=4.16e-05 mcm4l1f_cc_w_0_170_s_0_450=3.77e-11 mcm4l1f_cf_w_0_170_s_0_450=9.18e-12
+  mcm4l1f_ca_w_0_170_s_0_540=4.16e-05 mcm4l1f_cc_w_0_170_s_0_540=3.27e-11 mcm4l1f_cf_w_0_170_s_0_540=1.09e-11
+  mcm4l1f_ca_w_0_170_s_0_720=4.16e-05 mcm4l1f_cc_w_0_170_s_0_720=2.59e-11 mcm4l1f_cf_w_0_170_s_0_720=1.37e-11
+  mcm4l1f_ca_w_0_170_s_1_080=4.16e-05 mcm4l1f_cc_w_0_170_s_1_080=1.75e-11 mcm4l1f_cf_w_0_170_s_1_080=1.83e-11
+  mcm4l1f_ca_w_0_170_s_1_980=4.16e-05 mcm4l1f_cc_w_0_170_s_1_980=7.68e-12 mcm4l1f_cf_w_0_170_s_1_980=2.55e-11
+  mcm4l1f_ca_w_0_170_s_4_500=4.16e-05 mcm4l1f_cc_w_0_170_s_4_500=1.10e-12 mcm4l1f_cf_w_0_170_s_4_500=3.13e-11
+  mcm4l1f_ca_w_1_360_s_0_180=4.16e-05 mcm4l1f_cc_w_1_360_s_0_180=8.59e-11 mcm4l1f_cf_w_1_360_s_0_180=4.15e-12
+  mcm4l1f_ca_w_1_360_s_0_225=4.16e-05 mcm4l1f_cc_w_1_360_s_0_225=7.57e-11 mcm4l1f_cf_w_1_360_s_0_225=5.03e-12
+  mcm4l1f_ca_w_1_360_s_0_270=4.16e-05 mcm4l1f_cc_w_1_360_s_0_270=6.80e-11 mcm4l1f_cf_w_1_360_s_0_270=5.91e-12
+  mcm4l1f_ca_w_1_360_s_0_360=4.16e-05 mcm4l1f_cc_w_1_360_s_0_360=5.70e-11 mcm4l1f_cf_w_1_360_s_0_360=7.62e-12
+  mcm4l1f_ca_w_1_360_s_0_450=4.16e-05 mcm4l1f_cc_w_1_360_s_0_450=4.93e-11 mcm4l1f_cf_w_1_360_s_0_450=9.27e-12
+  mcm4l1f_ca_w_1_360_s_0_540=4.16e-05 mcm4l1f_cc_w_1_360_s_0_540=4.34e-11 mcm4l1f_cf_w_1_360_s_0_540=1.08e-11
+  mcm4l1f_ca_w_1_360_s_0_720=4.16e-05 mcm4l1f_cc_w_1_360_s_0_720=3.48e-11 mcm4l1f_cf_w_1_360_s_0_720=1.38e-11
+  mcm4l1f_ca_w_1_360_s_1_080=4.16e-05 mcm4l1f_cc_w_1_360_s_1_080=2.41e-11 mcm4l1f_cf_w_1_360_s_1_080=1.89e-11
+  mcm4l1f_ca_w_1_360_s_1_980=4.16e-05 mcm4l1f_cc_w_1_360_s_1_980=1.11e-11 mcm4l1f_cf_w_1_360_s_1_980=2.76e-11
+  mcm4l1f_ca_w_1_360_s_4_500=4.16e-05 mcm4l1f_cc_w_1_360_s_4_500=1.73e-12 mcm4l1f_cf_w_1_360_s_4_500=3.58e-11
+  mcm4l1d_ca_w_0_170_s_0_180=5.81e-05 mcm4l1d_cc_w_0_170_s_0_180=6.56e-11 mcm4l1d_cf_w_0_170_s_0_180=5.75e-12
+  mcm4l1d_ca_w_0_170_s_0_225=5.81e-05 mcm4l1d_cc_w_0_170_s_0_225=5.66e-11 mcm4l1d_cf_w_0_170_s_0_225=6.96e-12
+  mcm4l1d_ca_w_0_170_s_0_270=5.81e-05 mcm4l1d_cc_w_0_170_s_0_270=5.04e-11 mcm4l1d_cf_w_0_170_s_0_270=8.11e-12
+  mcm4l1d_ca_w_0_170_s_0_360=5.81e-05 mcm4l1d_cc_w_0_170_s_0_360=4.08e-11 mcm4l1d_cf_w_0_170_s_0_360=1.05e-11
+  mcm4l1d_ca_w_0_170_s_0_450=5.81e-05 mcm4l1d_cc_w_0_170_s_0_450=3.46e-11 mcm4l1d_cf_w_0_170_s_0_450=1.25e-11
+  mcm4l1d_ca_w_0_170_s_0_540=5.81e-05 mcm4l1d_cc_w_0_170_s_0_540=2.95e-11 mcm4l1d_cf_w_0_170_s_0_540=1.46e-11
+  mcm4l1d_ca_w_0_170_s_0_720=5.81e-05 mcm4l1d_cc_w_0_170_s_0_720=2.26e-11 mcm4l1d_cf_w_0_170_s_0_720=1.81e-11
+  mcm4l1d_ca_w_0_170_s_1_080=5.81e-05 mcm4l1d_cc_w_0_170_s_1_080=1.42e-11 mcm4l1d_cf_w_0_170_s_1_080=2.35e-11
+  mcm4l1d_ca_w_0_170_s_1_980=5.81e-05 mcm4l1d_cc_w_0_170_s_1_980=5.39e-12 mcm4l1d_cf_w_0_170_s_1_980=3.06e-11
+  mcm4l1d_ca_w_0_170_s_4_500=5.81e-05 mcm4l1d_cc_w_0_170_s_4_500=6.20e-13 mcm4l1d_cf_w_0_170_s_4_500=3.50e-11
+  mcm4l1d_ca_w_1_360_s_0_180=5.81e-05 mcm4l1d_cc_w_1_360_s_0_180=8.13e-11 mcm4l1d_cf_w_1_360_s_0_180=5.74e-12
+  mcm4l1d_ca_w_1_360_s_0_225=5.81e-05 mcm4l1d_cc_w_1_360_s_0_225=7.11e-11 mcm4l1d_cf_w_1_360_s_0_225=6.94e-12
+  mcm4l1d_ca_w_1_360_s_0_270=5.81e-05 mcm4l1d_cc_w_1_360_s_0_270=6.35e-11 mcm4l1d_cf_w_1_360_s_0_270=8.13e-12
+  mcm4l1d_ca_w_1_360_s_0_360=5.81e-05 mcm4l1d_cc_w_1_360_s_0_360=5.24e-11 mcm4l1d_cf_w_1_360_s_0_360=1.04e-11
+  mcm4l1d_ca_w_1_360_s_0_450=5.81e-05 mcm4l1d_cc_w_1_360_s_0_450=4.47e-11 mcm4l1d_cf_w_1_360_s_0_450=1.26e-11
+  mcm4l1d_ca_w_1_360_s_0_540=5.81e-05 mcm4l1d_cc_w_1_360_s_0_540=3.89e-11 mcm4l1d_cf_w_1_360_s_0_540=1.46e-11
+  mcm4l1d_ca_w_1_360_s_0_720=5.81e-05 mcm4l1d_cc_w_1_360_s_0_720=3.04e-11 mcm4l1d_cf_w_1_360_s_0_720=1.83e-11
+  mcm4l1d_ca_w_1_360_s_1_080=5.81e-05 mcm4l1d_cc_w_1_360_s_1_080=2.00e-11 mcm4l1d_cf_w_1_360_s_1_080=2.44e-11
+  mcm4l1d_ca_w_1_360_s_1_980=5.81e-05 mcm4l1d_cc_w_1_360_s_1_980=8.35e-12 mcm4l1d_cf_w_1_360_s_1_980=3.33e-11
+  mcm4l1d_ca_w_1_360_s_4_500=5.81e-05 mcm4l1d_cc_w_1_360_s_4_500=1.07e-12 mcm4l1d_cf_w_1_360_s_4_500=4.00e-11
+  mcm4l1p1_ca_w_0_170_s_0_180=8.13e-05 mcm4l1p1_cc_w_0_170_s_0_180=6.27e-11 mcm4l1p1_cf_w_0_170_s_0_180=7.94e-12
+  mcm4l1p1_ca_w_0_170_s_0_225=8.13e-05 mcm4l1p1_cc_w_0_170_s_0_225=5.36e-11 mcm4l1p1_cf_w_0_170_s_0_225=9.56e-12
+  mcm4l1p1_ca_w_0_170_s_0_270=8.13e-05 mcm4l1p1_cc_w_0_170_s_0_270=4.72e-11 mcm4l1p1_cf_w_0_170_s_0_270=1.11e-11
+  mcm4l1p1_ca_w_0_170_s_0_360=8.13e-05 mcm4l1p1_cc_w_0_170_s_0_360=3.74e-11 mcm4l1p1_cf_w_0_170_s_0_360=1.43e-11
+  mcm4l1p1_ca_w_0_170_s_0_450=8.13e-05 mcm4l1p1_cc_w_0_170_s_0_450=3.12e-11 mcm4l1p1_cf_w_0_170_s_0_450=1.67e-11
+  mcm4l1p1_ca_w_0_170_s_0_540=8.13e-05 mcm4l1p1_cc_w_0_170_s_0_540=2.60e-11 mcm4l1p1_cf_w_0_170_s_0_540=1.94e-11
+  mcm4l1p1_ca_w_0_170_s_0_720=8.13e-05 mcm4l1p1_cc_w_0_170_s_0_720=1.91e-11 mcm4l1p1_cf_w_0_170_s_0_720=2.36e-11
+  mcm4l1p1_ca_w_0_170_s_1_080=8.13e-05 mcm4l1p1_cc_w_0_170_s_1_080=1.11e-11 mcm4l1p1_cf_w_0_170_s_1_080=2.94e-11
+  mcm4l1p1_ca_w_0_170_s_1_980=8.13e-05 mcm4l1p1_cc_w_0_170_s_1_980=3.73e-12 mcm4l1p1_cf_w_0_170_s_1_980=3.59e-11
+  mcm4l1p1_ca_w_0_170_s_4_500=8.13e-05 mcm4l1p1_cc_w_0_170_s_4_500=3.70e-13 mcm4l1p1_cf_w_0_170_s_4_500=3.90e-11
+  mcm4l1p1_ca_w_1_360_s_0_180=8.13e-05 mcm4l1p1_cc_w_1_360_s_0_180=7.68e-11 mcm4l1p1_cf_w_1_360_s_0_180=7.98e-12
+  mcm4l1p1_ca_w_1_360_s_0_225=8.13e-05 mcm4l1p1_cc_w_1_360_s_0_225=6.68e-11 mcm4l1p1_cf_w_1_360_s_0_225=9.62e-12
+  mcm4l1p1_ca_w_1_360_s_0_270=8.13e-05 mcm4l1p1_cc_w_1_360_s_0_270=5.91e-11 mcm4l1p1_cf_w_1_360_s_0_270=1.12e-11
+  mcm4l1p1_ca_w_1_360_s_0_360=8.13e-05 mcm4l1p1_cc_w_1_360_s_0_360=4.82e-11 mcm4l1p1_cf_w_1_360_s_0_360=1.42e-11
+  mcm4l1p1_ca_w_1_360_s_0_450=8.13e-05 mcm4l1p1_cc_w_1_360_s_0_450=4.04e-11 mcm4l1p1_cf_w_1_360_s_0_450=1.70e-11
+  mcm4l1p1_ca_w_1_360_s_0_540=8.13e-05 mcm4l1p1_cc_w_1_360_s_0_540=3.47e-11 mcm4l1p1_cf_w_1_360_s_0_540=1.95e-11
+  mcm4l1p1_ca_w_1_360_s_0_720=8.13e-05 mcm4l1p1_cc_w_1_360_s_0_720=2.65e-11 mcm4l1p1_cf_w_1_360_s_0_720=2.40e-11
+  mcm4l1p1_ca_w_1_360_s_1_080=8.13e-05 mcm4l1p1_cc_w_1_360_s_1_080=1.66e-11 mcm4l1p1_cf_w_1_360_s_1_080=3.06e-11
+  mcm4l1p1_ca_w_1_360_s_1_980=8.13e-05 mcm4l1p1_cc_w_1_360_s_1_980=6.33e-12 mcm4l1p1_cf_w_1_360_s_1_980=3.93e-11
+  mcm4l1p1_ca_w_1_360_s_4_500=8.13e-05 mcm4l1p1_cc_w_1_360_s_4_500=7.25e-13 mcm4l1p1_cf_w_1_360_s_4_500=4.46e-11
+  mcm5l1f_ca_w_0_170_s_0_180=3.85e-05 mcm5l1f_cc_w_0_170_s_0_180=6.83e-11 mcm5l1f_cf_w_0_170_s_0_180=3.85e-12
+  mcm5l1f_ca_w_0_170_s_0_225=3.85e-05 mcm5l1f_cc_w_0_170_s_0_225=5.93e-11 mcm5l1f_cf_w_0_170_s_0_225=4.65e-12
+  mcm5l1f_ca_w_0_170_s_0_270=3.85e-05 mcm5l1f_cc_w_0_170_s_0_270=5.35e-11 mcm5l1f_cf_w_0_170_s_0_270=5.46e-12
+  mcm5l1f_ca_w_0_170_s_0_360=3.85e-05 mcm5l1f_cc_w_0_170_s_0_360=4.42e-11 mcm5l1f_cf_w_0_170_s_0_360=7.18e-12
+  mcm5l1f_ca_w_0_170_s_0_450=3.85e-05 mcm5l1f_cc_w_0_170_s_0_450=3.85e-11 mcm5l1f_cf_w_0_170_s_0_450=8.51e-12
+  mcm5l1f_ca_w_0_170_s_0_540=3.85e-05 mcm5l1f_cc_w_0_170_s_0_540=3.35e-11 mcm5l1f_cf_w_0_170_s_0_540=1.01e-11
+  mcm5l1f_ca_w_0_170_s_0_720=3.85e-05 mcm5l1f_cc_w_0_170_s_0_720=2.69e-11 mcm5l1f_cf_w_0_170_s_0_720=1.28e-11
+  mcm5l1f_ca_w_0_170_s_1_080=3.85e-05 mcm5l1f_cc_w_0_170_s_1_080=1.86e-11 mcm5l1f_cf_w_0_170_s_1_080=1.73e-11
+  mcm5l1f_ca_w_0_170_s_1_980=3.85e-05 mcm5l1f_cc_w_0_170_s_1_980=8.77e-12 mcm5l1f_cf_w_0_170_s_1_980=2.42e-11
+  mcm5l1f_ca_w_0_170_s_4_500=3.85e-05 mcm5l1f_cc_w_0_170_s_4_500=1.60e-12 mcm5l1f_cf_w_0_170_s_4_500=3.06e-11
+  mcm5l1f_ca_w_1_360_s_0_180=3.85e-05 mcm5l1f_cc_w_1_360_s_0_180=8.77e-11 mcm5l1f_cf_w_1_360_s_0_180=3.84e-12
+  mcm5l1f_ca_w_1_360_s_0_225=3.85e-05 mcm5l1f_cc_w_1_360_s_0_225=7.75e-11 mcm5l1f_cf_w_1_360_s_0_225=4.66e-12
+  mcm5l1f_ca_w_1_360_s_0_270=3.85e-05 mcm5l1f_cc_w_1_360_s_0_270=7.00e-11 mcm5l1f_cf_w_1_360_s_0_270=5.47e-12
+  mcm5l1f_ca_w_1_360_s_0_360=3.85e-05 mcm5l1f_cc_w_1_360_s_0_360=5.91e-11 mcm5l1f_cf_w_1_360_s_0_360=7.06e-12
+  mcm5l1f_ca_w_1_360_s_0_450=3.85e-05 mcm5l1f_cc_w_1_360_s_0_450=5.14e-11 mcm5l1f_cf_w_1_360_s_0_450=8.59e-12
+  mcm5l1f_ca_w_1_360_s_0_540=3.85e-05 mcm5l1f_cc_w_1_360_s_0_540=4.56e-11 mcm5l1f_cf_w_1_360_s_0_540=1.01e-11
+  mcm5l1f_ca_w_1_360_s_0_720=3.85e-05 mcm5l1f_cc_w_1_360_s_0_720=3.71e-11 mcm5l1f_cf_w_1_360_s_0_720=1.28e-11
+  mcm5l1f_ca_w_1_360_s_1_080=3.85e-05 mcm5l1f_cc_w_1_360_s_1_080=2.64e-11 mcm5l1f_cf_w_1_360_s_1_080=1.77e-11
+  mcm5l1f_ca_w_1_360_s_1_980=3.85e-05 mcm5l1f_cc_w_1_360_s_1_980=1.32e-11 mcm5l1f_cf_w_1_360_s_1_980=2.62e-11
+  mcm5l1f_ca_w_1_360_s_4_500=3.85e-05 mcm5l1f_cc_w_1_360_s_4_500=2.76e-12 mcm5l1f_cf_w_1_360_s_4_500=3.52e-11
+  mcm5l1d_ca_w_0_170_s_0_180=5.50e-05 mcm5l1d_cc_w_0_170_s_0_180=6.59e-11 mcm5l1d_cf_w_0_170_s_0_180=5.44e-12
+  mcm5l1d_ca_w_0_170_s_0_225=5.50e-05 mcm5l1d_cc_w_0_170_s_0_225=5.71e-11 mcm5l1d_cf_w_0_170_s_0_225=6.59e-12
+  mcm5l1d_ca_w_0_170_s_0_270=5.50e-05 mcm5l1d_cc_w_0_170_s_0_270=5.09e-11 mcm5l1d_cf_w_0_170_s_0_270=7.68e-12
+  mcm5l1d_ca_w_0_170_s_0_360=5.50e-05 mcm5l1d_cc_w_0_170_s_0_360=4.13e-11 mcm5l1d_cf_w_0_170_s_0_360=9.99e-12
+  mcm5l1d_ca_w_0_170_s_0_450=5.50e-05 mcm5l1d_cc_w_0_170_s_0_450=3.54e-11 mcm5l1d_cf_w_0_170_s_0_450=1.18e-11
+  mcm5l1d_ca_w_0_170_s_0_540=5.50e-05 mcm5l1d_cc_w_0_170_s_0_540=3.03e-11 mcm5l1d_cf_w_0_170_s_0_540=1.39e-11
+  mcm5l1d_ca_w_0_170_s_0_720=5.50e-05 mcm5l1d_cc_w_0_170_s_0_720=2.34e-11 mcm5l1d_cf_w_0_170_s_0_720=1.73e-11
+  mcm5l1d_ca_w_0_170_s_1_080=5.50e-05 mcm5l1d_cc_w_0_170_s_1_080=1.51e-11 mcm5l1d_cf_w_0_170_s_1_080=2.26e-11
+  mcm5l1d_ca_w_0_170_s_1_980=5.50e-05 mcm5l1d_cc_w_0_170_s_1_980=6.25e-12 mcm5l1d_cf_w_0_170_s_1_980=2.97e-11
+  mcm5l1d_ca_w_0_170_s_4_500=5.50e-05 mcm5l1d_cc_w_0_170_s_4_500=9.55e-13 mcm5l1d_cf_w_0_170_s_4_500=3.46e-11
+  mcm5l1d_ca_w_1_360_s_0_180=5.50e-05 mcm5l1d_cc_w_1_360_s_0_180=8.32e-11 mcm5l1d_cf_w_1_360_s_0_180=5.43e-12
+  mcm5l1d_ca_w_1_360_s_0_225=5.50e-05 mcm5l1d_cc_w_1_360_s_0_225=7.30e-11 mcm5l1d_cf_w_1_360_s_0_225=6.58e-12
+  mcm5l1d_ca_w_1_360_s_0_270=5.50e-05 mcm5l1d_cc_w_1_360_s_0_270=6.55e-11 mcm5l1d_cf_w_1_360_s_0_270=7.70e-12
+  mcm5l1d_ca_w_1_360_s_0_360=5.50e-05 mcm5l1d_cc_w_1_360_s_0_360=5.45e-11 mcm5l1d_cf_w_1_360_s_0_360=9.87e-12
+  mcm5l1d_ca_w_1_360_s_0_450=5.50e-05 mcm5l1d_cc_w_1_360_s_0_450=4.68e-11 mcm5l1d_cf_w_1_360_s_0_450=1.19e-11
+  mcm5l1d_ca_w_1_360_s_0_540=5.50e-05 mcm5l1d_cc_w_1_360_s_0_540=4.10e-11 mcm5l1d_cf_w_1_360_s_0_540=1.39e-11
+  mcm5l1d_ca_w_1_360_s_0_720=5.50e-05 mcm5l1d_cc_w_1_360_s_0_720=3.26e-11 mcm5l1d_cf_w_1_360_s_0_720=1.74e-11
+  mcm5l1d_ca_w_1_360_s_1_080=5.50e-05 mcm5l1d_cc_w_1_360_s_1_080=2.22e-11 mcm5l1d_cf_w_1_360_s_1_080=2.33e-11
+  mcm5l1d_ca_w_1_360_s_1_980=5.50e-05 mcm5l1d_cc_w_1_360_s_1_980=1.02e-11 mcm5l1d_cf_w_1_360_s_1_980=3.24e-11
+  mcm5l1d_ca_w_1_360_s_4_500=5.50e-05 mcm5l1d_cc_w_1_360_s_4_500=1.86e-12 mcm5l1d_cf_w_1_360_s_4_500=4.00e-11
+  mcm5l1p1_ca_w_0_170_s_0_180=7.81e-05 mcm5l1p1_cc_w_0_170_s_0_180=6.32e-11 mcm5l1p1_cf_w_0_170_s_0_180=7.63e-12
+  mcm5l1p1_ca_w_0_170_s_0_225=7.81e-05 mcm5l1p1_cc_w_0_170_s_0_225=5.41e-11 mcm5l1p1_cf_w_0_170_s_0_225=9.19e-12
+  mcm5l1p1_ca_w_0_170_s_0_270=7.81e-05 mcm5l1p1_cc_w_0_170_s_0_270=4.77e-11 mcm5l1p1_cf_w_0_170_s_0_270=1.07e-11
+  mcm5l1p1_ca_w_0_170_s_0_360=7.81e-05 mcm5l1p1_cc_w_0_170_s_0_360=3.80e-11 mcm5l1p1_cf_w_0_170_s_0_360=1.38e-11
+  mcm5l1p1_ca_w_0_170_s_0_450=7.81e-05 mcm5l1p1_cc_w_0_170_s_0_450=3.19e-11 mcm5l1p1_cf_w_0_170_s_0_450=1.61e-11
+  mcm5l1p1_ca_w_0_170_s_0_540=7.81e-05 mcm5l1p1_cc_w_0_170_s_0_540=2.67e-11 mcm5l1p1_cf_w_0_170_s_0_540=1.88e-11
+  mcm5l1p1_ca_w_0_170_s_0_720=7.81e-05 mcm5l1p1_cc_w_0_170_s_0_720=1.98e-11 mcm5l1p1_cf_w_0_170_s_0_720=2.28e-11
+  mcm5l1p1_ca_w_0_170_s_1_080=7.81e-05 mcm5l1p1_cc_w_0_170_s_1_080=1.19e-11 mcm5l1p1_cf_w_0_170_s_1_080=2.86e-11
+  mcm5l1p1_ca_w_0_170_s_1_980=7.81e-05 mcm5l1p1_cc_w_0_170_s_1_980=4.38e-12 mcm5l1p1_cf_w_0_170_s_1_980=3.52e-11
+  mcm5l1p1_ca_w_0_170_s_4_500=7.81e-05 mcm5l1p1_cc_w_0_170_s_4_500=5.96e-13 mcm5l1p1_cf_w_0_170_s_4_500=3.88e-11
+  mcm5l1p1_ca_w_1_360_s_0_180=7.81e-05 mcm5l1p1_cc_w_1_360_s_0_180=7.88e-11 mcm5l1p1_cf_w_1_360_s_0_180=7.69e-12
+  mcm5l1p1_ca_w_1_360_s_0_225=7.81e-05 mcm5l1p1_cc_w_1_360_s_0_225=6.87e-11 mcm5l1p1_cf_w_1_360_s_0_225=9.25e-12
+  mcm5l1p1_ca_w_1_360_s_0_270=7.81e-05 mcm5l1p1_cc_w_1_360_s_0_270=6.11e-11 mcm5l1p1_cf_w_1_360_s_0_270=1.08e-11
+  mcm5l1p1_ca_w_1_360_s_0_360=7.81e-05 mcm5l1p1_cc_w_1_360_s_0_360=5.02e-11 mcm5l1p1_cf_w_1_360_s_0_360=1.37e-11
+  mcm5l1p1_ca_w_1_360_s_0_450=7.81e-05 mcm5l1p1_cc_w_1_360_s_0_450=4.26e-11 mcm5l1p1_cf_w_1_360_s_0_450=1.64e-11
+  mcm5l1p1_ca_w_1_360_s_0_540=7.81e-05 mcm5l1p1_cc_w_1_360_s_0_540=3.68e-11 mcm5l1p1_cf_w_1_360_s_0_540=1.88e-11
+  mcm5l1p1_ca_w_1_360_s_0_720=7.81e-05 mcm5l1p1_cc_w_1_360_s_0_720=2.86e-11 mcm5l1p1_cf_w_1_360_s_0_720=2.32e-11
+  mcm5l1p1_ca_w_1_360_s_1_080=7.81e-05 mcm5l1p1_cc_w_1_360_s_1_080=1.87e-11 mcm5l1p1_cf_w_1_360_s_1_080=2.98e-11
+  mcm5l1p1_ca_w_1_360_s_1_980=7.81e-05 mcm5l1p1_cc_w_1_360_s_1_980=7.95e-12 mcm5l1p1_cf_w_1_360_s_1_980=3.87e-11
+  mcm5l1p1_ca_w_1_360_s_4_500=7.81e-05 mcm5l1p1_cc_w_1_360_s_4_500=1.34e-12 mcm5l1p1_cf_w_1_360_s_4_500=4.50e-11
+  mcrdll1f_ca_w_0_170_s_0_180=3.36e-05 mcrdll1f_cc_w_0_170_s_0_180=6.88e-11 mcrdll1f_cf_w_0_170_s_0_180=3.36e-12
+  mcrdll1f_ca_w_0_170_s_0_225=3.36e-05 mcrdll1f_cc_w_0_170_s_0_225=6.01e-11 mcrdll1f_cf_w_0_170_s_0_225=4.07e-12
+  mcrdll1f_ca_w_0_170_s_0_270=3.36e-05 mcrdll1f_cc_w_0_170_s_0_270=5.43e-11 mcrdll1f_cf_w_0_170_s_0_270=4.78e-12
+  mcrdll1f_ca_w_0_170_s_0_360=3.36e-05 mcrdll1f_cc_w_0_170_s_0_360=4.52e-11 mcrdll1f_cf_w_0_170_s_0_360=6.31e-12
+  mcrdll1f_ca_w_0_170_s_0_450=3.36e-05 mcrdll1f_cc_w_0_170_s_0_450=3.96e-11 mcrdll1f_cf_w_0_170_s_0_450=7.46e-12
+  mcrdll1f_ca_w_0_170_s_0_540=3.36e-05 mcrdll1f_cc_w_0_170_s_0_540=3.48e-11 mcrdll1f_cf_w_0_170_s_0_540=8.95e-12
+  mcrdll1f_ca_w_0_170_s_0_720=3.36e-05 mcrdll1f_cc_w_0_170_s_0_720=2.83e-11 mcrdll1f_cf_w_0_170_s_0_720=1.14e-11
+  mcrdll1f_ca_w_0_170_s_1_080=3.36e-05 mcrdll1f_cc_w_0_170_s_1_080=2.02e-11 mcrdll1f_cf_w_0_170_s_1_080=1.55e-11
+  mcrdll1f_ca_w_0_170_s_1_980=3.36e-05 mcrdll1f_cc_w_0_170_s_1_980=1.08e-11 mcrdll1f_cf_w_0_170_s_1_980=2.21e-11
+  mcrdll1f_ca_w_0_170_s_4_500=3.36e-05 mcrdll1f_cc_w_0_170_s_4_500=2.88e-12 mcrdll1f_cf_w_0_170_s_4_500=2.91e-11
+  mcrdll1f_ca_w_1_360_s_0_180=3.36e-05 mcrdll1f_cc_w_1_360_s_0_180=9.08e-11 mcrdll1f_cf_w_1_360_s_0_180=3.36e-12
+  mcrdll1f_ca_w_1_360_s_0_225=3.36e-05 mcrdll1f_cc_w_1_360_s_0_225=8.07e-11 mcrdll1f_cf_w_1_360_s_0_225=4.08e-12
+  mcrdll1f_ca_w_1_360_s_0_270=3.36e-05 mcrdll1f_cc_w_1_360_s_0_270=7.32e-11 mcrdll1f_cf_w_1_360_s_0_270=4.79e-12
+  mcrdll1f_ca_w_1_360_s_0_360=3.36e-05 mcrdll1f_cc_w_1_360_s_0_360=6.24e-11 mcrdll1f_cf_w_1_360_s_0_360=6.20e-12
+  mcrdll1f_ca_w_1_360_s_0_450=3.36e-05 mcrdll1f_cc_w_1_360_s_0_450=5.49e-11 mcrdll1f_cf_w_1_360_s_0_450=7.54e-12
+  mcrdll1f_ca_w_1_360_s_0_540=3.36e-05 mcrdll1f_cc_w_1_360_s_0_540=4.92e-11 mcrdll1f_cf_w_1_360_s_0_540=8.84e-12
+  mcrdll1f_ca_w_1_360_s_0_720=3.36e-05 mcrdll1f_cc_w_1_360_s_0_720=4.09e-11 mcrdll1f_cf_w_1_360_s_0_720=1.13e-11
+  mcrdll1f_ca_w_1_360_s_1_080=3.36e-05 mcrdll1f_cc_w_1_360_s_1_080=3.05e-11 mcrdll1f_cf_w_1_360_s_1_080=1.57e-11
+  mcrdll1f_ca_w_1_360_s_1_980=3.36e-05 mcrdll1f_cc_w_1_360_s_1_980=1.74e-11 mcrdll1f_cf_w_1_360_s_1_980=2.39e-11
+  mcrdll1f_ca_w_1_360_s_4_500=3.36e-05 mcrdll1f_cc_w_1_360_s_4_500=5.54e-12 mcrdll1f_cf_w_1_360_s_4_500=3.39e-11
+  mcrdll1d_ca_w_0_170_s_0_180=5.02e-05 mcrdll1d_cc_w_0_170_s_0_180=6.66e-11 mcrdll1d_cf_w_0_170_s_0_180=4.96e-12
+  mcrdll1d_ca_w_0_170_s_0_225=5.02e-05 mcrdll1d_cc_w_0_170_s_0_225=5.77e-11 mcrdll1d_cf_w_0_170_s_0_225=5.99e-12
+  mcrdll1d_ca_w_0_170_s_0_270=5.02e-05 mcrdll1d_cc_w_0_170_s_0_270=5.17e-11 mcrdll1d_cf_w_0_170_s_0_270=7.00e-12
+  mcrdll1d_ca_w_0_170_s_0_360=5.02e-05 mcrdll1d_cc_w_0_170_s_0_360=4.23e-11 mcrdll1d_cf_w_0_170_s_0_360=9.15e-12
+  mcrdll1d_ca_w_0_170_s_0_450=5.02e-05 mcrdll1d_cc_w_0_170_s_0_450=3.65e-11 mcrdll1d_cf_w_0_170_s_0_450=1.08e-11
+  mcrdll1d_ca_w_0_170_s_0_540=5.02e-05 mcrdll1d_cc_w_0_170_s_0_540=3.14e-11 mcrdll1d_cf_w_0_170_s_0_540=1.28e-11
+  mcrdll1d_ca_w_0_170_s_0_720=5.02e-05 mcrdll1d_cc_w_0_170_s_0_720=2.47e-11 mcrdll1d_cf_w_0_170_s_0_720=1.60e-11
+  mcrdll1d_ca_w_0_170_s_1_080=5.02e-05 mcrdll1d_cc_w_0_170_s_1_080=1.66e-11 mcrdll1d_cf_w_0_170_s_1_080=2.11e-11
+  mcrdll1d_ca_w_0_170_s_1_980=5.02e-05 mcrdll1d_cc_w_0_170_s_1_980=7.79e-12 mcrdll1d_cf_w_0_170_s_1_980=2.81e-11
+  mcrdll1d_ca_w_0_170_s_4_500=5.02e-05 mcrdll1d_cc_w_0_170_s_4_500=1.80e-12 mcrdll1d_cf_w_0_170_s_4_500=3.37e-11
+  mcrdll1d_ca_w_1_360_s_0_180=5.02e-05 mcrdll1d_cc_w_1_360_s_0_180=8.62e-11 mcrdll1d_cf_w_1_360_s_0_180=4.96e-12
+  mcrdll1d_ca_w_1_360_s_0_225=5.02e-05 mcrdll1d_cc_w_1_360_s_0_225=7.62e-11 mcrdll1d_cf_w_1_360_s_0_225=6.00e-12
+  mcrdll1d_ca_w_1_360_s_0_270=5.02e-05 mcrdll1d_cc_w_1_360_s_0_270=6.87e-11 mcrdll1d_cf_w_1_360_s_0_270=7.03e-12
+  mcrdll1d_ca_w_1_360_s_0_360=5.02e-05 mcrdll1d_cc_w_1_360_s_0_360=5.78e-11 mcrdll1d_cf_w_1_360_s_0_360=9.03e-12
+  mcrdll1d_ca_w_1_360_s_0_450=5.02e-05 mcrdll1d_cc_w_1_360_s_0_450=5.03e-11 mcrdll1d_cf_w_1_360_s_0_450=1.09e-11
+  mcrdll1d_ca_w_1_360_s_0_540=5.02e-05 mcrdll1d_cc_w_1_360_s_0_540=4.46e-11 mcrdll1d_cf_w_1_360_s_0_540=1.27e-11
+  mcrdll1d_ca_w_1_360_s_0_720=5.02e-05 mcrdll1d_cc_w_1_360_s_0_720=3.63e-11 mcrdll1d_cf_w_1_360_s_0_720=1.60e-11
+  mcrdll1d_ca_w_1_360_s_1_080=5.02e-05 mcrdll1d_cc_w_1_360_s_1_080=2.62e-11 mcrdll1d_cf_w_1_360_s_1_080=2.16e-11
+  mcrdll1d_ca_w_1_360_s_1_980=5.02e-05 mcrdll1d_cc_w_1_360_s_1_980=1.39e-11 mcrdll1d_cf_w_1_360_s_1_980=3.07e-11
+  mcrdll1d_ca_w_1_360_s_4_500=5.02e-05 mcrdll1d_cc_w_1_360_s_4_500=4.00e-12 mcrdll1d_cf_w_1_360_s_4_500=3.96e-11
+  mcrdll1p1_ca_w_0_170_s_0_180=7.33e-05 mcrdll1p1_cc_w_0_170_s_0_180=6.39e-11 mcrdll1p1_cf_w_0_170_s_0_180=7.16e-12
+  mcrdll1p1_ca_w_0_170_s_0_225=7.33e-05 mcrdll1p1_cc_w_0_170_s_0_225=5.48e-11 mcrdll1p1_cf_w_0_170_s_0_225=8.61e-12
+  mcrdll1p1_ca_w_0_170_s_0_270=7.33e-05 mcrdll1p1_cc_w_0_170_s_0_270=4.86e-11 mcrdll1p1_cf_w_0_170_s_0_270=1.00e-11
+  mcrdll1p1_ca_w_0_170_s_0_360=7.33e-05 mcrdll1p1_cc_w_0_170_s_0_360=3.89e-11 mcrdll1p1_cf_w_0_170_s_0_360=1.29e-11
+  mcrdll1p1_ca_w_0_170_s_0_450=7.33e-05 mcrdll1p1_cc_w_0_170_s_0_450=3.30e-11 mcrdll1p1_cf_w_0_170_s_0_450=1.52e-11
+  mcrdll1p1_ca_w_0_170_s_0_540=7.33e-05 mcrdll1p1_cc_w_0_170_s_0_540=2.78e-11 mcrdll1p1_cf_w_0_170_s_0_540=1.77e-11
+  mcrdll1p1_ca_w_0_170_s_0_720=7.33e-05 mcrdll1p1_cc_w_0_170_s_0_720=2.11e-11 mcrdll1p1_cf_w_0_170_s_0_720=2.17e-11
+  mcrdll1p1_ca_w_0_170_s_1_080=7.33e-05 mcrdll1p1_cc_w_0_170_s_1_080=1.32e-11 mcrdll1p1_cf_w_0_170_s_1_080=2.74e-11
+  mcrdll1p1_ca_w_0_170_s_1_980=7.33e-05 mcrdll1p1_cc_w_0_170_s_1_980=5.59e-12 mcrdll1p1_cf_w_0_170_s_1_980=3.41e-11
+  mcrdll1p1_ca_w_0_170_s_4_500=7.33e-05 mcrdll1p1_cc_w_0_170_s_4_500=1.19e-12 mcrdll1p1_cf_w_0_170_s_4_500=3.83e-11
+  mcrdll1p1_ca_w_1_360_s_0_180=7.33e-05 mcrdll1p1_cc_w_1_360_s_0_180=8.18e-11 mcrdll1p1_cf_w_1_360_s_0_180=7.21e-12
+  mcrdll1p1_ca_w_1_360_s_0_225=7.33e-05 mcrdll1p1_cc_w_1_360_s_0_225=7.19e-11 mcrdll1p1_cf_w_1_360_s_0_225=8.68e-12
+  mcrdll1p1_ca_w_1_360_s_0_270=7.33e-05 mcrdll1p1_cc_w_1_360_s_0_270=6.43e-11 mcrdll1p1_cf_w_1_360_s_0_270=1.01e-11
+  mcrdll1p1_ca_w_1_360_s_0_360=7.33e-05 mcrdll1p1_cc_w_1_360_s_0_360=5.35e-11 mcrdll1p1_cf_w_1_360_s_0_360=1.28e-11
+  mcrdll1p1_ca_w_1_360_s_0_450=7.33e-05 mcrdll1p1_cc_w_1_360_s_0_450=4.60e-11 mcrdll1p1_cf_w_1_360_s_0_450=1.54e-11
+  mcrdll1p1_ca_w_1_360_s_0_540=7.33e-05 mcrdll1p1_cc_w_1_360_s_0_540=4.03e-11 mcrdll1p1_cf_w_1_360_s_0_540=1.78e-11
+  mcrdll1p1_ca_w_1_360_s_0_720=7.33e-05 mcrdll1p1_cc_w_1_360_s_0_720=3.22e-11 mcrdll1p1_cf_w_1_360_s_0_720=2.19e-11
+  mcrdll1p1_ca_w_1_360_s_1_080=7.33e-05 mcrdll1p1_cc_w_1_360_s_1_080=2.24e-11 mcrdll1p1_cf_w_1_360_s_1_080=2.84e-11
+  mcrdll1p1_ca_w_1_360_s_1_980=7.33e-05 mcrdll1p1_cc_w_1_360_s_1_980=1.11e-11 mcrdll1p1_cf_w_1_360_s_1_980=3.77e-11
+  mcrdll1p1_ca_w_1_360_s_4_500=7.33e-05 mcrdll1p1_cc_w_1_360_s_4_500=3.00e-12 mcrdll1p1_cf_w_1_360_s_4_500=4.53e-11
+  mcm2m1f_ca_w_0_140_s_0_140=1.12e-04 mcm2m1f_cc_w_0_140_s_0_140=8.26e-11 mcm2m1f_cf_w_0_140_s_0_140=8.34e-12
+  mcm2m1f_ca_w_0_140_s_0_175=1.12e-04 mcm2m1f_cc_w_0_140_s_0_175=8.06e-11 mcm2m1f_cf_w_0_140_s_0_175=1.00e-11
+  mcm2m1f_ca_w_0_140_s_0_210=1.12e-04 mcm2m1f_cc_w_0_140_s_0_210=7.70e-11 mcm2m1f_cf_w_0_140_s_0_210=1.18e-11
+  mcm2m1f_ca_w_0_140_s_0_280=1.12e-04 mcm2m1f_cc_w_0_140_s_0_280=6.72e-11 mcm2m1f_cf_w_0_140_s_0_280=1.50e-11
+  mcm2m1f_ca_w_0_140_s_0_350=1.12e-04 mcm2m1f_cc_w_0_140_s_0_350=5.65e-11 mcm2m1f_cf_w_0_140_s_0_350=1.81e-11
+  mcm2m1f_ca_w_0_140_s_0_420=1.12e-04 mcm2m1f_cc_w_0_140_s_0_420=4.77e-11 mcm2m1f_cf_w_0_140_s_0_420=2.11e-11
+  mcm2m1f_ca_w_0_140_s_0_560=1.12e-04 mcm2m1f_cc_w_0_140_s_0_560=3.53e-11 mcm2m1f_cf_w_0_140_s_0_560=2.61e-11
+  mcm2m1f_ca_w_0_140_s_0_840=1.12e-04 mcm2m1f_cc_w_0_140_s_0_840=2.11e-11 mcm2m1f_cf_w_0_140_s_0_840=3.43e-11
+  mcm2m1f_ca_w_0_140_s_1_540=1.12e-04 mcm2m1f_cc_w_0_140_s_1_540=7.08e-12 mcm2m1f_cf_w_0_140_s_1_540=4.54e-11
+  mcm2m1f_ca_w_0_140_s_3_500=1.12e-04 mcm2m1f_cc_w_0_140_s_3_500=5.50e-13 mcm2m1f_cf_w_0_140_s_3_500=5.18e-11
+  mcm2m1f_ca_w_1_120_s_0_140=1.12e-04 mcm2m1f_cc_w_1_120_s_0_140=9.41e-11 mcm2m1f_cf_w_1_120_s_0_140=8.39e-12
+  mcm2m1f_ca_w_1_120_s_0_175=1.12e-04 mcm2m1f_cc_w_1_120_s_0_175=9.12e-11 mcm2m1f_cf_w_1_120_s_0_175=1.01e-11
+  mcm2m1f_ca_w_1_120_s_0_210=1.12e-04 mcm2m1f_cc_w_1_120_s_0_210=8.62e-11 mcm2m1f_cf_w_1_120_s_0_210=1.18e-11
+  mcm2m1f_ca_w_1_120_s_0_280=1.12e-04 mcm2m1f_cc_w_1_120_s_0_280=7.45e-11 mcm2m1f_cf_w_1_120_s_0_280=1.51e-11
+  mcm2m1f_ca_w_1_120_s_0_350=1.12e-04 mcm2m1f_cc_w_1_120_s_0_350=6.32e-11 mcm2m1f_cf_w_1_120_s_0_350=1.82e-11
+  mcm2m1f_ca_w_1_120_s_0_420=1.12e-04 mcm2m1f_cc_w_1_120_s_0_420=5.36e-11 mcm2m1f_cf_w_1_120_s_0_420=2.12e-11
+  mcm2m1f_ca_w_1_120_s_0_560=1.12e-04 mcm2m1f_cc_w_1_120_s_0_560=3.98e-11 mcm2m1f_cf_w_1_120_s_0_560=2.65e-11
+  mcm2m1f_ca_w_1_120_s_0_840=1.12e-04 mcm2m1f_cc_w_1_120_s_0_840=2.42e-11 mcm2m1f_cf_w_1_120_s_0_840=3.49e-11
+  mcm2m1f_ca_w_1_120_s_1_540=1.12e-04 mcm2m1f_cc_w_1_120_s_1_540=8.50e-12 mcm2m1f_cf_w_1_120_s_1_540=4.68e-11
+  mcm2m1f_ca_w_1_120_s_3_500=1.12e-04 mcm2m1f_cc_w_1_120_s_3_500=6.85e-13 mcm2m1f_cf_w_1_120_s_3_500=5.43e-11
+  mcm2m1d_ca_w_0_140_s_0_140=1.19e-04 mcm2m1d_cc_w_0_140_s_0_140=8.21e-11 mcm2m1d_cf_w_0_140_s_0_140=8.87e-12
+  mcm2m1d_ca_w_0_140_s_0_175=1.19e-04 mcm2m1d_cc_w_0_140_s_0_175=7.97e-11 mcm2m1d_cf_w_0_140_s_0_175=1.07e-11
+  mcm2m1d_ca_w_0_140_s_0_210=1.19e-04 mcm2m1d_cc_w_0_140_s_0_210=7.60e-11 mcm2m1d_cf_w_0_140_s_0_210=1.25e-11
+  mcm2m1d_ca_w_0_140_s_0_280=1.19e-04 mcm2m1d_cc_w_0_140_s_0_280=6.59e-11 mcm2m1d_cf_w_0_140_s_0_280=1.60e-11
+  mcm2m1d_ca_w_0_140_s_0_350=1.19e-04 mcm2m1d_cc_w_0_140_s_0_350=5.52e-11 mcm2m1d_cf_w_0_140_s_0_350=1.93e-11
+  mcm2m1d_ca_w_0_140_s_0_420=1.19e-04 mcm2m1d_cc_w_0_140_s_0_420=4.61e-11 mcm2m1d_cf_w_0_140_s_0_420=2.25e-11
+  mcm2m1d_ca_w_0_140_s_0_560=1.19e-04 mcm2m1d_cc_w_0_140_s_0_560=3.36e-11 mcm2m1d_cf_w_0_140_s_0_560=2.79e-11
+  mcm2m1d_ca_w_0_140_s_0_840=1.19e-04 mcm2m1d_cc_w_0_140_s_0_840=1.93e-11 mcm2m1d_cf_w_0_140_s_0_840=3.65e-11
+  mcm2m1d_ca_w_0_140_s_1_540=1.19e-04 mcm2m1d_cc_w_0_140_s_1_540=5.78e-12 mcm2m1d_cf_w_0_140_s_1_540=4.75e-11
+  mcm2m1d_ca_w_0_140_s_3_500=1.19e-04 mcm2m1d_cc_w_0_140_s_3_500=3.20e-13 mcm2m1d_cf_w_0_140_s_3_500=5.30e-11
+  mcm2m1d_ca_w_1_120_s_0_140=1.19e-04 mcm2m1d_cc_w_1_120_s_0_140=9.20e-11 mcm2m1d_cf_w_1_120_s_0_140=8.95e-12
+  mcm2m1d_ca_w_1_120_s_0_175=1.19e-04 mcm2m1d_cc_w_1_120_s_0_175=8.86e-11 mcm2m1d_cf_w_1_120_s_0_175=1.08e-11
+  mcm2m1d_ca_w_1_120_s_0_210=1.19e-04 mcm2m1d_cc_w_1_120_s_0_210=8.36e-11 mcm2m1d_cf_w_1_120_s_0_210=1.26e-11
+  mcm2m1d_ca_w_1_120_s_0_280=1.19e-04 mcm2m1d_cc_w_1_120_s_0_280=7.18e-11 mcm2m1d_cf_w_1_120_s_0_280=1.61e-11
+  mcm2m1d_ca_w_1_120_s_0_350=1.19e-04 mcm2m1d_cc_w_1_120_s_0_350=6.05e-11 mcm2m1d_cf_w_1_120_s_0_350=1.94e-11
+  mcm2m1d_ca_w_1_120_s_0_420=1.19e-04 mcm2m1d_cc_w_1_120_s_0_420=5.09e-11 mcm2m1d_cf_w_1_120_s_0_420=2.26e-11
+  mcm2m1d_ca_w_1_120_s_0_560=1.19e-04 mcm2m1d_cc_w_1_120_s_0_560=3.71e-11 mcm2m1d_cf_w_1_120_s_0_560=2.82e-11
+  mcm2m1d_ca_w_1_120_s_0_840=1.19e-04 mcm2m1d_cc_w_1_120_s_0_840=2.15e-11 mcm2m1d_cf_w_1_120_s_0_840=3.71e-11
+  mcm2m1d_ca_w_1_120_s_1_540=1.19e-04 mcm2m1d_cc_w_1_120_s_1_540=6.60e-12 mcm2m1d_cf_w_1_120_s_1_540=4.87e-11
+  mcm2m1d_ca_w_1_120_s_3_500=1.19e-04 mcm2m1d_cc_w_1_120_s_3_500=3.60e-13 mcm2m1d_cf_w_1_120_s_3_500=5.51e-11
+  mcm2m1p1_ca_w_0_140_s_0_140=1.26e-04 mcm2m1p1_cc_w_0_140_s_0_140=8.13e-11 mcm2m1p1_cf_w_0_140_s_0_140=9.42e-12
+  mcm2m1p1_ca_w_0_140_s_0_175=1.26e-04 mcm2m1p1_cc_w_0_140_s_0_175=7.88e-11 mcm2m1p1_cf_w_0_140_s_0_175=1.14e-11
+  mcm2m1p1_ca_w_0_140_s_0_210=1.26e-04 mcm2m1p1_cc_w_0_140_s_0_210=7.50e-11 mcm2m1p1_cf_w_0_140_s_0_210=1.33e-11
+  mcm2m1p1_ca_w_0_140_s_0_280=1.26e-04 mcm2m1p1_cc_w_0_140_s_0_280=6.48e-11 mcm2m1p1_cf_w_0_140_s_0_280=1.70e-11
+  mcm2m1p1_ca_w_0_140_s_0_350=1.26e-04 mcm2m1p1_cc_w_0_140_s_0_350=5.39e-11 mcm2m1p1_cf_w_0_140_s_0_350=2.06e-11
+  mcm2m1p1_ca_w_0_140_s_0_420=1.26e-04 mcm2m1p1_cc_w_0_140_s_0_420=4.47e-11 mcm2m1p1_cf_w_0_140_s_0_420=2.40e-11
+  mcm2m1p1_ca_w_0_140_s_0_560=1.26e-04 mcm2m1p1_cc_w_0_140_s_0_560=3.21e-11 mcm2m1p1_cf_w_0_140_s_0_560=2.96e-11
+  mcm2m1p1_ca_w_0_140_s_0_840=1.26e-04 mcm2m1p1_cc_w_0_140_s_0_840=1.78e-11 mcm2m1p1_cf_w_0_140_s_0_840=3.86e-11
+  mcm2m1p1_ca_w_0_140_s_1_540=1.26e-04 mcm2m1p1_cc_w_0_140_s_1_540=4.71e-12 mcm2m1p1_cf_w_0_140_s_1_540=4.97e-11
+  mcm2m1p1_ca_w_0_140_s_3_500=1.26e-04 mcm2m1p1_cc_w_0_140_s_3_500=2.05e-13 mcm2m1p1_cf_w_0_140_s_3_500=5.41e-11
+  mcm2m1p1_ca_w_1_120_s_0_140=1.26e-04 mcm2m1p1_cc_w_1_120_s_0_140=8.96e-11 mcm2m1p1_cf_w_1_120_s_0_140=9.53e-12
+  mcm2m1p1_ca_w_1_120_s_0_175=1.26e-04 mcm2m1p1_cc_w_1_120_s_0_175=8.62e-11 mcm2m1p1_cf_w_1_120_s_0_175=1.15e-11
+  mcm2m1p1_ca_w_1_120_s_0_210=1.26e-04 mcm2m1p1_cc_w_1_120_s_0_210=8.13e-11 mcm2m1p1_cf_w_1_120_s_0_210=1.34e-11
+  mcm2m1p1_ca_w_1_120_s_0_280=1.26e-04 mcm2m1p1_cc_w_1_120_s_0_280=6.94e-11 mcm2m1p1_cf_w_1_120_s_0_280=1.71e-11
+  mcm2m1p1_ca_w_1_120_s_0_350=1.26e-04 mcm2m1p1_cc_w_1_120_s_0_350=5.78e-11 mcm2m1p1_cf_w_1_120_s_0_350=2.07e-11
+  mcm2m1p1_ca_w_1_120_s_0_420=1.26e-04 mcm2m1p1_cc_w_1_120_s_0_420=4.84e-11 mcm2m1p1_cf_w_1_120_s_0_420=2.41e-11
+  mcm2m1p1_ca_w_1_120_s_0_560=1.26e-04 mcm2m1p1_cc_w_1_120_s_0_560=3.47e-11 mcm2m1p1_cf_w_1_120_s_0_560=3.00e-11
+  mcm2m1p1_ca_w_1_120_s_0_840=1.26e-04 mcm2m1p1_cc_w_1_120_s_0_840=1.94e-11 mcm2m1p1_cf_w_1_120_s_0_840=3.92e-11
+  mcm2m1p1_ca_w_1_120_s_1_540=1.26e-04 mcm2m1p1_cc_w_1_120_s_1_540=5.20e-12 mcm2m1p1_cf_w_1_120_s_1_540=5.08e-11
+  mcm2m1p1_ca_w_1_120_s_3_500=1.26e-04 mcm2m1p1_cc_w_1_120_s_3_500=2.35e-13 mcm2m1p1_cf_w_1_120_s_3_500=5.58e-11
+  mcm2m1l1_ca_w_0_140_s_0_140=1.78e-04 mcm2m1l1_cc_w_0_140_s_0_140=7.58e-11 mcm2m1l1_cf_w_0_140_s_0_140=1.32e-11
+  mcm2m1l1_ca_w_0_140_s_0_175=1.78e-04 mcm2m1l1_cc_w_0_140_s_0_175=7.34e-11 mcm2m1l1_cf_w_0_140_s_0_175=1.61e-11
+  mcm2m1l1_ca_w_0_140_s_0_210=1.78e-04 mcm2m1l1_cc_w_0_140_s_0_210=6.93e-11 mcm2m1l1_cf_w_0_140_s_0_210=1.88e-11
+  mcm2m1l1_ca_w_0_140_s_0_280=1.78e-04 mcm2m1l1_cc_w_0_140_s_0_280=5.77e-11 mcm2m1l1_cf_w_0_140_s_0_280=2.41e-11
+  mcm2m1l1_ca_w_0_140_s_0_350=1.78e-04 mcm2m1l1_cc_w_0_140_s_0_350=4.66e-11 mcm2m1l1_cf_w_0_140_s_0_350=2.90e-11
+  mcm2m1l1_ca_w_0_140_s_0_420=1.78e-04 mcm2m1l1_cc_w_0_140_s_0_420=3.73e-11 mcm2m1l1_cf_w_0_140_s_0_420=3.36e-11
+  mcm2m1l1_ca_w_0_140_s_0_560=1.78e-04 mcm2m1l1_cc_w_0_140_s_0_560=2.45e-11 mcm2m1l1_cf_w_0_140_s_0_560=4.11e-11
+  mcm2m1l1_ca_w_0_140_s_0_840=1.78e-04 mcm2m1l1_cc_w_0_140_s_0_840=1.10e-11 mcm2m1l1_cf_w_0_140_s_0_840=5.14e-11
+  mcm2m1l1_ca_w_0_140_s_1_540=1.78e-04 mcm2m1l1_cc_w_0_140_s_1_540=1.64e-12 mcm2m1l1_cf_w_0_140_s_1_540=6.06e-11
+  mcm2m1l1_ca_w_0_140_s_3_500=1.78e-04 mcm2m1l1_cc_w_0_140_s_3_500=7.00e-14 mcm2m1l1_cf_w_0_140_s_3_500=6.27e-11
+  mcm2m1l1_ca_w_1_120_s_0_140=1.78e-04 mcm2m1l1_cc_w_1_120_s_0_140=7.92e-11 mcm2m1l1_cf_w_1_120_s_0_140=1.33e-11
+  mcm2m1l1_ca_w_1_120_s_0_175=1.78e-04 mcm2m1l1_cc_w_1_120_s_0_175=7.61e-11 mcm2m1l1_cf_w_1_120_s_0_175=1.62e-11
+  mcm2m1l1_ca_w_1_120_s_0_210=1.78e-04 mcm2m1l1_cc_w_1_120_s_0_210=7.14e-11 mcm2m1l1_cf_w_1_120_s_0_210=1.89e-11
+  mcm2m1l1_ca_w_1_120_s_0_280=1.78e-04 mcm2m1l1_cc_w_1_120_s_0_280=5.93e-11 mcm2m1l1_cf_w_1_120_s_0_280=2.42e-11
+  mcm2m1l1_ca_w_1_120_s_0_350=1.78e-04 mcm2m1l1_cc_w_1_120_s_0_350=4.79e-11 mcm2m1l1_cf_w_1_120_s_0_350=2.92e-11
+  mcm2m1l1_ca_w_1_120_s_0_420=1.78e-04 mcm2m1l1_cc_w_1_120_s_0_420=3.82e-11 mcm2m1l1_cf_w_1_120_s_0_420=3.37e-11
+  mcm2m1l1_ca_w_1_120_s_0_560=1.78e-04 mcm2m1l1_cc_w_1_120_s_0_560=2.51e-11 mcm2m1l1_cf_w_1_120_s_0_560=4.14e-11
+  mcm2m1l1_ca_w_1_120_s_0_840=1.78e-04 mcm2m1l1_cc_w_1_120_s_0_840=1.14e-11 mcm2m1l1_cf_w_1_120_s_0_840=5.19e-11
+  mcm2m1l1_ca_w_1_120_s_1_540=1.78e-04 mcm2m1l1_cc_w_1_120_s_1_540=1.65e-12 mcm2m1l1_cf_w_1_120_s_1_540=6.13e-11
+  mcm2m1l1_ca_w_1_120_s_3_500=1.78e-04 mcm2m1l1_cc_w_1_120_s_3_500=5.00e-14 mcm2m1l1_cf_w_1_120_s_3_500=6.34e-11
+  mcm3m1f_ca_w_0_140_s_0_140=4.93e-05 mcm3m1f_cc_w_0_140_s_0_140=8.88e-11 mcm3m1f_cf_w_0_140_s_0_140=3.90e-12
+  mcm3m1f_ca_w_0_140_s_0_175=4.93e-05 mcm3m1f_cc_w_0_140_s_0_175=8.68e-11 mcm3m1f_cf_w_0_140_s_0_175=4.73e-12
+  mcm3m1f_ca_w_0_140_s_0_210=4.93e-05 mcm3m1f_cc_w_0_140_s_0_210=8.36e-11 mcm3m1f_cf_w_0_140_s_0_210=5.59e-12
+  mcm3m1f_ca_w_0_140_s_0_280=4.93e-05 mcm3m1f_cc_w_0_140_s_0_280=7.48e-11 mcm3m1f_cf_w_0_140_s_0_280=7.20e-12
+  mcm3m1f_ca_w_0_140_s_0_350=4.93e-05 mcm3m1f_cc_w_0_140_s_0_350=6.47e-11 mcm3m1f_cf_w_0_140_s_0_350=8.80e-12
+  mcm3m1f_ca_w_0_140_s_0_420=4.93e-05 mcm3m1f_cc_w_0_140_s_0_420=5.64e-11 mcm3m1f_cf_w_0_140_s_0_420=1.04e-11
+  mcm3m1f_ca_w_0_140_s_0_560=4.93e-05 mcm3m1f_cc_w_0_140_s_0_560=4.44e-11 mcm3m1f_cf_w_0_140_s_0_560=1.34e-11
+  mcm3m1f_ca_w_0_140_s_0_840=4.93e-05 mcm3m1f_cc_w_0_140_s_0_840=3.03e-11 mcm3m1f_cf_w_0_140_s_0_840=1.87e-11
+  mcm3m1f_ca_w_0_140_s_1_540=4.93e-05 mcm3m1f_cc_w_0_140_s_1_540=1.37e-11 mcm3m1f_cf_w_0_140_s_1_540=2.83e-11
+  mcm3m1f_ca_w_0_140_s_3_500=4.93e-05 mcm3m1f_cc_w_0_140_s_3_500=1.99e-12 mcm3m1f_cf_w_0_140_s_3_500=3.82e-11
+  mcm3m1f_ca_w_1_120_s_0_140=4.93e-05 mcm3m1f_cc_w_1_120_s_0_140=1.08e-10 mcm3m1f_cf_w_1_120_s_0_140=3.93e-12
+  mcm3m1f_ca_w_1_120_s_0_175=4.93e-05 mcm3m1f_cc_w_1_120_s_0_175=1.03e-10 mcm3m1f_cf_w_1_120_s_0_175=4.77e-12
+  mcm3m1f_ca_w_1_120_s_0_210=4.93e-05 mcm3m1f_cc_w_1_120_s_0_210=9.87e-11 mcm3m1f_cf_w_1_120_s_0_210=5.58e-12
+  mcm3m1f_ca_w_1_120_s_0_280=4.93e-05 mcm3m1f_cc_w_1_120_s_0_280=8.69e-11 mcm3m1f_cf_w_1_120_s_0_280=7.26e-12
+  mcm3m1f_ca_w_1_120_s_0_350=4.93e-05 mcm3m1f_cc_w_1_120_s_0_350=7.56e-11 mcm3m1f_cf_w_1_120_s_0_350=8.85e-12
+  mcm3m1f_ca_w_1_120_s_0_420=4.93e-05 mcm3m1f_cc_w_1_120_s_0_420=6.60e-11 mcm3m1f_cf_w_1_120_s_0_420=1.05e-11
+  mcm3m1f_ca_w_1_120_s_0_560=4.93e-05 mcm3m1f_cc_w_1_120_s_0_560=5.20e-11 mcm3m1f_cf_w_1_120_s_0_560=1.35e-11
+  mcm3m1f_ca_w_1_120_s_0_840=4.93e-05 mcm3m1f_cc_w_1_120_s_0_840=3.53e-11 mcm3m1f_cf_w_1_120_s_0_840=1.90e-11
+  mcm3m1f_ca_w_1_120_s_1_540=4.93e-05 mcm3m1f_cc_w_1_120_s_1_540=1.62e-11 mcm3m1f_cf_w_1_120_s_1_540=2.94e-11
+  mcm3m1f_ca_w_1_120_s_3_500=4.93e-05 mcm3m1f_cc_w_1_120_s_3_500=2.41e-12 mcm3m1f_cf_w_1_120_s_3_500=4.08e-11
+  mcm3m1d_ca_w_0_140_s_0_140=5.62e-05 mcm3m1d_cc_w_0_140_s_0_140=8.80e-11 mcm3m1d_cf_w_0_140_s_0_140=4.44e-12
+  mcm3m1d_ca_w_0_140_s_0_175=5.62e-05 mcm3m1d_cc_w_0_140_s_0_175=8.59e-11 mcm3m1d_cf_w_0_140_s_0_175=5.39e-12
+  mcm3m1d_ca_w_0_140_s_0_210=5.62e-05 mcm3m1d_cc_w_0_140_s_0_210=8.31e-11 mcm3m1d_cf_w_0_140_s_0_210=6.38e-12
+  mcm3m1d_ca_w_0_140_s_0_280=5.62e-05 mcm3m1d_cc_w_0_140_s_0_280=7.37e-11 mcm3m1d_cf_w_0_140_s_0_280=8.21e-12
+  mcm3m1d_ca_w_0_140_s_0_350=5.62e-05 mcm3m1d_cc_w_0_140_s_0_350=6.33e-11 mcm3m1d_cf_w_0_140_s_0_350=1.00e-11
+  mcm3m1d_ca_w_0_140_s_0_420=5.62e-05 mcm3m1d_cc_w_0_140_s_0_420=5.51e-11 mcm3m1d_cf_w_0_140_s_0_420=1.19e-11
+  mcm3m1d_ca_w_0_140_s_0_560=5.62e-05 mcm3m1d_cc_w_0_140_s_0_560=4.28e-11 mcm3m1d_cf_w_0_140_s_0_560=1.52e-11
+  mcm3m1d_ca_w_0_140_s_0_840=5.62e-05 mcm3m1d_cc_w_0_140_s_0_840=2.84e-11 mcm3m1d_cf_w_0_140_s_0_840=2.11e-11
+  mcm3m1d_ca_w_0_140_s_1_540=5.62e-05 mcm3m1d_cc_w_0_140_s_1_540=1.19e-11 mcm3m1d_cf_w_0_140_s_1_540=3.14e-11
+  mcm3m1d_ca_w_0_140_s_3_500=5.62e-05 mcm3m1d_cc_w_0_140_s_3_500=1.36e-12 mcm3m1d_cf_w_0_140_s_3_500=4.06e-11
+  mcm3m1d_ca_w_1_120_s_0_140=5.62e-05 mcm3m1d_cc_w_1_120_s_0_140=1.05e-10 mcm3m1d_cf_w_1_120_s_0_140=4.48e-12
+  mcm3m1d_ca_w_1_120_s_0_175=5.62e-05 mcm3m1d_cc_w_1_120_s_0_175=1.01e-10 mcm3m1d_cf_w_1_120_s_0_175=5.45e-12
+  mcm3m1d_ca_w_1_120_s_0_210=5.62e-05 mcm3m1d_cc_w_1_120_s_0_210=9.59e-11 mcm3m1d_cf_w_1_120_s_0_210=6.39e-12
+  mcm3m1d_ca_w_1_120_s_0_280=5.62e-05 mcm3m1d_cc_w_1_120_s_0_280=8.42e-11 mcm3m1d_cf_w_1_120_s_0_280=8.27e-12
+  mcm3m1d_ca_w_1_120_s_0_350=5.62e-05 mcm3m1d_cc_w_1_120_s_0_350=7.28e-11 mcm3m1d_cf_w_1_120_s_0_350=1.01e-11
+  mcm3m1d_ca_w_1_120_s_0_420=5.62e-05 mcm3m1d_cc_w_1_120_s_0_420=6.31e-11 mcm3m1d_cf_w_1_120_s_0_420=1.19e-11
+  mcm3m1d_ca_w_1_120_s_0_560=5.62e-05 mcm3m1d_cc_w_1_120_s_0_560=4.91e-11 mcm3m1d_cf_w_1_120_s_0_560=1.53e-11
+  mcm3m1d_ca_w_1_120_s_0_840=5.62e-05 mcm3m1d_cc_w_1_120_s_0_840=3.24e-11 mcm3m1d_cf_w_1_120_s_0_840=2.14e-11
+  mcm3m1d_ca_w_1_120_s_1_540=5.62e-05 mcm3m1d_cc_w_1_120_s_1_540=1.39e-11 mcm3m1d_cf_w_1_120_s_1_540=3.24e-11
+  mcm3m1d_ca_w_1_120_s_3_500=5.62e-05 mcm3m1d_cc_w_1_120_s_3_500=1.58e-12 mcm3m1d_cf_w_1_120_s_3_500=4.30e-11
+  mcm3m1p1_ca_w_0_140_s_0_140=6.31e-05 mcm3m1p1_cc_w_0_140_s_0_140=8.73e-11 mcm3m1p1_cf_w_0_140_s_0_140=4.99e-12
+  mcm3m1p1_ca_w_0_140_s_0_175=6.31e-05 mcm3m1p1_cc_w_0_140_s_0_175=8.64e-11 mcm3m1p1_cf_w_0_140_s_0_175=6.06e-12
+  mcm3m1p1_ca_w_0_140_s_0_210=6.31e-05 mcm3m1p1_cc_w_0_140_s_0_210=8.20e-11 mcm3m1p1_cf_w_0_140_s_0_210=7.18e-12
+  mcm3m1p1_ca_w_0_140_s_0_280=6.31e-05 mcm3m1p1_cc_w_0_140_s_0_280=7.25e-11 mcm3m1p1_cf_w_0_140_s_0_280=9.24e-12
+  mcm3m1p1_ca_w_0_140_s_0_350=6.31e-05 mcm3m1p1_cc_w_0_140_s_0_350=6.22e-11 mcm3m1p1_cf_w_0_140_s_0_350=1.13e-11
+  mcm3m1p1_ca_w_0_140_s_0_420=6.31e-05 mcm3m1p1_cc_w_0_140_s_0_420=5.35e-11 mcm3m1p1_cf_w_0_140_s_0_420=1.32e-11
+  mcm3m1p1_ca_w_0_140_s_0_560=6.31e-05 mcm3m1p1_cc_w_0_140_s_0_560=4.13e-11 mcm3m1p1_cf_w_0_140_s_0_560=1.70e-11
+  mcm3m1p1_ca_w_0_140_s_0_840=6.31e-05 mcm3m1p1_cc_w_0_140_s_0_840=2.66e-11 mcm3m1p1_cf_w_0_140_s_0_840=2.34e-11
+  mcm3m1p1_ca_w_0_140_s_1_540=6.31e-05 mcm3m1p1_cc_w_0_140_s_1_540=1.04e-11 mcm3m1p1_cf_w_0_140_s_1_540=3.41e-11
+  mcm3m1p1_ca_w_0_140_s_3_500=6.31e-05 mcm3m1p1_cc_w_0_140_s_3_500=9.80e-13 mcm3m1p1_cf_w_0_140_s_3_500=4.27e-11
+  mcm3m1p1_ca_w_1_120_s_0_140=6.31e-05 mcm3m1p1_cc_w_1_120_s_0_140=1.02e-10 mcm3m1p1_cf_w_1_120_s_0_140=5.09e-12
+  mcm3m1p1_ca_w_1_120_s_0_175=6.31e-05 mcm3m1p1_cc_w_1_120_s_0_175=9.85e-11 mcm3m1p1_cf_w_1_120_s_0_175=6.18e-12
+  mcm3m1p1_ca_w_1_120_s_0_210=6.31e-05 mcm3m1p1_cc_w_1_120_s_0_210=9.37e-11 mcm3m1p1_cf_w_1_120_s_0_210=7.22e-12
+  mcm3m1p1_ca_w_1_120_s_0_280=6.31e-05 mcm3m1p1_cc_w_1_120_s_0_280=8.19e-11 mcm3m1p1_cf_w_1_120_s_0_280=9.34e-12
+  mcm3m1p1_ca_w_1_120_s_0_350=6.31e-05 mcm3m1p1_cc_w_1_120_s_0_350=7.03e-11 mcm3m1p1_cf_w_1_120_s_0_350=1.14e-11
+  mcm3m1p1_ca_w_1_120_s_0_420=6.31e-05 mcm3m1p1_cc_w_1_120_s_0_420=6.08e-11 mcm3m1p1_cf_w_1_120_s_0_420=1.34e-11
+  mcm3m1p1_ca_w_1_120_s_0_560=6.31e-05 mcm3m1p1_cc_w_1_120_s_0_560=4.66e-11 mcm3m1p1_cf_w_1_120_s_0_560=1.71e-11
+  mcm3m1p1_ca_w_1_120_s_0_840=6.31e-05 mcm3m1p1_cc_w_1_120_s_0_840=3.01e-11 mcm3m1p1_cf_w_1_120_s_0_840=2.38e-11
+  mcm3m1p1_ca_w_1_120_s_1_540=6.31e-05 mcm3m1p1_cc_w_1_120_s_1_540=1.20e-11 mcm3m1p1_cf_w_1_120_s_1_540=3.53e-11
+  mcm3m1p1_ca_w_1_120_s_3_500=6.31e-05 mcm3m1p1_cc_w_1_120_s_3_500=1.15e-12 mcm3m1p1_cf_w_1_120_s_3_500=4.49e-11
+  mcm3m1l1_ca_w_0_140_s_0_140=1.15e-04 mcm3m1l1_cc_w_0_140_s_0_140=8.14e-11 mcm3m1l1_cf_w_0_140_s_0_140=8.80e-12
+  mcm3m1l1_ca_w_0_140_s_0_175=1.15e-04 mcm3m1l1_cc_w_0_140_s_0_175=7.97e-11 mcm3m1l1_cf_w_0_140_s_0_175=1.08e-11
+  mcm3m1l1_ca_w_0_140_s_0_210=1.15e-04 mcm3m1l1_cc_w_0_140_s_0_210=7.60e-11 mcm3m1l1_cf_w_0_140_s_0_210=1.27e-11
+  mcm3m1l1_ca_w_0_140_s_0_280=1.15e-04 mcm3m1l1_cc_w_0_140_s_0_280=6.55e-11 mcm3m1l1_cf_w_0_140_s_0_280=1.64e-11
+  mcm3m1l1_ca_w_0_140_s_0_350=1.15e-04 mcm3m1l1_cc_w_0_140_s_0_350=5.47e-11 mcm3m1l1_cf_w_0_140_s_0_350=1.98e-11
+  mcm3m1l1_ca_w_0_140_s_0_420=1.15e-04 mcm3m1l1_cc_w_0_140_s_0_420=4.57e-11 mcm3m1l1_cf_w_0_140_s_0_420=2.30e-11
+  mcm3m1l1_ca_w_0_140_s_0_560=1.15e-04 mcm3m1l1_cc_w_0_140_s_0_560=3.33e-11 mcm3m1l1_cf_w_0_140_s_0_560=2.89e-11
+  mcm3m1l1_ca_w_0_140_s_0_840=1.15e-04 mcm3m1l1_cc_w_0_140_s_0_840=1.90e-11 mcm3m1l1_cf_w_0_140_s_0_840=3.77e-11
+  mcm3m1l1_ca_w_0_140_s_1_540=1.15e-04 mcm3m1l1_cc_w_0_140_s_1_540=5.50e-12 mcm3m1l1_cf_w_0_140_s_1_540=4.88e-11
+  mcm3m1l1_ca_w_0_140_s_3_500=1.15e-04 mcm3m1l1_cc_w_0_140_s_3_500=2.60e-13 mcm3m1l1_cf_w_0_140_s_3_500=5.42e-11
+  mcm3m1l1_ca_w_1_120_s_0_140=1.15e-04 mcm3m1l1_cc_w_1_120_s_0_140=9.25e-11 mcm3m1l1_cf_w_1_120_s_0_140=8.90e-12
+  mcm3m1l1_ca_w_1_120_s_0_175=1.15e-04 mcm3m1l1_cc_w_1_120_s_0_175=8.80e-11 mcm3m1l1_cf_w_1_120_s_0_175=1.09e-11
+  mcm3m1l1_ca_w_1_120_s_0_210=1.15e-04 mcm3m1l1_cc_w_1_120_s_0_210=8.36e-11 mcm3m1l1_cf_w_1_120_s_0_210=1.27e-11
+  mcm3m1l1_ca_w_1_120_s_0_280=1.15e-04 mcm3m1l1_cc_w_1_120_s_0_280=7.15e-11 mcm3m1l1_cf_w_1_120_s_0_280=1.65e-11
+  mcm3m1l1_ca_w_1_120_s_0_350=1.15e-04 mcm3m1l1_cc_w_1_120_s_0_350=6.02e-11 mcm3m1l1_cf_w_1_120_s_0_350=1.99e-11
+  mcm3m1l1_ca_w_1_120_s_0_420=1.15e-04 mcm3m1l1_cc_w_1_120_s_0_420=5.04e-11 mcm3m1l1_cf_w_1_120_s_0_420=2.32e-11
+  mcm3m1l1_ca_w_1_120_s_0_560=1.15e-04 mcm3m1l1_cc_w_1_120_s_0_560=3.68e-11 mcm3m1l1_cf_w_1_120_s_0_560=2.90e-11
+  mcm3m1l1_ca_w_1_120_s_0_840=1.15e-04 mcm3m1l1_cc_w_1_120_s_0_840=2.13e-11 mcm3m1l1_cf_w_1_120_s_0_840=3.82e-11
+  mcm3m1l1_ca_w_1_120_s_1_540=1.15e-04 mcm3m1l1_cc_w_1_120_s_1_540=6.41e-12 mcm3m1l1_cf_w_1_120_s_1_540=5.02e-11
+  mcm3m1l1_ca_w_1_120_s_3_500=1.15e-04 mcm3m1l1_cc_w_1_120_s_3_500=3.05e-13 mcm3m1l1_cf_w_1_120_s_3_500=5.62e-11
+  mcm4m1f_ca_w_0_140_s_0_140=3.51e-05 mcm4m1f_cc_w_0_140_s_0_140=9.07e-11 mcm4m1f_cf_w_0_140_s_0_140=2.81e-12
+  mcm4m1f_ca_w_0_140_s_0_175=3.51e-05 mcm4m1f_cc_w_0_140_s_0_175=9.01e-11 mcm4m1f_cf_w_0_140_s_0_175=3.41e-12
+  mcm4m1f_ca_w_0_140_s_0_210=3.51e-05 mcm4m1f_cc_w_0_140_s_0_210=8.55e-11 mcm4m1f_cf_w_0_140_s_0_210=4.04e-12
+  mcm4m1f_ca_w_0_140_s_0_280=3.51e-05 mcm4m1f_cc_w_0_140_s_0_280=7.74e-11 mcm4m1f_cf_w_0_140_s_0_280=5.21e-12
+  mcm4m1f_ca_w_0_140_s_0_350=3.51e-05 mcm4m1f_cc_w_0_140_s_0_350=6.73e-11 mcm4m1f_cf_w_0_140_s_0_350=6.37e-12
+  mcm4m1f_ca_w_0_140_s_0_420=3.51e-05 mcm4m1f_cc_w_0_140_s_0_420=5.90e-11 mcm4m1f_cf_w_0_140_s_0_420=7.57e-12
+  mcm4m1f_ca_w_0_140_s_0_560=3.51e-05 mcm4m1f_cc_w_0_140_s_0_560=4.79e-11 mcm4m1f_cf_w_0_140_s_0_560=9.79e-12
+  mcm4m1f_ca_w_0_140_s_0_840=3.51e-05 mcm4m1f_cc_w_0_140_s_0_840=3.45e-11 mcm4m1f_cf_w_0_140_s_0_840=1.39e-11
+  mcm4m1f_ca_w_0_140_s_1_540=3.51e-05 mcm4m1f_cc_w_0_140_s_1_540=1.81e-11 mcm4m1f_cf_w_0_140_s_1_540=2.20e-11
+  mcm4m1f_ca_w_0_140_s_3_500=3.51e-05 mcm4m1f_cc_w_0_140_s_3_500=4.16e-12 mcm4m1f_cf_w_0_140_s_3_500=3.26e-11
+  mcm4m1f_ca_w_1_120_s_0_140=3.51e-05 mcm4m1f_cc_w_1_120_s_0_140=1.13e-10 mcm4m1f_cf_w_1_120_s_0_140=2.84e-12
+  mcm4m1f_ca_w_1_120_s_0_175=3.51e-05 mcm4m1f_cc_w_1_120_s_0_175=1.09e-10 mcm4m1f_cf_w_1_120_s_0_175=3.45e-12
+  mcm4m1f_ca_w_1_120_s_0_210=3.51e-05 mcm4m1f_cc_w_1_120_s_0_210=1.05e-10 mcm4m1f_cf_w_1_120_s_0_210=4.04e-12
+  mcm4m1f_ca_w_1_120_s_0_280=3.51e-05 mcm4m1f_cc_w_1_120_s_0_280=9.29e-11 mcm4m1f_cf_w_1_120_s_0_280=5.25e-12
+  mcm4m1f_ca_w_1_120_s_0_350=3.51e-05 mcm4m1f_cc_w_1_120_s_0_350=8.16e-11 mcm4m1f_cf_w_1_120_s_0_350=6.43e-12
+  mcm4m1f_ca_w_1_120_s_0_420=3.51e-05 mcm4m1f_cc_w_1_120_s_0_420=7.21e-11 mcm4m1f_cf_w_1_120_s_0_420=7.61e-12
+  mcm4m1f_ca_w_1_120_s_0_560=3.51e-05 mcm4m1f_cc_w_1_120_s_0_560=5.83e-11 mcm4m1f_cf_w_1_120_s_0_560=9.82e-12
+  mcm4m1f_ca_w_1_120_s_0_840=3.51e-05 mcm4m1f_cc_w_1_120_s_0_840=4.17e-11 mcm4m1f_cf_w_1_120_s_0_840=1.40e-11
+  mcm4m1f_ca_w_1_120_s_1_540=3.51e-05 mcm4m1f_cc_w_1_120_s_1_540=2.23e-11 mcm4m1f_cf_w_1_120_s_1_540=2.27e-11
+  mcm4m1f_ca_w_1_120_s_3_500=3.51e-05 mcm4m1f_cc_w_1_120_s_3_500=5.32e-12 mcm4m1f_cf_w_1_120_s_3_500=3.52e-11
+  mcm4m1d_ca_w_0_140_s_0_140=4.20e-05 mcm4m1d_cc_w_0_140_s_0_140=8.99e-11 mcm4m1d_cf_w_0_140_s_0_140=3.35e-12
+  mcm4m1d_ca_w_0_140_s_0_175=4.20e-05 mcm4m1d_cc_w_0_140_s_0_175=8.92e-11 mcm4m1d_cf_w_0_140_s_0_175=4.07e-12
+  mcm4m1d_ca_w_0_140_s_0_210=4.20e-05 mcm4m1d_cc_w_0_140_s_0_210=8.46e-11 mcm4m1d_cf_w_0_140_s_0_210=4.81e-12
+  mcm4m1d_ca_w_0_140_s_0_280=4.20e-05 mcm4m1d_cc_w_0_140_s_0_280=7.62e-11 mcm4m1d_cf_w_0_140_s_0_280=6.22e-12
+  mcm4m1d_ca_w_0_140_s_0_350=4.20e-05 mcm4m1d_cc_w_0_140_s_0_350=6.61e-11 mcm4m1d_cf_w_0_140_s_0_350=7.60e-12
+  mcm4m1d_ca_w_0_140_s_0_420=4.20e-05 mcm4m1d_cc_w_0_140_s_0_420=5.77e-11 mcm4m1d_cf_w_0_140_s_0_420=9.00e-12
+  mcm4m1d_ca_w_0_140_s_0_560=4.20e-05 mcm4m1d_cc_w_0_140_s_0_560=4.64e-11 mcm4m1d_cf_w_0_140_s_0_560=1.16e-11
+  mcm4m1d_ca_w_0_140_s_0_840=4.20e-05 mcm4m1d_cc_w_0_140_s_0_840=3.24e-11 mcm4m1d_cf_w_0_140_s_0_840=1.63e-11
+  mcm4m1d_ca_w_0_140_s_1_540=4.20e-05 mcm4m1d_cc_w_0_140_s_1_540=1.60e-11 mcm4m1d_cf_w_0_140_s_1_540=2.53e-11
+  mcm4m1d_ca_w_0_140_s_3_500=4.20e-05 mcm4m1d_cc_w_0_140_s_3_500=3.15e-12 mcm4m1d_cf_w_0_140_s_3_500=3.58e-11
+  mcm4m1d_ca_w_1_120_s_0_140=4.20e-05 mcm4m1d_cc_w_1_120_s_0_140=1.10e-10 mcm4m1d_cf_w_1_120_s_0_140=3.39e-12
+  mcm4m1d_ca_w_1_120_s_0_175=4.20e-05 mcm4m1d_cc_w_1_120_s_0_175=1.06e-10 mcm4m1d_cf_w_1_120_s_0_175=4.12e-12
+  mcm4m1d_ca_w_1_120_s_0_210=4.20e-05 mcm4m1d_cc_w_1_120_s_0_210=1.02e-10 mcm4m1d_cf_w_1_120_s_0_210=4.84e-12
+  mcm4m1d_ca_w_1_120_s_0_280=4.20e-05 mcm4m1d_cc_w_1_120_s_0_280=9.03e-11 mcm4m1d_cf_w_1_120_s_0_280=6.27e-12
+  mcm4m1d_ca_w_1_120_s_0_350=4.20e-05 mcm4m1d_cc_w_1_120_s_0_350=7.88e-11 mcm4m1d_cf_w_1_120_s_0_350=7.67e-12
+  mcm4m1d_ca_w_1_120_s_0_420=4.20e-05 mcm4m1d_cc_w_1_120_s_0_420=6.96e-11 mcm4m1d_cf_w_1_120_s_0_420=9.04e-12
+  mcm4m1d_ca_w_1_120_s_0_560=4.20e-05 mcm4m1d_cc_w_1_120_s_0_560=5.53e-11 mcm4m1d_cf_w_1_120_s_0_560=1.17e-11
+  mcm4m1d_ca_w_1_120_s_0_840=4.20e-05 mcm4m1d_cc_w_1_120_s_0_840=3.88e-11 mcm4m1d_cf_w_1_120_s_0_840=1.65e-11
+  mcm4m1d_ca_w_1_120_s_1_540=4.20e-05 mcm4m1d_cc_w_1_120_s_1_540=1.97e-11 mcm4m1d_cf_w_1_120_s_1_540=2.61e-11
+  mcm4m1d_ca_w_1_120_s_3_500=4.20e-05 mcm4m1d_cc_w_1_120_s_3_500=4.05e-12 mcm4m1d_cf_w_1_120_s_3_500=3.84e-11
+  mcm4m1p1_ca_w_0_140_s_0_140=4.90e-05 mcm4m1p1_cc_w_0_140_s_0_140=8.92e-11 mcm4m1p1_cf_w_0_140_s_0_140=3.90e-12
+  mcm4m1p1_ca_w_0_140_s_0_175=4.90e-05 mcm4m1p1_cc_w_0_140_s_0_175=8.84e-11 mcm4m1p1_cf_w_0_140_s_0_175=4.74e-12
+  mcm4m1p1_ca_w_0_140_s_0_210=4.90e-05 mcm4m1p1_cc_w_0_140_s_0_210=8.35e-11 mcm4m1p1_cf_w_0_140_s_0_210=5.61e-12
+  mcm4m1p1_ca_w_0_140_s_0_280=4.90e-05 mcm4m1p1_cc_w_0_140_s_0_280=7.48e-11 mcm4m1p1_cf_w_0_140_s_0_280=7.23e-12
+  mcm4m1p1_ca_w_0_140_s_0_350=4.90e-05 mcm4m1p1_cc_w_0_140_s_0_350=6.50e-11 mcm4m1p1_cf_w_0_140_s_0_350=8.85e-12
+  mcm4m1p1_ca_w_0_140_s_0_420=4.90e-05 mcm4m1p1_cc_w_0_140_s_0_420=5.63e-11 mcm4m1p1_cf_w_0_140_s_0_420=1.04e-11
+  mcm4m1p1_ca_w_0_140_s_0_560=4.90e-05 mcm4m1p1_cc_w_0_140_s_0_560=4.47e-11 mcm4m1p1_cf_w_0_140_s_0_560=1.34e-11
+  mcm4m1p1_ca_w_0_140_s_0_840=4.90e-05 mcm4m1p1_cc_w_0_140_s_0_840=3.06e-11 mcm4m1p1_cf_w_0_140_s_0_840=1.87e-11
+  mcm4m1p1_ca_w_0_140_s_1_540=4.90e-05 mcm4m1p1_cc_w_0_140_s_1_540=1.44e-11 mcm4m1p1_cf_w_0_140_s_1_540=2.84e-11
+  mcm4m1p1_ca_w_0_140_s_3_500=4.90e-05 mcm4m1p1_cc_w_0_140_s_3_500=2.48e-12 mcm4m1p1_cf_w_0_140_s_3_500=3.84e-11
+  mcm4m1p1_ca_w_1_120_s_0_140=4.90e-05 mcm4m1p1_cc_w_1_120_s_0_140=1.07e-10 mcm4m1p1_cf_w_1_120_s_0_140=4.01e-12
+  mcm4m1p1_ca_w_1_120_s_0_175=4.90e-05 mcm4m1p1_cc_w_1_120_s_0_175=1.04e-10 mcm4m1p1_cf_w_1_120_s_0_175=4.85e-12
+  mcm4m1p1_ca_w_1_120_s_0_210=4.90e-05 mcm4m1p1_cc_w_1_120_s_0_210=9.97e-11 mcm4m1p1_cf_w_1_120_s_0_210=5.68e-12
+  mcm4m1p1_ca_w_1_120_s_0_280=4.90e-05 mcm4m1p1_cc_w_1_120_s_0_280=8.78e-11 mcm4m1p1_cf_w_1_120_s_0_280=7.35e-12
+  mcm4m1p1_ca_w_1_120_s_0_350=4.90e-05 mcm4m1p1_cc_w_1_120_s_0_350=7.64e-11 mcm4m1p1_cf_w_1_120_s_0_350=8.96e-12
+  mcm4m1p1_ca_w_1_120_s_0_420=4.90e-05 mcm4m1p1_cc_w_1_120_s_0_420=6.69e-11 mcm4m1p1_cf_w_1_120_s_0_420=1.05e-11
+  mcm4m1p1_ca_w_1_120_s_0_560=4.90e-05 mcm4m1p1_cc_w_1_120_s_0_560=5.30e-11 mcm4m1p1_cf_w_1_120_s_0_560=1.36e-11
+  mcm4m1p1_ca_w_1_120_s_0_840=4.90e-05 mcm4m1p1_cc_w_1_120_s_0_840=3.65e-11 mcm4m1p1_cf_w_1_120_s_0_840=1.90e-11
+  mcm4m1p1_ca_w_1_120_s_1_540=4.90e-05 mcm4m1p1_cc_w_1_120_s_1_540=1.77e-11 mcm4m1p1_cf_w_1_120_s_1_540=2.93e-11
+  mcm4m1p1_ca_w_1_120_s_3_500=4.90e-05 mcm4m1p1_cc_w_1_120_s_3_500=3.25e-12 mcm4m1p1_cf_w_1_120_s_3_500=4.11e-11
+  mcm4m1l1_ca_w_0_140_s_0_140=1.01e-04 mcm4m1l1_cc_w_0_140_s_0_140=8.36e-11 mcm4m1l1_cf_w_0_140_s_0_140=7.71e-12
+  mcm4m1l1_ca_w_0_140_s_0_175=1.01e-04 mcm4m1l1_cc_w_0_140_s_0_175=8.16e-11 mcm4m1l1_cf_w_0_140_s_0_175=9.44e-12
+  mcm4m1l1_ca_w_0_140_s_0_210=1.01e-04 mcm4m1l1_cc_w_0_140_s_0_210=7.75e-11 mcm4m1l1_cf_w_0_140_s_0_210=1.12e-11
+  mcm4m1l1_ca_w_0_140_s_0_280=1.01e-04 mcm4m1l1_cc_w_0_140_s_0_280=6.80e-11 mcm4m1l1_cf_w_0_140_s_0_280=1.44e-11
+  mcm4m1l1_ca_w_0_140_s_0_350=1.01e-04 mcm4m1l1_cc_w_0_140_s_0_350=5.76e-11 mcm4m1l1_cf_w_0_140_s_0_350=1.74e-11
+  mcm4m1l1_ca_w_0_140_s_0_420=1.01e-04 mcm4m1l1_cc_w_0_140_s_0_420=4.89e-11 mcm4m1l1_cf_w_0_140_s_0_420=2.03e-11
+  mcm4m1l1_ca_w_0_140_s_0_560=1.01e-04 mcm4m1l1_cc_w_0_140_s_0_560=3.66e-11 mcm4m1l1_cf_w_0_140_s_0_560=2.54e-11
+  mcm4m1l1_ca_w_0_140_s_0_840=1.01e-04 mcm4m1l1_cc_w_0_140_s_0_840=2.26e-11 mcm4m1l1_cf_w_0_140_s_0_840=3.35e-11
+  mcm4m1l1_ca_w_0_140_s_1_540=1.01e-04 mcm4m1l1_cc_w_0_140_s_1_540=8.46e-12 mcm4m1l1_cf_w_0_140_s_1_540=4.47e-11
+  mcm4m1l1_ca_w_0_140_s_3_500=1.01e-04 mcm4m1l1_cc_w_0_140_s_3_500=9.85e-13 mcm4m1l1_cf_w_0_140_s_3_500=5.18e-11
+  mcm4m1l1_ca_w_1_120_s_0_140=1.01e-04 mcm4m1l1_cc_w_1_120_s_0_140=9.72e-11 mcm4m1l1_cf_w_1_120_s_0_140=7.81e-12
+  mcm4m1l1_ca_w_1_120_s_0_175=1.01e-04 mcm4m1l1_cc_w_1_120_s_0_175=9.37e-11 mcm4m1l1_cf_w_1_120_s_0_175=9.56e-12
+  mcm4m1l1_ca_w_1_120_s_0_210=1.01e-04 mcm4m1l1_cc_w_1_120_s_0_210=8.94e-11 mcm4m1l1_cf_w_1_120_s_0_210=1.12e-11
+  mcm4m1l1_ca_w_1_120_s_0_280=1.01e-04 mcm4m1l1_cc_w_1_120_s_0_280=7.75e-11 mcm4m1l1_cf_w_1_120_s_0_280=1.45e-11
+  mcm4m1l1_ca_w_1_120_s_0_350=1.01e-04 mcm4m1l1_cc_w_1_120_s_0_350=6.62e-11 mcm4m1l1_cf_w_1_120_s_0_350=1.75e-11
+  mcm4m1l1_ca_w_1_120_s_0_420=1.01e-04 mcm4m1l1_cc_w_1_120_s_0_420=5.69e-11 mcm4m1l1_cf_w_1_120_s_0_420=2.04e-11
+  mcm4m1l1_ca_w_1_120_s_0_560=1.01e-04 mcm4m1l1_cc_w_1_120_s_0_560=4.31e-11 mcm4m1l1_cf_w_1_120_s_0_560=2.55e-11
+  mcm4m1l1_ca_w_1_120_s_0_840=1.01e-04 mcm4m1l1_cc_w_1_120_s_0_840=2.74e-11 mcm4m1l1_cf_w_1_120_s_0_840=3.38e-11
+  mcm4m1l1_ca_w_1_120_s_1_540=1.01e-04 mcm4m1l1_cc_w_1_120_s_1_540=1.11e-11 mcm4m1l1_cf_w_1_120_s_1_540=4.60e-11
+  mcm4m1l1_ca_w_1_120_s_3_500=1.01e-04 mcm4m1l1_cc_w_1_120_s_3_500=1.46e-12 mcm4m1l1_cf_w_1_120_s_3_500=5.51e-11
+  mcm5m1f_ca_w_0_140_s_0_140=3.03e-05 mcm5m1f_cc_w_0_140_s_0_140=9.13e-11 mcm5m1f_cf_w_0_140_s_0_140=2.43e-12
+  mcm5m1f_ca_w_0_140_s_0_175=3.03e-05 mcm5m1f_cc_w_0_140_s_0_175=9.09e-11 mcm5m1f_cf_w_0_140_s_0_175=2.95e-12
+  mcm5m1f_ca_w_0_140_s_0_210=3.03e-05 mcm5m1f_cc_w_0_140_s_0_210=8.63e-11 mcm5m1f_cf_w_0_140_s_0_210=3.49e-12
+  mcm5m1f_ca_w_0_140_s_0_280=3.03e-05 mcm5m1f_cc_w_0_140_s_0_280=7.82e-11 mcm5m1f_cf_w_0_140_s_0_280=4.51e-12
+  mcm5m1f_ca_w_0_140_s_0_350=3.03e-05 mcm5m1f_cc_w_0_140_s_0_350=6.84e-11 mcm5m1f_cf_w_0_140_s_0_350=5.52e-12
+  mcm5m1f_ca_w_0_140_s_0_420=3.03e-05 mcm5m1f_cc_w_0_140_s_0_420=6.03e-11 mcm5m1f_cf_w_0_140_s_0_420=6.58e-12
+  mcm5m1f_ca_w_0_140_s_0_560=3.03e-05 mcm5m1f_cc_w_0_140_s_0_560=4.92e-11 mcm5m1f_cf_w_0_140_s_0_560=8.50e-12
+  mcm5m1f_ca_w_0_140_s_0_840=3.03e-05 mcm5m1f_cc_w_0_140_s_0_840=3.61e-11 mcm5m1f_cf_w_0_140_s_0_840=1.21e-11
+  mcm5m1f_ca_w_0_140_s_1_540=3.03e-05 mcm5m1f_cc_w_0_140_s_1_540=2.02e-11 mcm5m1f_cf_w_0_140_s_1_540=1.95e-11
+  mcm5m1f_ca_w_0_140_s_3_500=3.03e-05 mcm5m1f_cc_w_0_140_s_3_500=5.72e-12 mcm5m1f_cf_w_0_140_s_3_500=3.02e-11
+  mcm5m1f_ca_w_1_120_s_0_140=3.03e-05 mcm5m1f_cc_w_1_120_s_0_140=1.15e-10 mcm5m1f_cf_w_1_120_s_0_140=2.46e-12
+  mcm5m1f_ca_w_1_120_s_0_175=3.03e-05 mcm5m1f_cc_w_1_120_s_0_175=1.11e-10 mcm5m1f_cf_w_1_120_s_0_175=2.99e-12
+  mcm5m1f_ca_w_1_120_s_0_210=3.03e-05 mcm5m1f_cc_w_1_120_s_0_210=1.07e-10 mcm5m1f_cf_w_1_120_s_0_210=3.50e-12
+  mcm5m1f_ca_w_1_120_s_0_280=3.03e-05 mcm5m1f_cc_w_1_120_s_0_280=9.54e-11 mcm5m1f_cf_w_1_120_s_0_280=4.55e-12
+  mcm5m1f_ca_w_1_120_s_0_350=3.03e-05 mcm5m1f_cc_w_1_120_s_0_350=8.41e-11 mcm5m1f_cf_w_1_120_s_0_350=5.58e-12
+  mcm5m1f_ca_w_1_120_s_0_420=3.03e-05 mcm5m1f_cc_w_1_120_s_0_420=7.45e-11 mcm5m1f_cf_w_1_120_s_0_420=6.59e-12
+  mcm5m1f_ca_w_1_120_s_0_560=3.03e-05 mcm5m1f_cc_w_1_120_s_0_560=6.12e-11 mcm5m1f_cf_w_1_120_s_0_560=8.53e-12
+  mcm5m1f_ca_w_1_120_s_0_840=3.03e-05 mcm5m1f_cc_w_1_120_s_0_840=4.48e-11 mcm5m1f_cf_w_1_120_s_0_840=1.22e-11
+  mcm5m1f_ca_w_1_120_s_1_540=3.03e-05 mcm5m1f_cc_w_1_120_s_1_540=2.55e-11 mcm5m1f_cf_w_1_120_s_1_540=2.00e-11
+  mcm5m1f_ca_w_1_120_s_3_500=3.03e-05 mcm5m1f_cc_w_1_120_s_3_500=7.62e-12 mcm5m1f_cf_w_1_120_s_3_500=3.24e-11
+  mcm5m1d_ca_w_0_140_s_0_140=3.72e-05 mcm5m1d_cc_w_0_140_s_0_140=9.05e-11 mcm5m1d_cf_w_0_140_s_0_140=2.97e-12
+  mcm5m1d_ca_w_0_140_s_0_175=3.72e-05 mcm5m1d_cc_w_0_140_s_0_175=9.00e-11 mcm5m1d_cf_w_0_140_s_0_175=3.61e-12
+  mcm5m1d_ca_w_0_140_s_0_210=3.72e-05 mcm5m1d_cc_w_0_140_s_0_210=8.53e-11 mcm5m1d_cf_w_0_140_s_0_210=4.27e-12
+  mcm5m1d_ca_w_0_140_s_0_280=3.72e-05 mcm5m1d_cc_w_0_140_s_0_280=7.68e-11 mcm5m1d_cf_w_0_140_s_0_280=5.51e-12
+  mcm5m1d_ca_w_0_140_s_0_350=3.72e-05 mcm5m1d_cc_w_0_140_s_0_350=6.68e-11 mcm5m1d_cf_w_0_140_s_0_350=6.74e-12
+  mcm5m1d_ca_w_0_140_s_0_420=3.72e-05 mcm5m1d_cc_w_0_140_s_0_420=5.90e-11 mcm5m1d_cf_w_0_140_s_0_420=8.02e-12
+  mcm5m1d_ca_w_0_140_s_0_560=3.72e-05 mcm5m1d_cc_w_0_140_s_0_560=4.74e-11 mcm5m1d_cf_w_0_140_s_0_560=1.03e-11
+  mcm5m1d_ca_w_0_140_s_0_840=3.72e-05 mcm5m1d_cc_w_0_140_s_0_840=3.41e-11 mcm5m1d_cf_w_0_140_s_0_840=1.46e-11
+  mcm5m1d_ca_w_0_140_s_1_540=3.72e-05 mcm5m1d_cc_w_0_140_s_1_540=1.80e-11 mcm5m1d_cf_w_0_140_s_1_540=2.29e-11
+  mcm5m1d_ca_w_0_140_s_3_500=3.72e-05 mcm5m1d_cc_w_0_140_s_3_500=4.46e-12 mcm5m1d_cf_w_0_140_s_3_500=3.35e-11
+  mcm5m1d_ca_w_1_120_s_0_140=3.72e-05 mcm5m1d_cc_w_1_120_s_0_140=1.12e-10 mcm5m1d_cf_w_1_120_s_0_140=3.02e-12
+  mcm5m1d_ca_w_1_120_s_0_175=3.72e-05 mcm5m1d_cc_w_1_120_s_0_175=1.08e-10 mcm5m1d_cf_w_1_120_s_0_175=3.66e-12
+  mcm5m1d_ca_w_1_120_s_0_210=3.72e-05 mcm5m1d_cc_w_1_120_s_0_210=1.05e-10 mcm5m1d_cf_w_1_120_s_0_210=4.30e-12
+  mcm5m1d_ca_w_1_120_s_0_280=3.72e-05 mcm5m1d_cc_w_1_120_s_0_280=9.27e-11 mcm5m1d_cf_w_1_120_s_0_280=5.57e-12
+  mcm5m1d_ca_w_1_120_s_0_350=3.72e-05 mcm5m1d_cc_w_1_120_s_0_350=8.16e-11 mcm5m1d_cf_w_1_120_s_0_350=6.82e-12
+  mcm5m1d_ca_w_1_120_s_0_420=3.72e-05 mcm5m1d_cc_w_1_120_s_0_420=7.22e-11 mcm5m1d_cf_w_1_120_s_0_420=8.04e-12
+  mcm5m1d_ca_w_1_120_s_0_560=3.72e-05 mcm5m1d_cc_w_1_120_s_0_560=5.83e-11 mcm5m1d_cf_w_1_120_s_0_560=1.04e-11
+  mcm5m1d_ca_w_1_120_s_0_840=3.72e-05 mcm5m1d_cc_w_1_120_s_0_840=4.19e-11 mcm5m1d_cf_w_1_120_s_0_840=1.48e-11
+  mcm5m1d_ca_w_1_120_s_1_540=3.72e-05 mcm5m1d_cc_w_1_120_s_1_540=2.28e-11 mcm5m1d_cf_w_1_120_s_1_540=2.36e-11
+  mcm5m1d_ca_w_1_120_s_3_500=3.72e-05 mcm5m1d_cc_w_1_120_s_3_500=6.06e-12 mcm5m1d_cf_w_1_120_s_3_500=3.61e-11
+  mcm5m1p1_ca_w_0_140_s_0_140=4.42e-05 mcm5m1p1_cc_w_0_140_s_0_140=8.97e-11 mcm5m1p1_cf_w_0_140_s_0_140=3.52e-12
+  mcm5m1p1_ca_w_0_140_s_0_175=4.42e-05 mcm5m1p1_cc_w_0_140_s_0_175=8.91e-11 mcm5m1p1_cf_w_0_140_s_0_175=4.28e-12
+  mcm5m1p1_ca_w_0_140_s_0_210=4.42e-05 mcm5m1p1_cc_w_0_140_s_0_210=8.44e-11 mcm5m1p1_cf_w_0_140_s_0_210=5.06e-12
+  mcm5m1p1_ca_w_0_140_s_0_280=4.42e-05 mcm5m1p1_cc_w_0_140_s_0_280=7.54e-11 mcm5m1p1_cf_w_0_140_s_0_280=6.55e-12
+  mcm5m1p1_ca_w_0_140_s_0_350=4.42e-05 mcm5m1p1_cc_w_0_140_s_0_350=6.59e-11 mcm5m1p1_cf_w_0_140_s_0_350=8.00e-12
+  mcm5m1p1_ca_w_0_140_s_0_420=4.42e-05 mcm5m1p1_cc_w_0_140_s_0_420=5.76e-11 mcm5m1p1_cf_w_0_140_s_0_420=9.47e-12
+  mcm5m1p1_ca_w_0_140_s_0_560=4.42e-05 mcm5m1p1_cc_w_0_140_s_0_560=4.59e-11 mcm5m1p1_cf_w_0_140_s_0_560=1.22e-11
+  mcm5m1p1_ca_w_0_140_s_0_840=4.42e-05 mcm5m1p1_cc_w_0_140_s_0_840=3.22e-11 mcm5m1p1_cf_w_0_140_s_0_840=1.70e-11
+  mcm5m1p1_ca_w_0_140_s_1_540=4.42e-05 mcm5m1p1_cc_w_0_140_s_1_540=1.63e-11 mcm5m1p1_cf_w_0_140_s_1_540=2.61e-11
+  mcm5m1p1_ca_w_0_140_s_3_500=4.42e-05 mcm5m1p1_cc_w_0_140_s_3_500=3.63e-12 mcm5m1p1_cf_w_0_140_s_3_500=3.65e-11
+  mcm5m1p1_ca_w_1_120_s_0_140=4.42e-05 mcm5m1p1_cc_w_1_120_s_0_140=1.10e-10 mcm5m1p1_cf_w_1_120_s_0_140=3.64e-12
+  mcm5m1p1_ca_w_1_120_s_0_175=4.42e-05 mcm5m1p1_cc_w_1_120_s_0_175=1.06e-10 mcm5m1p1_cf_w_1_120_s_0_175=4.40e-12
+  mcm5m1p1_ca_w_1_120_s_0_210=4.42e-05 mcm5m1p1_cc_w_1_120_s_0_210=1.02e-10 mcm5m1p1_cf_w_1_120_s_0_210=5.15e-12
+  mcm5m1p1_ca_w_1_120_s_0_280=4.42e-05 mcm5m1p1_cc_w_1_120_s_0_280=9.04e-11 mcm5m1p1_cf_w_1_120_s_0_280=6.65e-12
+  mcm5m1p1_ca_w_1_120_s_0_350=4.42e-05 mcm5m1p1_cc_w_1_120_s_0_350=7.91e-11 mcm5m1p1_cf_w_1_120_s_0_350=8.12e-12
+  mcm5m1p1_ca_w_1_120_s_0_420=4.42e-05 mcm5m1p1_cc_w_1_120_s_0_420=6.97e-11 mcm5m1p1_cf_w_1_120_s_0_420=9.54e-12
+  mcm5m1p1_ca_w_1_120_s_0_560=4.42e-05 mcm5m1p1_cc_w_1_120_s_0_560=5.59e-11 mcm5m1p1_cf_w_1_120_s_0_560=1.23e-11
+  mcm5m1p1_ca_w_1_120_s_0_840=4.42e-05 mcm5m1p1_cc_w_1_120_s_0_840=3.95e-11 mcm5m1p1_cf_w_1_120_s_0_840=1.73e-11
+  mcm5m1p1_ca_w_1_120_s_1_540=4.42e-05 mcm5m1p1_cc_w_1_120_s_1_540=2.07e-11 mcm5m1p1_cf_w_1_120_s_1_540=2.69e-11
+  mcm5m1p1_ca_w_1_120_s_3_500=4.42e-05 mcm5m1p1_cc_w_1_120_s_3_500=5.08e-12 mcm5m1p1_cf_w_1_120_s_3_500=3.92e-11
+  mcm5m1l1_ca_w_0_140_s_0_140=9.59e-05 mcm5m1l1_cc_w_0_140_s_0_140=8.43e-11 mcm5m1l1_cf_w_0_140_s_0_140=7.32e-12
+  mcm5m1l1_ca_w_0_140_s_0_175=9.59e-05 mcm5m1l1_cc_w_0_140_s_0_175=8.30e-11 mcm5m1l1_cf_w_0_140_s_0_175=8.98e-12
+  mcm5m1l1_ca_w_0_140_s_0_210=9.59e-05 mcm5m1l1_cc_w_0_140_s_0_210=7.83e-11 mcm5m1l1_cf_w_0_140_s_0_210=1.06e-11
+  mcm5m1l1_ca_w_0_140_s_0_280=9.59e-05 mcm5m1l1_cc_w_0_140_s_0_280=6.89e-11 mcm5m1l1_cf_w_0_140_s_0_280=1.37e-11
+  mcm5m1l1_ca_w_0_140_s_0_350=9.59e-05 mcm5m1l1_cc_w_0_140_s_0_350=5.86e-11 mcm5m1l1_cf_w_0_140_s_0_350=1.65e-11
+  mcm5m1l1_ca_w_0_140_s_0_420=9.59e-05 mcm5m1l1_cc_w_0_140_s_0_420=5.00e-11 mcm5m1l1_cf_w_0_140_s_0_420=1.93e-11
+  mcm5m1l1_ca_w_0_140_s_0_560=9.59e-05 mcm5m1l1_cc_w_0_140_s_0_560=3.78e-11 mcm5m1l1_cf_w_0_140_s_0_560=2.42e-11
+  mcm5m1l1_ca_w_0_140_s_0_840=9.59e-05 mcm5m1l1_cc_w_0_140_s_0_840=2.41e-11 mcm5m1l1_cf_w_0_140_s_0_840=3.19e-11
+  mcm5m1l1_ca_w_0_140_s_1_540=9.59e-05 mcm5m1l1_cc_w_0_140_s_1_540=9.91e-12 mcm5m1l1_cf_w_0_140_s_1_540=4.30e-11
+  mcm5m1l1_ca_w_0_140_s_3_500=9.59e-05 mcm5m1l1_cc_w_0_140_s_3_500=1.65e-12 mcm5m1l1_cf_w_0_140_s_3_500=5.08e-11
+  mcm5m1l1_ca_w_1_120_s_0_140=9.59e-05 mcm5m1l1_cc_w_1_120_s_0_140=9.95e-11 mcm5m1l1_cf_w_1_120_s_0_140=7.45e-12
+  mcm5m1l1_ca_w_1_120_s_0_175=9.59e-05 mcm5m1l1_cc_w_1_120_s_0_175=9.63e-11 mcm5m1l1_cf_w_1_120_s_0_175=9.10e-12
+  mcm5m1l1_ca_w_1_120_s_0_210=9.59e-05 mcm5m1l1_cc_w_1_120_s_0_210=9.18e-11 mcm5m1l1_cf_w_1_120_s_0_210=1.07e-11
+  mcm5m1l1_ca_w_1_120_s_0_280=9.59e-05 mcm5m1l1_cc_w_1_120_s_0_280=8.00e-11 mcm5m1l1_cf_w_1_120_s_0_280=1.38e-11
+  mcm5m1l1_ca_w_1_120_s_0_350=9.59e-05 mcm5m1l1_cc_w_1_120_s_0_350=6.89e-11 mcm5m1l1_cf_w_1_120_s_0_350=1.67e-11
+  mcm5m1l1_ca_w_1_120_s_0_420=9.59e-05 mcm5m1l1_cc_w_1_120_s_0_420=5.93e-11 mcm5m1l1_cf_w_1_120_s_0_420=1.94e-11
+  mcm5m1l1_ca_w_1_120_s_0_560=9.59e-05 mcm5m1l1_cc_w_1_120_s_0_560=4.59e-11 mcm5m1l1_cf_w_1_120_s_0_560=2.43e-11
+  mcm5m1l1_ca_w_1_120_s_0_840=9.59e-05 mcm5m1l1_cc_w_1_120_s_0_840=3.04e-11 mcm5m1l1_cf_w_1_120_s_0_840=3.22e-11
+  mcm5m1l1_ca_w_1_120_s_1_540=9.59e-05 mcm5m1l1_cc_w_1_120_s_1_540=1.38e-11 mcm5m1l1_cf_w_1_120_s_1_540=4.43e-11
+  mcm5m1l1_ca_w_1_120_s_3_500=9.59e-05 mcm5m1l1_cc_w_1_120_s_3_500=2.66e-12 mcm5m1l1_cf_w_1_120_s_3_500=5.45e-11
+  mcrdlm1f_ca_w_0_140_s_0_140=2.43e-05 mcrdlm1f_cc_w_0_140_s_0_140=9.20e-11 mcrdlm1f_cf_w_0_140_s_0_140=1.94e-12
+  mcrdlm1f_ca_w_0_140_s_0_175=2.43e-05 mcrdlm1f_cc_w_0_140_s_0_175=9.07e-11 mcrdlm1f_cf_w_0_140_s_0_175=2.36e-12
+  mcrdlm1f_ca_w_0_140_s_0_210=2.43e-05 mcrdlm1f_cc_w_0_140_s_0_210=8.67e-11 mcrdlm1f_cf_w_0_140_s_0_210=2.80e-12
+  mcrdlm1f_ca_w_0_140_s_0_280=2.43e-05 mcrdlm1f_cc_w_0_140_s_0_280=7.88e-11 mcrdlm1f_cf_w_0_140_s_0_280=3.62e-12
+  mcrdlm1f_ca_w_0_140_s_0_350=2.43e-05 mcrdlm1f_cc_w_0_140_s_0_350=6.92e-11 mcrdlm1f_cf_w_0_140_s_0_350=4.43e-12
+  mcrdlm1f_ca_w_0_140_s_0_420=2.43e-05 mcrdlm1f_cc_w_0_140_s_0_420=6.16e-11 mcrdlm1f_cf_w_0_140_s_0_420=5.27e-12
+  mcrdlm1f_ca_w_0_140_s_0_560=2.43e-05 mcrdlm1f_cc_w_0_140_s_0_560=5.08e-11 mcrdlm1f_cf_w_0_140_s_0_560=6.84e-12
+  mcrdlm1f_ca_w_0_140_s_0_840=2.43e-05 mcrdlm1f_cc_w_0_140_s_0_840=3.82e-11 mcrdlm1f_cf_w_0_140_s_0_840=9.75e-12
+  mcrdlm1f_ca_w_0_140_s_1_540=2.43e-05 mcrdlm1f_cc_w_0_140_s_1_540=2.33e-11 mcrdlm1f_cf_w_0_140_s_1_540=1.60e-11
+  mcrdlm1f_ca_w_0_140_s_3_500=2.43e-05 mcrdlm1f_cc_w_0_140_s_3_500=8.88e-12 mcrdlm1f_cf_w_0_140_s_3_500=2.62e-11
+  mcrdlm1f_ca_w_1_120_s_0_140=2.43e-05 mcrdlm1f_cc_w_1_120_s_0_140=1.18e-10 mcrdlm1f_cf_w_1_120_s_0_140=1.98e-12
+  mcrdlm1f_ca_w_1_120_s_0_175=2.43e-05 mcrdlm1f_cc_w_1_120_s_0_175=1.14e-10 mcrdlm1f_cf_w_1_120_s_0_175=2.40e-12
+  mcrdlm1f_ca_w_1_120_s_0_210=2.43e-05 mcrdlm1f_cc_w_1_120_s_0_210=1.11e-10 mcrdlm1f_cf_w_1_120_s_0_210=2.82e-12
+  mcrdlm1f_ca_w_1_120_s_0_280=2.43e-05 mcrdlm1f_cc_w_1_120_s_0_280=9.89e-11 mcrdlm1f_cf_w_1_120_s_0_280=3.66e-12
+  mcrdlm1f_ca_w_1_120_s_0_350=2.43e-05 mcrdlm1f_cc_w_1_120_s_0_350=8.78e-11 mcrdlm1f_cf_w_1_120_s_0_350=4.48e-12
+  mcrdlm1f_ca_w_1_120_s_0_420=2.43e-05 mcrdlm1f_cc_w_1_120_s_0_420=7.86e-11 mcrdlm1f_cf_w_1_120_s_0_420=5.29e-12
+  mcrdlm1f_ca_w_1_120_s_0_560=2.43e-05 mcrdlm1f_cc_w_1_120_s_0_560=6.52e-11 mcrdlm1f_cf_w_1_120_s_0_560=6.87e-12
+  mcrdlm1f_ca_w_1_120_s_0_840=2.43e-05 mcrdlm1f_cc_w_1_120_s_0_840=4.93e-11 mcrdlm1f_cf_w_1_120_s_0_840=9.86e-12
+  mcrdlm1f_ca_w_1_120_s_1_540=2.43e-05 mcrdlm1f_cc_w_1_120_s_1_540=3.09e-11 mcrdlm1f_cf_w_1_120_s_1_540=1.64e-11
+  mcrdlm1f_ca_w_1_120_s_3_500=2.43e-05 mcrdlm1f_cc_w_1_120_s_3_500=1.26e-11 mcrdlm1f_cf_w_1_120_s_3_500=2.80e-11
+  mcrdlm1d_ca_w_0_140_s_0_140=3.12e-05 mcrdlm1d_cc_w_0_140_s_0_140=9.12e-11 mcrdlm1d_cf_w_0_140_s_0_140=2.49e-12
+  mcrdlm1d_ca_w_0_140_s_0_175=3.12e-05 mcrdlm1d_cc_w_0_140_s_0_175=8.98e-11 mcrdlm1d_cf_w_0_140_s_0_175=3.03e-12
+  mcrdlm1d_ca_w_0_140_s_0_210=3.12e-05 mcrdlm1d_cc_w_0_140_s_0_210=8.57e-11 mcrdlm1d_cf_w_0_140_s_0_210=3.58e-12
+  mcrdlm1d_ca_w_0_140_s_0_280=3.12e-05 mcrdlm1d_cc_w_0_140_s_0_280=7.77e-11 mcrdlm1d_cf_w_0_140_s_0_280=4.63e-12
+  mcrdlm1d_ca_w_0_140_s_0_350=3.12e-05 mcrdlm1d_cc_w_0_140_s_0_350=6.79e-11 mcrdlm1d_cf_w_0_140_s_0_350=5.66e-12
+  mcrdlm1d_ca_w_0_140_s_0_420=3.12e-05 mcrdlm1d_cc_w_0_140_s_0_420=6.01e-11 mcrdlm1d_cf_w_0_140_s_0_420=6.71e-12
+  mcrdlm1d_ca_w_0_140_s_0_560=3.12e-05 mcrdlm1d_cc_w_0_140_s_0_560=4.91e-11 mcrdlm1d_cf_w_0_140_s_0_560=8.67e-12
+  mcrdlm1d_ca_w_0_140_s_0_840=3.12e-05 mcrdlm1d_cc_w_0_140_s_0_840=3.63e-11 mcrdlm1d_cf_w_0_140_s_0_840=1.22e-11
+  mcrdlm1d_ca_w_0_140_s_1_540=3.12e-05 mcrdlm1d_cc_w_0_140_s_1_540=2.10e-11 mcrdlm1d_cf_w_0_140_s_1_540=1.96e-11
+  mcrdlm1d_ca_w_0_140_s_3_500=3.12e-05 mcrdlm1d_cc_w_0_140_s_3_500=7.18e-12 mcrdlm1d_cf_w_0_140_s_3_500=3.02e-11
+  mcrdlm1d_ca_w_1_120_s_0_140=3.12e-05 mcrdlm1d_cc_w_1_120_s_0_140=1.15e-10 mcrdlm1d_cf_w_1_120_s_0_140=2.54e-12
+  mcrdlm1d_ca_w_1_120_s_0_175=3.12e-05 mcrdlm1d_cc_w_1_120_s_0_175=1.12e-10 mcrdlm1d_cf_w_1_120_s_0_175=3.09e-12
+  mcrdlm1d_ca_w_1_120_s_0_210=3.12e-05 mcrdlm1d_cc_w_1_120_s_0_210=1.08e-10 mcrdlm1d_cf_w_1_120_s_0_210=3.62e-12
+  mcrdlm1d_ca_w_1_120_s_0_280=3.12e-05 mcrdlm1d_cc_w_1_120_s_0_280=9.62e-11 mcrdlm1d_cf_w_1_120_s_0_280=4.69e-12
+  mcrdlm1d_ca_w_1_120_s_0_350=3.12e-05 mcrdlm1d_cc_w_1_120_s_0_350=8.51e-11 mcrdlm1d_cf_w_1_120_s_0_350=5.73e-12
+  mcrdlm1d_ca_w_1_120_s_0_420=3.12e-05 mcrdlm1d_cc_w_1_120_s_0_420=7.57e-11 mcrdlm1d_cf_w_1_120_s_0_420=6.76e-12
+  mcrdlm1d_ca_w_1_120_s_0_560=3.12e-05 mcrdlm1d_cc_w_1_120_s_0_560=6.23e-11 mcrdlm1d_cf_w_1_120_s_0_560=8.74e-12
+  mcrdlm1d_ca_w_1_120_s_0_840=3.12e-05 mcrdlm1d_cc_w_1_120_s_0_840=4.65e-11 mcrdlm1d_cf_w_1_120_s_0_840=1.24e-11
+  mcrdlm1d_ca_w_1_120_s_1_540=3.12e-05 mcrdlm1d_cc_w_1_120_s_1_540=2.80e-11 mcrdlm1d_cf_w_1_120_s_1_540=2.02e-11
+  mcrdlm1d_ca_w_1_120_s_3_500=3.12e-05 mcrdlm1d_cc_w_1_120_s_3_500=1.06e-11 mcrdlm1d_cf_w_1_120_s_3_500=3.25e-11
+  mcrdlm1p1_ca_w_0_140_s_0_140=3.81e-05 mcrdlm1p1_cc_w_0_140_s_0_140=9.04e-11 mcrdlm1p1_cf_w_0_140_s_0_140=3.04e-12
+  mcrdlm1p1_ca_w_0_140_s_0_175=3.81e-05 mcrdlm1p1_cc_w_0_140_s_0_175=8.90e-11 mcrdlm1p1_cf_w_0_140_s_0_175=3.70e-12
+  mcrdlm1p1_ca_w_0_140_s_0_210=3.81e-05 mcrdlm1p1_cc_w_0_140_s_0_210=8.47e-11 mcrdlm1p1_cf_w_0_140_s_0_210=4.36e-12
+  mcrdlm1p1_ca_w_0_140_s_0_280=3.81e-05 mcrdlm1p1_cc_w_0_140_s_0_280=7.66e-11 mcrdlm1p1_cf_w_0_140_s_0_280=5.65e-12
+  mcrdlm1p1_ca_w_0_140_s_0_350=3.81e-05 mcrdlm1p1_cc_w_0_140_s_0_350=6.67e-11 mcrdlm1p1_cf_w_0_140_s_0_350=6.90e-12
+  mcrdlm1p1_ca_w_0_140_s_0_420=3.81e-05 mcrdlm1p1_cc_w_0_140_s_0_420=5.86e-11 mcrdlm1p1_cf_w_0_140_s_0_420=8.15e-12
+  mcrdlm1p1_ca_w_0_140_s_0_560=3.81e-05 mcrdlm1p1_cc_w_0_140_s_0_560=4.76e-11 mcrdlm1p1_cf_w_0_140_s_0_560=1.05e-11
+  mcrdlm1p1_ca_w_0_140_s_0_840=3.81e-05 mcrdlm1p1_cc_w_0_140_s_0_840=3.44e-11 mcrdlm1p1_cf_w_0_140_s_0_840=1.47e-11
+  mcrdlm1p1_ca_w_0_140_s_1_540=3.81e-05 mcrdlm1p1_cc_w_0_140_s_1_540=1.91e-11 mcrdlm1p1_cf_w_0_140_s_1_540=2.30e-11
+  mcrdlm1p1_ca_w_0_140_s_3_500=3.81e-05 mcrdlm1p1_cc_w_0_140_s_3_500=6.01e-12 mcrdlm1p1_cf_w_0_140_s_3_500=3.36e-11
+  mcrdlm1p1_ca_w_1_120_s_0_140=3.81e-05 mcrdlm1p1_cc_w_1_120_s_0_140=1.13e-10 mcrdlm1p1_cf_w_1_120_s_0_140=3.15e-12
+  mcrdlm1p1_ca_w_1_120_s_0_175=3.81e-05 mcrdlm1p1_cc_w_1_120_s_0_175=1.10e-10 mcrdlm1p1_cf_w_1_120_s_0_175=3.82e-12
+  mcrdlm1p1_ca_w_1_120_s_0_210=3.81e-05 mcrdlm1p1_cc_w_1_120_s_0_210=1.05e-10 mcrdlm1p1_cf_w_1_120_s_0_210=4.45e-12
+  mcrdlm1p1_ca_w_1_120_s_0_280=3.81e-05 mcrdlm1p1_cc_w_1_120_s_0_280=9.37e-11 mcrdlm1p1_cf_w_1_120_s_0_280=5.76e-12
+  mcrdlm1p1_ca_w_1_120_s_0_350=3.81e-05 mcrdlm1p1_cc_w_1_120_s_0_350=8.26e-11 mcrdlm1p1_cf_w_1_120_s_0_350=7.02e-12
+  mcrdlm1p1_ca_w_1_120_s_0_420=3.81e-05 mcrdlm1p1_cc_w_1_120_s_0_420=7.33e-11 mcrdlm1p1_cf_w_1_120_s_0_420=8.26e-12
+  mcrdlm1p1_ca_w_1_120_s_0_560=3.81e-05 mcrdlm1p1_cc_w_1_120_s_0_560=5.98e-11 mcrdlm1p1_cf_w_1_120_s_0_560=1.06e-11
+  mcrdlm1p1_ca_w_1_120_s_0_840=3.81e-05 mcrdlm1p1_cc_w_1_120_s_0_840=4.42e-11 mcrdlm1p1_cf_w_1_120_s_0_840=1.49e-11
+  mcrdlm1p1_ca_w_1_120_s_1_540=3.81e-05 mcrdlm1p1_cc_w_1_120_s_1_540=2.58e-11 mcrdlm1p1_cf_w_1_120_s_1_540=2.36e-11
+  mcrdlm1p1_ca_w_1_120_s_3_500=3.81e-05 mcrdlm1p1_cc_w_1_120_s_3_500=9.23e-12 mcrdlm1p1_cf_w_1_120_s_3_500=3.62e-11
+  mcrdlm1l1_ca_w_0_140_s_0_140=8.99e-05 mcrdlm1l1_cc_w_0_140_s_0_140=8.50e-11 mcrdlm1l1_cf_w_0_140_s_0_140=6.84e-12
+  mcrdlm1l1_ca_w_0_140_s_0_175=8.99e-05 mcrdlm1l1_cc_w_0_140_s_0_175=8.36e-11 mcrdlm1l1_cf_w_0_140_s_0_175=8.40e-12
+  mcrdlm1l1_ca_w_0_140_s_0_210=8.99e-05 mcrdlm1l1_cc_w_0_140_s_0_210=7.92e-11 mcrdlm1l1_cf_w_0_140_s_0_210=9.94e-12
+  mcrdlm1l1_ca_w_0_140_s_0_280=8.99e-05 mcrdlm1l1_cc_w_0_140_s_0_280=6.99e-11 mcrdlm1l1_cf_w_0_140_s_0_280=1.28e-11
+  mcrdlm1l1_ca_w_0_140_s_0_350=8.99e-05 mcrdlm1l1_cc_w_0_140_s_0_350=5.95e-11 mcrdlm1l1_cf_w_0_140_s_0_350=1.54e-11
+  mcrdlm1l1_ca_w_0_140_s_0_420=8.99e-05 mcrdlm1l1_cc_w_0_140_s_0_420=5.11e-11 mcrdlm1l1_cf_w_0_140_s_0_420=1.80e-11
+  mcrdlm1l1_ca_w_0_140_s_0_560=8.99e-05 mcrdlm1l1_cc_w_0_140_s_0_560=3.95e-11 mcrdlm1l1_cf_w_0_140_s_0_560=2.26e-11
+  mcrdlm1l1_ca_w_0_140_s_0_840=8.99e-05 mcrdlm1l1_cc_w_0_140_s_0_840=2.62e-11 mcrdlm1l1_cf_w_0_140_s_0_840=2.98e-11
+  mcrdlm1l1_ca_w_0_140_s_1_540=8.99e-05 mcrdlm1l1_cc_w_0_140_s_1_540=1.21e-11 mcrdlm1l1_cf_w_0_140_s_1_540=4.07e-11
+  mcrdlm1l1_ca_w_0_140_s_3_500=8.99e-05 mcrdlm1l1_cc_w_0_140_s_3_500=3.03e-12 mcrdlm1l1_cf_w_0_140_s_3_500=4.94e-11
+  mcrdlm1l1_ca_w_1_120_s_0_140=8.99e-05 mcrdlm1l1_cc_w_1_120_s_0_140=1.02e-10 mcrdlm1l1_cf_w_1_120_s_0_140=6.96e-12
+  mcrdlm1l1_ca_w_1_120_s_0_175=8.99e-05 mcrdlm1l1_cc_w_1_120_s_0_175=1.00e-10 mcrdlm1l1_cf_w_1_120_s_0_175=8.52e-12
+  mcrdlm1l1_ca_w_1_120_s_0_210=8.99e-05 mcrdlm1l1_cc_w_1_120_s_0_210=9.51e-11 mcrdlm1l1_cf_w_1_120_s_0_210=1.00e-11
+  mcrdlm1l1_ca_w_1_120_s_0_280=8.99e-05 mcrdlm1l1_cc_w_1_120_s_0_280=8.35e-11 mcrdlm1l1_cf_w_1_120_s_0_280=1.29e-11
+  mcrdlm1l1_ca_w_1_120_s_0_350=8.99e-05 mcrdlm1l1_cc_w_1_120_s_0_350=7.27e-11 mcrdlm1l1_cf_w_1_120_s_0_350=1.56e-11
+  mcrdlm1l1_ca_w_1_120_s_0_420=8.99e-05 mcrdlm1l1_cc_w_1_120_s_0_420=6.32e-11 mcrdlm1l1_cf_w_1_120_s_0_420=1.81e-11
+  mcrdlm1l1_ca_w_1_120_s_0_560=8.99e-05 mcrdlm1l1_cc_w_1_120_s_0_560=4.99e-11 mcrdlm1l1_cf_w_1_120_s_0_560=2.26e-11
+  mcrdlm1l1_ca_w_1_120_s_0_840=8.99e-05 mcrdlm1l1_cc_w_1_120_s_0_840=3.48e-11 mcrdlm1l1_cf_w_1_120_s_0_840=3.02e-11
+  mcrdlm1l1_ca_w_1_120_s_1_540=8.99e-05 mcrdlm1l1_cc_w_1_120_s_1_540=1.83e-11 mcrdlm1l1_cf_w_1_120_s_1_540=4.18e-11
+  mcrdlm1l1_ca_w_1_120_s_3_500=8.99e-05 mcrdlm1l1_cc_w_1_120_s_3_500=5.53e-12 mcrdlm1l1_cf_w_1_120_s_3_500=5.33e-11
+  mcm3m2f_ca_w_0_140_s_0_140=7.98e-05 mcm3m2f_cc_w_0_140_s_0_140=8.54e-11 mcm3m2f_cf_w_0_140_s_0_140=6.07e-12
+  mcm3m2f_ca_w_0_140_s_0_175=7.98e-05 mcm3m2f_cc_w_0_140_s_0_175=8.44e-11 mcm3m2f_cf_w_0_140_s_0_175=7.33e-12
+  mcm3m2f_ca_w_0_140_s_0_210=7.98e-05 mcm3m2f_cc_w_0_140_s_0_210=8.04e-11 mcm3m2f_cf_w_0_140_s_0_210=8.61e-12
+  mcm3m2f_ca_w_0_140_s_0_280=7.98e-05 mcm3m2f_cc_w_0_140_s_0_280=7.08e-11 mcm3m2f_cf_w_0_140_s_0_280=1.10e-11
+  mcm3m2f_ca_w_0_140_s_0_350=7.98e-05 mcm3m2f_cc_w_0_140_s_0_350=6.06e-11 mcm3m2f_cf_w_0_140_s_0_350=1.33e-11
+  mcm3m2f_ca_w_0_140_s_0_420=7.98e-05 mcm3m2f_cc_w_0_140_s_0_420=5.15e-11 mcm3m2f_cf_w_0_140_s_0_420=1.57e-11
+  mcm3m2f_ca_w_0_140_s_0_560=7.98e-05 mcm3m2f_cc_w_0_140_s_0_560=3.95e-11 mcm3m2f_cf_w_0_140_s_0_560=1.98e-11
+  mcm3m2f_ca_w_0_140_s_0_840=7.98e-05 mcm3m2f_cc_w_0_140_s_0_840=2.52e-11 mcm3m2f_cf_w_0_140_s_0_840=2.66e-11
+  mcm3m2f_ca_w_0_140_s_1_540=7.98e-05 mcm3m2f_cc_w_0_140_s_1_540=1.01e-11 mcm3m2f_cf_w_0_140_s_1_540=3.74e-11
+  mcm3m2f_ca_w_0_140_s_3_500=7.98e-05 mcm3m2f_cc_w_0_140_s_3_500=1.26e-12 mcm3m2f_cf_w_0_140_s_3_500=4.55e-11
+  mcm3m2f_ca_w_1_120_s_0_140=7.98e-05 mcm3m2f_cc_w_1_120_s_0_140=9.99e-11 mcm3m2f_cf_w_1_120_s_0_140=6.12e-12
+  mcm3m2f_ca_w_1_120_s_0_175=7.98e-05 mcm3m2f_cc_w_1_120_s_0_175=9.68e-11 mcm3m2f_cf_w_1_120_s_0_175=7.39e-12
+  mcm3m2f_ca_w_1_120_s_0_210=7.98e-05 mcm3m2f_cc_w_1_120_s_0_210=9.22e-11 mcm3m2f_cf_w_1_120_s_0_210=8.62e-12
+  mcm3m2f_ca_w_1_120_s_0_280=7.98e-05 mcm3m2f_cc_w_1_120_s_0_280=8.04e-11 mcm3m2f_cf_w_1_120_s_0_280=1.11e-11
+  mcm3m2f_ca_w_1_120_s_0_350=7.98e-05 mcm3m2f_cc_w_1_120_s_0_350=6.90e-11 mcm3m2f_cf_w_1_120_s_0_350=1.35e-11
+  mcm3m2f_ca_w_1_120_s_0_420=7.98e-05 mcm3m2f_cc_w_1_120_s_0_420=5.95e-11 mcm3m2f_cf_w_1_120_s_0_420=1.58e-11
+  mcm3m2f_ca_w_1_120_s_0_560=7.98e-05 mcm3m2f_cc_w_1_120_s_0_560=4.57e-11 mcm3m2f_cf_w_1_120_s_0_560=2.00e-11
+  mcm3m2f_ca_w_1_120_s_0_840=7.98e-05 mcm3m2f_cc_w_1_120_s_0_840=2.97e-11 mcm3m2f_cf_w_1_120_s_0_840=2.71e-11
+  mcm3m2f_ca_w_1_120_s_1_540=7.98e-05 mcm3m2f_cc_w_1_120_s_1_540=1.24e-11 mcm3m2f_cf_w_1_120_s_1_540=3.85e-11
+  mcm3m2f_ca_w_1_120_s_3_500=7.98e-05 mcm3m2f_cc_w_1_120_s_3_500=1.62e-12 mcm3m2f_cf_w_1_120_s_3_500=4.83e-11
+  mcm3m2d_ca_w_0_140_s_0_140=8.28e-05 mcm3m2d_cc_w_0_140_s_0_140=8.54e-11 mcm3m2d_cf_w_0_140_s_0_140=6.31e-12
+  mcm3m2d_ca_w_0_140_s_0_175=8.28e-05 mcm3m2d_cc_w_0_140_s_0_175=8.36e-11 mcm3m2d_cf_w_0_140_s_0_175=7.62e-12
+  mcm3m2d_ca_w_0_140_s_0_210=8.28e-05 mcm3m2d_cc_w_0_140_s_0_210=8.00e-11 mcm3m2d_cf_w_0_140_s_0_210=8.95e-12
+  mcm3m2d_ca_w_0_140_s_0_280=8.28e-05 mcm3m2d_cc_w_0_140_s_0_280=7.03e-11 mcm3m2d_cf_w_0_140_s_0_280=1.14e-11
+  mcm3m2d_ca_w_0_140_s_0_350=8.28e-05 mcm3m2d_cc_w_0_140_s_0_350=5.99e-11 mcm3m2d_cf_w_0_140_s_0_350=1.39e-11
+  mcm3m2d_ca_w_0_140_s_0_420=8.28e-05 mcm3m2d_cc_w_0_140_s_0_420=5.09e-11 mcm3m2d_cf_w_0_140_s_0_420=1.63e-11
+  mcm3m2d_ca_w_0_140_s_0_560=8.28e-05 mcm3m2d_cc_w_0_140_s_0_560=3.88e-11 mcm3m2d_cf_w_0_140_s_0_560=2.05e-11
+  mcm3m2d_ca_w_0_140_s_0_840=8.28e-05 mcm3m2d_cc_w_0_140_s_0_840=2.45e-11 mcm3m2d_cf_w_0_140_s_0_840=2.77e-11
+  mcm3m2d_ca_w_0_140_s_1_540=8.28e-05 mcm3m2d_cc_w_0_140_s_1_540=9.24e-12 mcm3m2d_cf_w_0_140_s_1_540=3.85e-11
+  mcm3m2d_ca_w_0_140_s_3_500=8.28e-05 mcm3m2d_cc_w_0_140_s_3_500=9.55e-13 mcm3m2d_cf_w_0_140_s_3_500=4.62e-11
+  mcm3m2d_ca_w_1_120_s_0_140=8.28e-05 mcm3m2d_cc_w_1_120_s_0_140=9.87e-11 mcm3m2d_cf_w_1_120_s_0_140=6.35e-12
+  mcm3m2d_ca_w_1_120_s_0_175=8.28e-05 mcm3m2d_cc_w_1_120_s_0_175=9.55e-11 mcm3m2d_cf_w_1_120_s_0_175=7.69e-12
+  mcm3m2d_ca_w_1_120_s_0_210=8.28e-05 mcm3m2d_cc_w_1_120_s_0_210=9.06e-11 mcm3m2d_cf_w_1_120_s_0_210=8.97e-12
+  mcm3m2d_ca_w_1_120_s_0_280=8.28e-05 mcm3m2d_cc_w_1_120_s_0_280=7.88e-11 mcm3m2d_cf_w_1_120_s_0_280=1.15e-11
+  mcm3m2d_ca_w_1_120_s_0_350=8.28e-05 mcm3m2d_cc_w_1_120_s_0_350=6.76e-11 mcm3m2d_cf_w_1_120_s_0_350=1.40e-11
+  mcm3m2d_ca_w_1_120_s_0_420=8.28e-05 mcm3m2d_cc_w_1_120_s_0_420=5.80e-11 mcm3m2d_cf_w_1_120_s_0_420=1.64e-11
+  mcm3m2d_ca_w_1_120_s_0_560=8.28e-05 mcm3m2d_cc_w_1_120_s_0_560=4.42e-11 mcm3m2d_cf_w_1_120_s_0_560=2.08e-11
+  mcm3m2d_ca_w_1_120_s_0_840=8.28e-05 mcm3m2d_cc_w_1_120_s_0_840=2.80e-11 mcm3m2d_cf_w_1_120_s_0_840=2.81e-11
+  mcm3m2d_ca_w_1_120_s_1_540=8.28e-05 mcm3m2d_cc_w_1_120_s_1_540=1.11e-11 mcm3m2d_cf_w_1_120_s_1_540=3.97e-11
+  mcm3m2d_ca_w_1_120_s_3_500=8.28e-05 mcm3m2d_cc_w_1_120_s_3_500=1.19e-12 mcm3m2d_cf_w_1_120_s_3_500=4.88e-11
+  mcm3m2p1_ca_w_0_140_s_0_140=8.53e-05 mcm3m2p1_cc_w_0_140_s_0_140=8.48e-11 mcm3m2p1_cf_w_0_140_s_0_140=6.52e-12
+  mcm3m2p1_ca_w_0_140_s_0_175=8.53e-05 mcm3m2p1_cc_w_0_140_s_0_175=8.34e-11 mcm3m2p1_cf_w_0_140_s_0_175=7.86e-12
+  mcm3m2p1_ca_w_0_140_s_0_210=8.53e-05 mcm3m2p1_cc_w_0_140_s_0_210=7.96e-11 mcm3m2p1_cf_w_0_140_s_0_210=9.25e-12
+  mcm3m2p1_ca_w_0_140_s_0_280=8.53e-05 mcm3m2p1_cc_w_0_140_s_0_280=6.96e-11 mcm3m2p1_cf_w_0_140_s_0_280=1.18e-11
+  mcm3m2p1_ca_w_0_140_s_0_350=8.53e-05 mcm3m2p1_cc_w_0_140_s_0_350=5.94e-11 mcm3m2p1_cf_w_0_140_s_0_350=1.44e-11
+  mcm3m2p1_ca_w_0_140_s_0_420=8.53e-05 mcm3m2p1_cc_w_0_140_s_0_420=5.06e-11 mcm3m2p1_cf_w_0_140_s_0_420=1.68e-11
+  mcm3m2p1_ca_w_0_140_s_0_560=8.53e-05 mcm3m2p1_cc_w_0_140_s_0_560=3.82e-11 mcm3m2p1_cf_w_0_140_s_0_560=2.12e-11
+  mcm3m2p1_ca_w_0_140_s_0_840=8.53e-05 mcm3m2p1_cc_w_0_140_s_0_840=2.37e-11 mcm3m2p1_cf_w_0_140_s_0_840=2.86e-11
+  mcm3m2p1_ca_w_0_140_s_1_540=8.53e-05 mcm3m2p1_cc_w_0_140_s_1_540=8.63e-12 mcm3m2p1_cf_w_0_140_s_1_540=3.95e-11
+  mcm3m2p1_ca_w_0_140_s_3_500=8.53e-05 mcm3m2p1_cc_w_0_140_s_3_500=7.70e-13 mcm3m2p1_cf_w_0_140_s_3_500=4.68e-11
+  mcm3m2p1_ca_w_1_120_s_0_140=8.53e-05 mcm3m2p1_cc_w_1_120_s_0_140=9.75e-11 mcm3m2p1_cf_w_1_120_s_0_140=6.58e-12
+  mcm3m2p1_ca_w_1_120_s_0_175=8.53e-05 mcm3m2p1_cc_w_1_120_s_0_175=9.44e-11 mcm3m2p1_cf_w_1_120_s_0_175=7.95e-12
+  mcm3m2p1_ca_w_1_120_s_0_210=8.53e-05 mcm3m2p1_cc_w_1_120_s_0_210=8.98e-11 mcm3m2p1_cf_w_1_120_s_0_210=9.29e-12
+  mcm3m2p1_ca_w_1_120_s_0_280=8.53e-05 mcm3m2p1_cc_w_1_120_s_0_280=7.76e-11 mcm3m2p1_cf_w_1_120_s_0_280=1.19e-11
+  mcm3m2p1_ca_w_1_120_s_0_350=8.53e-05 mcm3m2p1_cc_w_1_120_s_0_350=6.67e-11 mcm3m2p1_cf_w_1_120_s_0_350=1.45e-11
+  mcm3m2p1_ca_w_1_120_s_0_420=8.53e-05 mcm3m2p1_cc_w_1_120_s_0_420=5.68e-11 mcm3m2p1_cf_w_1_120_s_0_420=1.70e-11
+  mcm3m2p1_ca_w_1_120_s_0_560=8.53e-05 mcm3m2p1_cc_w_1_120_s_0_560=4.29e-11 mcm3m2p1_cf_w_1_120_s_0_560=2.14e-11
+  mcm3m2p1_ca_w_1_120_s_0_840=8.53e-05 mcm3m2p1_cc_w_1_120_s_0_840=2.68e-11 mcm3m2p1_cf_w_1_120_s_0_840=2.89e-11
+  mcm3m2p1_ca_w_1_120_s_1_540=8.53e-05 mcm3m2p1_cc_w_1_120_s_1_540=1.01e-11 mcm3m2p1_cf_w_1_120_s_1_540=4.07e-11
+  mcm3m2p1_ca_w_1_120_s_3_500=8.53e-05 mcm3m2p1_cc_w_1_120_s_3_500=8.95e-13 mcm3m2p1_cf_w_1_120_s_3_500=4.92e-11
+  mcm3m2l1_ca_w_0_140_s_0_140=9.58e-05 mcm3m2l1_cc_w_0_140_s_0_140=8.43e-11 mcm3m2l1_cf_w_0_140_s_0_140=7.32e-12
+  mcm3m2l1_ca_w_0_140_s_0_175=9.58e-05 mcm3m2l1_cc_w_0_140_s_0_175=8.20e-11 mcm3m2l1_cf_w_0_140_s_0_175=8.86e-12
+  mcm3m2l1_ca_w_0_140_s_0_210=9.58e-05 mcm3m2l1_cc_w_0_140_s_0_210=7.82e-11 mcm3m2l1_cf_w_0_140_s_0_210=1.04e-11
+  mcm3m2l1_ca_w_0_140_s_0_280=9.58e-05 mcm3m2l1_cc_w_0_140_s_0_280=6.79e-11 mcm3m2l1_cf_w_0_140_s_0_280=1.33e-11
+  mcm3m2l1_ca_w_0_140_s_0_350=9.58e-05 mcm3m2l1_cc_w_0_140_s_0_350=5.74e-11 mcm3m2l1_cf_w_0_140_s_0_350=1.62e-11
+  mcm3m2l1_ca_w_0_140_s_0_420=9.58e-05 mcm3m2l1_cc_w_0_140_s_0_420=4.86e-11 mcm3m2l1_cf_w_0_140_s_0_420=1.90e-11
+  mcm3m2l1_ca_w_0_140_s_0_560=9.58e-05 mcm3m2l1_cc_w_0_140_s_0_560=3.56e-11 mcm3m2l1_cf_w_0_140_s_0_560=2.38e-11
+  mcm3m2l1_ca_w_0_140_s_0_840=9.58e-05 mcm3m2l1_cc_w_0_140_s_0_840=2.10e-11 mcm3m2l1_cf_w_0_140_s_0_840=3.18e-11
+  mcm3m2l1_ca_w_0_140_s_1_540=9.58e-05 mcm3m2l1_cc_w_0_140_s_1_540=6.45e-12 mcm3m2l1_cf_w_0_140_s_1_540=4.31e-11
+  mcm3m2l1_ca_w_0_140_s_3_500=9.58e-05 mcm3m2l1_cc_w_0_140_s_3_500=3.50e-13 mcm3m2l1_cf_w_0_140_s_3_500=4.90e-11
+  mcm3m2l1_ca_w_1_120_s_0_140=9.58e-05 mcm3m2l1_cc_w_1_120_s_0_140=9.41e-11 mcm3m2l1_cf_w_1_120_s_0_140=7.37e-12
+  mcm3m2l1_ca_w_1_120_s_0_175=9.58e-05 mcm3m2l1_cc_w_1_120_s_0_175=9.06e-11 mcm3m2l1_cf_w_1_120_s_0_175=8.93e-12
+  mcm3m2l1_ca_w_1_120_s_0_210=9.58e-05 mcm3m2l1_cc_w_1_120_s_0_210=8.59e-11 mcm3m2l1_cf_w_1_120_s_0_210=1.04e-11
+  mcm3m2l1_ca_w_1_120_s_0_280=9.58e-05 mcm3m2l1_cc_w_1_120_s_0_280=7.38e-11 mcm3m2l1_cf_w_1_120_s_0_280=1.34e-11
+  mcm3m2l1_ca_w_1_120_s_0_350=9.58e-05 mcm3m2l1_cc_w_1_120_s_0_350=6.24e-11 mcm3m2l1_cf_w_1_120_s_0_350=1.63e-11
+  mcm3m2l1_ca_w_1_120_s_0_420=9.58e-05 mcm3m2l1_cc_w_1_120_s_0_420=5.28e-11 mcm3m2l1_cf_w_1_120_s_0_420=1.90e-11
+  mcm3m2l1_ca_w_1_120_s_0_560=9.58e-05 mcm3m2l1_cc_w_1_120_s_0_560=3.87e-11 mcm3m2l1_cf_w_1_120_s_0_560=2.41e-11
+  mcm3m2l1_ca_w_1_120_s_0_840=9.58e-05 mcm3m2l1_cc_w_1_120_s_0_840=2.29e-11 mcm3m2l1_cf_w_1_120_s_0_840=3.23e-11
+  mcm3m2l1_ca_w_1_120_s_1_540=9.58e-05 mcm3m2l1_cc_w_1_120_s_1_540=7.13e-12 mcm3m2l1_cf_w_1_120_s_1_540=4.42e-11
+  mcm3m2l1_ca_w_1_120_s_3_500=9.58e-05 mcm3m2l1_cc_w_1_120_s_3_500=3.80e-13 mcm3m2l1_cf_w_1_120_s_3_500=5.08e-11
+  mcm3m2m1_ca_w_0_140_s_0_140=1.55e-04 mcm3m2m1_cc_w_0_140_s_0_140=7.77e-11 mcm3m2m1_cf_w_0_140_s_0_140=1.17e-11
+  mcm3m2m1_ca_w_0_140_s_0_175=1.55e-04 mcm3m2m1_cc_w_0_140_s_0_175=7.57e-11 mcm3m2m1_cf_w_0_140_s_0_175=1.43e-11
+  mcm3m2m1_ca_w_0_140_s_0_210=1.55e-04 mcm3m2m1_cc_w_0_140_s_0_210=7.14e-11 mcm3m2m1_cf_w_0_140_s_0_210=1.68e-11
+  mcm3m2m1_ca_w_0_140_s_0_280=1.55e-04 mcm3m2m1_cc_w_0_140_s_0_280=6.00e-11 mcm3m2m1_cf_w_0_140_s_0_280=2.15e-11
+  mcm3m2m1_ca_w_0_140_s_0_350=1.55e-04 mcm3m2m1_cc_w_0_140_s_0_350=4.93e-11 mcm3m2m1_cf_w_0_140_s_0_350=2.60e-11
+  mcm3m2m1_ca_w_0_140_s_0_420=1.55e-04 mcm3m2m1_cc_w_0_140_s_0_420=3.97e-11 mcm3m2m1_cf_w_0_140_s_0_420=3.02e-11
+  mcm3m2m1_ca_w_0_140_s_0_560=1.55e-04 mcm3m2m1_cc_w_0_140_s_0_560=2.70e-11 mcm3m2m1_cf_w_0_140_s_0_560=3.73e-11
+  mcm3m2m1_ca_w_0_140_s_0_840=1.55e-04 mcm3m2m1_cc_w_0_140_s_0_840=1.29e-11 mcm3m2m1_cf_w_0_140_s_0_840=4.73e-11
+  mcm3m2m1_ca_w_0_140_s_1_540=1.55e-04 mcm3m2m1_cc_w_0_140_s_1_540=2.29e-12 mcm3m2m1_cf_w_0_140_s_1_540=5.73e-11
+  mcm3m2m1_ca_w_0_140_s_3_500=1.55e-04 mcm3m2m1_cc_w_0_140_s_3_500=7.50e-14 mcm3m2m1_cf_w_0_140_s_3_500=6.01e-11
+  mcm3m2m1_ca_w_1_120_s_0_140=1.55e-04 mcm3m2m1_cc_w_1_120_s_0_140=8.27e-11 mcm3m2m1_cf_w_1_120_s_0_140=1.17e-11
+  mcm3m2m1_ca_w_1_120_s_0_175=1.55e-04 mcm3m2m1_cc_w_1_120_s_0_175=7.97e-11 mcm3m2m1_cf_w_1_120_s_0_175=1.43e-11
+  mcm3m2m1_ca_w_1_120_s_0_210=1.55e-04 mcm3m2m1_cc_w_1_120_s_0_210=7.41e-11 mcm3m2m1_cf_w_1_120_s_0_210=1.68e-11
+  mcm3m2m1_ca_w_1_120_s_0_280=1.55e-04 mcm3m2m1_cc_w_1_120_s_0_280=6.24e-11 mcm3m2m1_cf_w_1_120_s_0_280=2.16e-11
+  mcm3m2m1_ca_w_1_120_s_0_350=1.55e-04 mcm3m2m1_cc_w_1_120_s_0_350=5.07e-11 mcm3m2m1_cf_w_1_120_s_0_350=2.60e-11
+  mcm3m2m1_ca_w_1_120_s_0_420=1.55e-04 mcm3m2m1_cc_w_1_120_s_0_420=4.15e-11 mcm3m2m1_cf_w_1_120_s_0_420=3.03e-11
+  mcm3m2m1_ca_w_1_120_s_0_560=1.55e-04 mcm3m2m1_cc_w_1_120_s_0_560=2.82e-11 mcm3m2m1_cf_w_1_120_s_0_560=3.75e-11
+  mcm3m2m1_ca_w_1_120_s_0_840=1.55e-04 mcm3m2m1_cc_w_1_120_s_0_840=1.35e-11 mcm3m2m1_cf_w_1_120_s_0_840=4.79e-11
+  mcm3m2m1_ca_w_1_120_s_1_540=1.55e-04 mcm3m2m1_cc_w_1_120_s_1_540=2.35e-12 mcm3m2m1_cf_w_1_120_s_1_540=5.82e-11
+  mcm3m2m1_ca_w_1_120_s_3_500=1.55e-04 mcm3m2m1_cc_w_1_120_s_3_500=5.00e-14 mcm3m2m1_cf_w_1_120_s_3_500=6.09e-11
+  mcm4m2f_ca_w_0_140_s_0_140=3.35e-05 mcm4m2f_cc_w_0_140_s_0_140=9.08e-11 mcm4m2f_cf_w_0_140_s_0_140=2.67e-12
+  mcm4m2f_ca_w_0_140_s_0_175=3.35e-05 mcm4m2f_cc_w_0_140_s_0_175=9.02e-11 mcm4m2f_cf_w_0_140_s_0_175=3.24e-12
+  mcm4m2f_ca_w_0_140_s_0_210=3.35e-05 mcm4m2f_cc_w_0_140_s_0_210=8.57e-11 mcm4m2f_cf_w_0_140_s_0_210=3.85e-12
+  mcm4m2f_ca_w_0_140_s_0_280=3.35e-05 mcm4m2f_cc_w_0_140_s_0_280=7.75e-11 mcm4m2f_cf_w_0_140_s_0_280=4.96e-12
+  mcm4m2f_ca_w_0_140_s_0_350=3.35e-05 mcm4m2f_cc_w_0_140_s_0_350=6.74e-11 mcm4m2f_cf_w_0_140_s_0_350=6.06e-12
+  mcm4m2f_ca_w_0_140_s_0_420=3.35e-05 mcm4m2f_cc_w_0_140_s_0_420=5.91e-11 mcm4m2f_cf_w_0_140_s_0_420=7.19e-12
+  mcm4m2f_ca_w_0_140_s_0_560=3.35e-05 mcm4m2f_cc_w_0_140_s_0_560=4.78e-11 mcm4m2f_cf_w_0_140_s_0_560=9.31e-12
+  mcm4m2f_ca_w_0_140_s_0_840=3.35e-05 mcm4m2f_cc_w_0_140_s_0_840=3.46e-11 mcm4m2f_cf_w_0_140_s_0_840=1.32e-11
+  mcm4m2f_ca_w_0_140_s_1_540=3.35e-05 mcm4m2f_cc_w_0_140_s_1_540=1.83e-11 mcm4m2f_cf_w_0_140_s_1_540=2.11e-11
+  mcm4m2f_ca_w_0_140_s_3_500=3.35e-05 mcm4m2f_cc_w_0_140_s_3_500=4.27e-12 mcm4m2f_cf_w_0_140_s_3_500=3.16e-11
+  mcm4m2f_ca_w_1_120_s_0_140=3.35e-05 mcm4m2f_cc_w_1_120_s_0_140=1.13e-10 mcm4m2f_cf_w_1_120_s_0_140=2.69e-12
+  mcm4m2f_ca_w_1_120_s_0_175=3.35e-05 mcm4m2f_cc_w_1_120_s_0_175=1.09e-10 mcm4m2f_cf_w_1_120_s_0_175=3.27e-12
+  mcm4m2f_ca_w_1_120_s_0_210=3.35e-05 mcm4m2f_cc_w_1_120_s_0_210=1.05e-10 mcm4m2f_cf_w_1_120_s_0_210=3.84e-12
+  mcm4m2f_ca_w_1_120_s_0_280=3.35e-05 mcm4m2f_cc_w_1_120_s_0_280=9.29e-11 mcm4m2f_cf_w_1_120_s_0_280=4.98e-12
+  mcm4m2f_ca_w_1_120_s_0_350=3.35e-05 mcm4m2f_cc_w_1_120_s_0_350=8.17e-11 mcm4m2f_cf_w_1_120_s_0_350=6.10e-12
+  mcm4m2f_ca_w_1_120_s_0_420=3.35e-05 mcm4m2f_cc_w_1_120_s_0_420=7.18e-11 mcm4m2f_cf_w_1_120_s_0_420=7.21e-12
+  mcm4m2f_ca_w_1_120_s_0_560=3.35e-05 mcm4m2f_cc_w_1_120_s_0_560=5.83e-11 mcm4m2f_cf_w_1_120_s_0_560=9.35e-12
+  mcm4m2f_ca_w_1_120_s_0_840=3.35e-05 mcm4m2f_cc_w_1_120_s_0_840=4.17e-11 mcm4m2f_cf_w_1_120_s_0_840=1.34e-11
+  mcm4m2f_ca_w_1_120_s_1_540=3.35e-05 mcm4m2f_cc_w_1_120_s_1_540=2.23e-11 mcm4m2f_cf_w_1_120_s_1_540=2.18e-11
+  mcm4m2f_ca_w_1_120_s_3_500=3.35e-05 mcm4m2f_cc_w_1_120_s_3_500=5.36e-12 mcm4m2f_cf_w_1_120_s_3_500=3.40e-11
+  mcm4m2d_ca_w_0_140_s_0_140=3.65e-05 mcm4m2d_cc_w_0_140_s_0_140=9.04e-11 mcm4m2d_cf_w_0_140_s_0_140=2.91e-12
+  mcm4m2d_ca_w_0_140_s_0_175=3.65e-05 mcm4m2d_cc_w_0_140_s_0_175=8.98e-11 mcm4m2d_cf_w_0_140_s_0_175=3.53e-12
+  mcm4m2d_ca_w_0_140_s_0_210=3.65e-05 mcm4m2d_cc_w_0_140_s_0_210=8.53e-11 mcm4m2d_cf_w_0_140_s_0_210=4.19e-12
+  mcm4m2d_ca_w_0_140_s_0_280=3.65e-05 mcm4m2d_cc_w_0_140_s_0_280=7.70e-11 mcm4m2d_cf_w_0_140_s_0_280=5.40e-12
+  mcm4m2d_ca_w_0_140_s_0_350=3.65e-05 mcm4m2d_cc_w_0_140_s_0_350=6.68e-11 mcm4m2d_cf_w_0_140_s_0_350=6.60e-12
+  mcm4m2d_ca_w_0_140_s_0_420=3.65e-05 mcm4m2d_cc_w_0_140_s_0_420=5.89e-11 mcm4m2d_cf_w_0_140_s_0_420=7.86e-12
+  mcm4m2d_ca_w_0_140_s_0_560=3.65e-05 mcm4m2d_cc_w_0_140_s_0_560=4.74e-11 mcm4m2d_cf_w_0_140_s_0_560=1.01e-11
+  mcm4m2d_ca_w_0_140_s_0_840=3.65e-05 mcm4m2d_cc_w_0_140_s_0_840=3.35e-11 mcm4m2d_cf_w_0_140_s_0_840=1.43e-11
+  mcm4m2d_ca_w_0_140_s_1_540=3.65e-05 mcm4m2d_cc_w_0_140_s_1_540=1.72e-11 mcm4m2d_cf_w_0_140_s_1_540=2.26e-11
+  mcm4m2d_ca_w_0_140_s_3_500=3.65e-05 mcm4m2d_cc_w_0_140_s_3_500=3.59e-12 mcm4m2d_cf_w_0_140_s_3_500=3.31e-11
+  mcm4m2d_ca_w_1_120_s_0_140=3.65e-05 mcm4m2d_cc_w_1_120_s_0_140=1.11e-10 mcm4m2d_cf_w_1_120_s_0_140=2.94e-12
+  mcm4m2d_ca_w_1_120_s_0_175=3.65e-05 mcm4m2d_cc_w_1_120_s_0_175=1.08e-10 mcm4m2d_cf_w_1_120_s_0_175=3.56e-12
+  mcm4m2d_ca_w_1_120_s_0_210=3.65e-05 mcm4m2d_cc_w_1_120_s_0_210=1.03e-10 mcm4m2d_cf_w_1_120_s_0_210=4.19e-12
+  mcm4m2d_ca_w_1_120_s_0_280=3.65e-05 mcm4m2d_cc_w_1_120_s_0_280=9.15e-11 mcm4m2d_cf_w_1_120_s_0_280=5.43e-12
+  mcm4m2d_ca_w_1_120_s_0_350=3.65e-05 mcm4m2d_cc_w_1_120_s_0_350=8.02e-11 mcm4m2d_cf_w_1_120_s_0_350=6.65e-12
+  mcm4m2d_ca_w_1_120_s_0_420=3.65e-05 mcm4m2d_cc_w_1_120_s_0_420=7.06e-11 mcm4m2d_cf_w_1_120_s_0_420=7.89e-12
+  mcm4m2d_ca_w_1_120_s_0_560=3.65e-05 mcm4m2d_cc_w_1_120_s_0_560=5.67e-11 mcm4m2d_cf_w_1_120_s_0_560=1.02e-11
+  mcm4m2d_ca_w_1_120_s_0_840=3.65e-05 mcm4m2d_cc_w_1_120_s_0_840=4.00e-11 mcm4m2d_cf_w_1_120_s_0_840=1.45e-11
+  mcm4m2d_ca_w_1_120_s_1_540=3.65e-05 mcm4m2d_cc_w_1_120_s_1_540=2.08e-11 mcm4m2d_cf_w_1_120_s_1_540=2.34e-11
+  mcm4m2d_ca_w_1_120_s_3_500=3.65e-05 mcm4m2d_cc_w_1_120_s_3_500=4.48e-12 mcm4m2d_cf_w_1_120_s_3_500=3.55e-11
+  mcm4m2p1_ca_w_0_140_s_0_140=3.90e-05 mcm4m2p1_cc_w_0_140_s_0_140=9.01e-11 mcm4m2p1_cf_w_0_140_s_0_140=3.11e-12
+  mcm4m2p1_ca_w_0_140_s_0_175=3.90e-05 mcm4m2p1_cc_w_0_140_s_0_175=8.96e-11 mcm4m2p1_cf_w_0_140_s_0_175=3.77e-12
+  mcm4m2p1_ca_w_0_140_s_0_210=3.90e-05 mcm4m2p1_cc_w_0_140_s_0_210=8.50e-11 mcm4m2p1_cf_w_0_140_s_0_210=4.47e-12
+  mcm4m2p1_ca_w_0_140_s_0_280=3.90e-05 mcm4m2p1_cc_w_0_140_s_0_280=7.65e-11 mcm4m2p1_cf_w_0_140_s_0_280=5.77e-12
+  mcm4m2p1_ca_w_0_140_s_0_350=3.90e-05 mcm4m2p1_cc_w_0_140_s_0_350=6.63e-11 mcm4m2p1_cf_w_0_140_s_0_350=7.06e-12
+  mcm4m2p1_ca_w_0_140_s_0_420=3.90e-05 mcm4m2p1_cc_w_0_140_s_0_420=5.83e-11 mcm4m2p1_cf_w_0_140_s_0_420=8.37e-12
+  mcm4m2p1_ca_w_0_140_s_0_560=3.90e-05 mcm4m2p1_cc_w_0_140_s_0_560=4.68e-11 mcm4m2p1_cf_w_0_140_s_0_560=1.08e-11
+  mcm4m2p1_ca_w_0_140_s_0_840=3.90e-05 mcm4m2p1_cc_w_0_140_s_0_840=3.27e-11 mcm4m2p1_cf_w_0_140_s_0_840=1.52e-11
+  mcm4m2p1_ca_w_0_140_s_1_540=3.90e-05 mcm4m2p1_cc_w_0_140_s_1_540=1.63e-11 mcm4m2p1_cf_w_0_140_s_1_540=2.38e-11
+  mcm4m2p1_ca_w_0_140_s_3_500=3.90e-05 mcm4m2p1_cc_w_0_140_s_3_500=3.14e-12 mcm4m2p1_cf_w_0_140_s_3_500=3.44e-11
+  mcm4m2p1_ca_w_1_120_s_0_140=3.90e-05 mcm4m2p1_cc_w_1_120_s_0_140=1.10e-10 mcm4m2p1_cf_w_1_120_s_0_140=3.16e-12
+  mcm4m2p1_ca_w_1_120_s_0_175=3.90e-05 mcm4m2p1_cc_w_1_120_s_0_175=1.07e-10 mcm4m2p1_cf_w_1_120_s_0_175=3.84e-12
+  mcm4m2p1_ca_w_1_120_s_0_210=3.90e-05 mcm4m2p1_cc_w_1_120_s_0_210=1.02e-10 mcm4m2p1_cf_w_1_120_s_0_210=4.50e-12
+  mcm4m2p1_ca_w_1_120_s_0_280=3.90e-05 mcm4m2p1_cc_w_1_120_s_0_280=9.03e-11 mcm4m2p1_cf_w_1_120_s_0_280=5.82e-12
+  mcm4m2p1_ca_w_1_120_s_0_350=3.90e-05 mcm4m2p1_cc_w_1_120_s_0_350=7.91e-11 mcm4m2p1_cf_w_1_120_s_0_350=7.13e-12
+  mcm4m2p1_ca_w_1_120_s_0_420=3.90e-05 mcm4m2p1_cc_w_1_120_s_0_420=6.94e-11 mcm4m2p1_cf_w_1_120_s_0_420=8.41e-12
+  mcm4m2p1_ca_w_1_120_s_0_560=3.90e-05 mcm4m2p1_cc_w_1_120_s_0_560=5.54e-11 mcm4m2p1_cf_w_1_120_s_0_560=1.09e-11
+  mcm4m2p1_ca_w_1_120_s_0_840=3.90e-05 mcm4m2p1_cc_w_1_120_s_0_840=3.88e-11 mcm4m2p1_cf_w_1_120_s_0_840=1.55e-11
+  mcm4m2p1_ca_w_1_120_s_1_540=3.90e-05 mcm4m2p1_cc_w_1_120_s_1_540=1.96e-11 mcm4m2p1_cf_w_1_120_s_1_540=2.47e-11
+  mcm4m2p1_ca_w_1_120_s_3_500=3.90e-05 mcm4m2p1_cc_w_1_120_s_3_500=3.86e-12 mcm4m2p1_cf_w_1_120_s_3_500=3.67e-11
+  mcm4m2l1_ca_w_0_140_s_0_140=4.95e-05 mcm4m2l1_cc_w_0_140_s_0_140=8.89e-11 mcm4m2l1_cf_w_0_140_s_0_140=3.93e-12
+  mcm4m2l1_ca_w_0_140_s_0_175=4.95e-05 mcm4m2l1_cc_w_0_140_s_0_175=8.83e-11 mcm4m2l1_cf_w_0_140_s_0_175=4.77e-12
+  mcm4m2l1_ca_w_0_140_s_0_210=4.95e-05 mcm4m2l1_cc_w_0_140_s_0_210=8.35e-11 mcm4m2l1_cf_w_0_140_s_0_210=5.65e-12
+  mcm4m2l1_ca_w_0_140_s_0_280=4.95e-05 mcm4m2l1_cc_w_0_140_s_0_280=7.48e-11 mcm4m2l1_cf_w_0_140_s_0_280=7.29e-12
+  mcm4m2l1_ca_w_0_140_s_0_350=4.95e-05 mcm4m2l1_cc_w_0_140_s_0_350=6.46e-11 mcm4m2l1_cf_w_0_140_s_0_350=8.91e-12
+  mcm4m2l1_ca_w_0_140_s_0_420=4.95e-05 mcm4m2l1_cc_w_0_140_s_0_420=5.59e-11 mcm4m2l1_cf_w_0_140_s_0_420=1.05e-11
+  mcm4m2l1_ca_w_0_140_s_0_560=4.95e-05 mcm4m2l1_cc_w_0_140_s_0_560=4.41e-11 mcm4m2l1_cf_w_0_140_s_0_560=1.35e-11
+  mcm4m2l1_ca_w_0_140_s_0_840=4.95e-05 mcm4m2l1_cc_w_0_140_s_0_840=2.98e-11 mcm4m2l1_cf_w_0_140_s_0_840=1.89e-11
+  mcm4m2l1_ca_w_0_140_s_1_540=4.95e-05 mcm4m2l1_cc_w_0_140_s_1_540=1.35e-11 mcm4m2l1_cf_w_0_140_s_1_540=2.86e-11
+  mcm4m2l1_ca_w_0_140_s_3_500=4.95e-05 mcm4m2l1_cc_w_0_140_s_3_500=1.95e-12 mcm4m2l1_cf_w_0_140_s_3_500=3.84e-11
+  mcm4m2l1_ca_w_1_120_s_0_140=4.95e-05 mcm4m2l1_cc_w_1_120_s_0_140=1.06e-10 mcm4m2l1_cf_w_1_120_s_0_140=3.95e-12
+  mcm4m2l1_ca_w_1_120_s_0_175=4.95e-05 mcm4m2l1_cc_w_1_120_s_0_175=1.02e-10 mcm4m2l1_cf_w_1_120_s_0_175=4.80e-12
+  mcm4m2l1_ca_w_1_120_s_0_210=4.95e-05 mcm4m2l1_cc_w_1_120_s_0_210=9.84e-11 mcm4m2l1_cf_w_1_120_s_0_210=5.65e-12
+  mcm4m2l1_ca_w_1_120_s_0_280=4.95e-05 mcm4m2l1_cc_w_1_120_s_0_280=8.64e-11 mcm4m2l1_cf_w_1_120_s_0_280=7.32e-12
+  mcm4m2l1_ca_w_1_120_s_0_350=4.95e-05 mcm4m2l1_cc_w_1_120_s_0_350=7.48e-11 mcm4m2l1_cf_w_1_120_s_0_350=8.95e-12
+  mcm4m2l1_ca_w_1_120_s_0_420=4.95e-05 mcm4m2l1_cc_w_1_120_s_0_420=6.54e-11 mcm4m2l1_cf_w_1_120_s_0_420=1.06e-11
+  mcm4m2l1_ca_w_1_120_s_0_560=4.95e-05 mcm4m2l1_cc_w_1_120_s_0_560=5.13e-11 mcm4m2l1_cf_w_1_120_s_0_560=1.36e-11
+  mcm4m2l1_ca_w_1_120_s_0_840=4.95e-05 mcm4m2l1_cc_w_1_120_s_0_840=3.47e-11 mcm4m2l1_cf_w_1_120_s_0_840=1.92e-11
+  mcm4m2l1_ca_w_1_120_s_1_540=4.95e-05 mcm4m2l1_cc_w_1_120_s_1_540=1.59e-11 mcm4m2l1_cf_w_1_120_s_1_540=2.96e-11
+  mcm4m2l1_ca_w_1_120_s_3_500=4.95e-05 mcm4m2l1_cc_w_1_120_s_3_500=2.39e-12 mcm4m2l1_cf_w_1_120_s_3_500=4.09e-11
+  mcm4m2m1_ca_w_0_140_s_0_140=1.09e-04 mcm4m2m1_cc_w_0_140_s_0_140=8.24e-11 mcm4m2m1_cf_w_0_140_s_0_140=8.30e-12
+  mcm4m2m1_ca_w_0_140_s_0_175=1.09e-04 mcm4m2m1_cc_w_0_140_s_0_175=8.07e-11 mcm4m2m1_cf_w_0_140_s_0_175=1.02e-11
+  mcm4m2m1_ca_w_0_140_s_0_210=1.09e-04 mcm4m2m1_cc_w_0_140_s_0_210=7.70e-11 mcm4m2m1_cf_w_0_140_s_0_210=1.20e-11
+  mcm4m2m1_ca_w_0_140_s_0_280=1.09e-04 mcm4m2m1_cc_w_0_140_s_0_280=6.69e-11 mcm4m2m1_cf_w_0_140_s_0_280=1.55e-11
+  mcm4m2m1_ca_w_0_140_s_0_350=1.09e-04 mcm4m2m1_cc_w_0_140_s_0_350=5.62e-11 mcm4m2m1_cf_w_0_140_s_0_350=1.87e-11
+  mcm4m2m1_ca_w_0_140_s_0_420=1.09e-04 mcm4m2m1_cc_w_0_140_s_0_420=4.75e-11 mcm4m2m1_cf_w_0_140_s_0_420=2.18e-11
+  mcm4m2m1_ca_w_0_140_s_0_560=1.09e-04 mcm4m2m1_cc_w_0_140_s_0_560=3.51e-11 mcm4m2m1_cf_w_0_140_s_0_560=2.74e-11
+  mcm4m2m1_ca_w_0_140_s_0_840=1.09e-04 mcm4m2m1_cc_w_0_140_s_0_840=2.08e-11 mcm4m2m1_cf_w_0_140_s_0_840=3.57e-11
+  mcm4m2m1_ca_w_0_140_s_1_540=1.09e-04 mcm4m2m1_cc_w_0_140_s_1_540=7.01e-12 mcm4m2m1_cf_w_0_140_s_1_540=4.70e-11
+  mcm4m2m1_ca_w_0_140_s_3_500=1.09e-04 mcm4m2m1_cc_w_0_140_s_3_500=6.00e-13 mcm4m2m1_cf_w_0_140_s_3_500=5.34e-11
+  mcm4m2m1_ca_w_1_120_s_0_140=1.09e-04 mcm4m2m1_cc_w_1_120_s_0_140=9.48e-11 mcm4m2m1_cf_w_1_120_s_0_140=8.31e-12
+  mcm4m2m1_ca_w_1_120_s_0_175=1.09e-04 mcm4m2m1_cc_w_1_120_s_0_175=9.13e-11 mcm4m2m1_cf_w_1_120_s_0_175=1.02e-11
+  mcm4m2m1_ca_w_1_120_s_0_210=1.09e-04 mcm4m2m1_cc_w_1_120_s_0_210=8.67e-11 mcm4m2m1_cf_w_1_120_s_0_210=1.20e-11
+  mcm4m2m1_ca_w_1_120_s_0_280=1.09e-04 mcm4m2m1_cc_w_1_120_s_0_280=7.47e-11 mcm4m2m1_cf_w_1_120_s_0_280=1.55e-11
+  mcm4m2m1_ca_w_1_120_s_0_350=1.09e-04 mcm4m2m1_cc_w_1_120_s_0_350=6.33e-11 mcm4m2m1_cf_w_1_120_s_0_350=1.88e-11
+  mcm4m2m1_ca_w_1_120_s_0_420=1.09e-04 mcm4m2m1_cc_w_1_120_s_0_420=5.39e-11 mcm4m2m1_cf_w_1_120_s_0_420=2.19e-11
+  mcm4m2m1_ca_w_1_120_s_0_560=1.09e-04 mcm4m2m1_cc_w_1_120_s_0_560=4.01e-11 mcm4m2m1_cf_w_1_120_s_0_560=2.74e-11
+  mcm4m2m1_ca_w_1_120_s_0_840=1.09e-04 mcm4m2m1_cc_w_1_120_s_0_840=2.45e-11 mcm4m2m1_cf_w_1_120_s_0_840=3.61e-11
+  mcm4m2m1_ca_w_1_120_s_1_540=1.09e-04 mcm4m2m1_cc_w_1_120_s_1_540=8.82e-12 mcm4m2m1_cf_w_1_120_s_1_540=4.84e-11
+  mcm4m2m1_ca_w_1_120_s_3_500=1.09e-04 mcm4m2m1_cc_w_1_120_s_3_500=7.55e-13 mcm4m2m1_cf_w_1_120_s_3_500=5.62e-11
+  mcm5m2f_ca_w_0_140_s_0_140=2.54e-05 mcm5m2f_cc_w_0_140_s_0_140=9.19e-11 mcm5m2f_cf_w_0_140_s_0_140=2.04e-12
+  mcm5m2f_ca_w_0_140_s_0_175=2.54e-05 mcm5m2f_cc_w_0_140_s_0_175=9.15e-11 mcm5m2f_cf_w_0_140_s_0_175=2.47e-12
+  mcm5m2f_ca_w_0_140_s_0_210=2.54e-05 mcm5m2f_cc_w_0_140_s_0_210=8.70e-11 mcm5m2f_cf_w_0_140_s_0_210=2.93e-12
+  mcm5m2f_ca_w_0_140_s_0_280=2.54e-05 mcm5m2f_cc_w_0_140_s_0_280=7.85e-11 mcm5m2f_cf_w_0_140_s_0_280=3.80e-12
+  mcm5m2f_ca_w_0_140_s_0_350=2.54e-05 mcm5m2f_cc_w_0_140_s_0_350=6.91e-11 mcm5m2f_cf_w_0_140_s_0_350=4.64e-12
+  mcm5m2f_ca_w_0_140_s_0_420=2.54e-05 mcm5m2f_cc_w_0_140_s_0_420=6.12e-11 mcm5m2f_cf_w_0_140_s_0_420=5.54e-12
+  mcm5m2f_ca_w_0_140_s_0_560=2.54e-05 mcm5m2f_cc_w_0_140_s_0_560=5.02e-11 mcm5m2f_cf_w_0_140_s_0_560=7.18e-12
+  mcm5m2f_ca_w_0_140_s_0_840=2.54e-05 mcm5m2f_cc_w_0_140_s_0_840=3.73e-11 mcm5m2f_cf_w_0_140_s_0_840=1.03e-11
+  mcm5m2f_ca_w_0_140_s_1_540=2.54e-05 mcm5m2f_cc_w_0_140_s_1_540=2.16e-11 mcm5m2f_cf_w_0_140_s_1_540=1.68e-11
+  mcm5m2f_ca_w_0_140_s_3_500=2.54e-05 mcm5m2f_cc_w_0_140_s_3_500=6.62e-12 mcm5m2f_cf_w_0_140_s_3_500=2.72e-11
+  mcm5m2f_ca_w_1_120_s_0_140=2.54e-05 mcm5m2f_cc_w_1_120_s_0_140=1.16e-10 mcm5m2f_cf_w_1_120_s_0_140=2.05e-12
+  mcm5m2f_ca_w_1_120_s_0_175=2.54e-05 mcm5m2f_cc_w_1_120_s_0_175=1.12e-10 mcm5m2f_cf_w_1_120_s_0_175=2.50e-12
+  mcm5m2f_ca_w_1_120_s_0_210=2.54e-05 mcm5m2f_cc_w_1_120_s_0_210=1.09e-10 mcm5m2f_cf_w_1_120_s_0_210=2.94e-12
+  mcm5m2f_ca_w_1_120_s_0_280=2.54e-05 mcm5m2f_cc_w_1_120_s_0_280=9.68e-11 mcm5m2f_cf_w_1_120_s_0_280=3.81e-12
+  mcm5m2f_ca_w_1_120_s_0_350=2.54e-05 mcm5m2f_cc_w_1_120_s_0_350=8.54e-11 mcm5m2f_cf_w_1_120_s_0_350=4.67e-12
+  mcm5m2f_ca_w_1_120_s_0_420=2.54e-05 mcm5m2f_cc_w_1_120_s_0_420=7.61e-11 mcm5m2f_cf_w_1_120_s_0_420=5.53e-12
+  mcm5m2f_ca_w_1_120_s_0_560=2.54e-05 mcm5m2f_cc_w_1_120_s_0_560=6.26e-11 mcm5m2f_cf_w_1_120_s_0_560=7.20e-12
+  mcm5m2f_ca_w_1_120_s_0_840=2.54e-05 mcm5m2f_cc_w_1_120_s_0_840=4.63e-11 mcm5m2f_cf_w_1_120_s_0_840=1.04e-11
+  mcm5m2f_ca_w_1_120_s_1_540=2.54e-05 mcm5m2f_cc_w_1_120_s_1_540=2.71e-11 mcm5m2f_cf_w_1_120_s_1_540=1.73e-11
+  mcm5m2f_ca_w_1_120_s_3_500=2.54e-05 mcm5m2f_cc_w_1_120_s_3_500=8.59e-12 mcm5m2f_cf_w_1_120_s_3_500=2.92e-11
+  mcm5m2d_ca_w_0_140_s_0_140=2.84e-05 mcm5m2d_cc_w_0_140_s_0_140=9.15e-11 mcm5m2d_cf_w_0_140_s_0_140=2.27e-12
+  mcm5m2d_ca_w_0_140_s_0_175=2.84e-05 mcm5m2d_cc_w_0_140_s_0_175=9.11e-11 mcm5m2d_cf_w_0_140_s_0_175=2.76e-12
+  mcm5m2d_ca_w_0_140_s_0_210=2.84e-05 mcm5m2d_cc_w_0_140_s_0_210=8.65e-11 mcm5m2d_cf_w_0_140_s_0_210=3.27e-12
+  mcm5m2d_ca_w_0_140_s_0_280=2.84e-05 mcm5m2d_cc_w_0_140_s_0_280=7.81e-11 mcm5m2d_cf_w_0_140_s_0_280=4.24e-12
+  mcm5m2d_ca_w_0_140_s_0_350=2.84e-05 mcm5m2d_cc_w_0_140_s_0_350=6.85e-11 mcm5m2d_cf_w_0_140_s_0_350=5.18e-12
+  mcm5m2d_ca_w_0_140_s_0_420=2.84e-05 mcm5m2d_cc_w_0_140_s_0_420=6.05e-11 mcm5m2d_cf_w_0_140_s_0_420=6.18e-12
+  mcm5m2d_ca_w_0_140_s_0_560=2.84e-05 mcm5m2d_cc_w_0_140_s_0_560=4.94e-11 mcm5m2d_cf_w_0_140_s_0_560=7.99e-12
+  mcm5m2d_ca_w_0_140_s_0_840=2.84e-05 mcm5m2d_cc_w_0_140_s_0_840=3.63e-11 mcm5m2d_cf_w_0_140_s_0_840=1.14e-11
+  mcm5m2d_ca_w_0_140_s_1_540=2.84e-05 mcm5m2d_cc_w_0_140_s_1_540=2.04e-11 mcm5m2d_cf_w_0_140_s_1_540=1.85e-11
+  mcm5m2d_ca_w_0_140_s_3_500=2.84e-05 mcm5m2d_cc_w_0_140_s_3_500=5.74e-12 mcm5m2d_cf_w_0_140_s_3_500=2.90e-11
+  mcm5m2d_ca_w_1_120_s_0_140=2.84e-05 mcm5m2d_cc_w_1_120_s_0_140=1.15e-10 mcm5m2d_cf_w_1_120_s_0_140=2.30e-12
+  mcm5m2d_ca_w_1_120_s_0_175=2.84e-05 mcm5m2d_cc_w_1_120_s_0_175=1.11e-10 mcm5m2d_cf_w_1_120_s_0_175=2.79e-12
+  mcm5m2d_ca_w_1_120_s_0_210=2.84e-05 mcm5m2d_cc_w_1_120_s_0_210=1.07e-10 mcm5m2d_cf_w_1_120_s_0_210=3.28e-12
+  mcm5m2d_ca_w_1_120_s_0_280=2.84e-05 mcm5m2d_cc_w_1_120_s_0_280=9.54e-11 mcm5m2d_cf_w_1_120_s_0_280=4.26e-12
+  mcm5m2d_ca_w_1_120_s_0_350=2.84e-05 mcm5m2d_cc_w_1_120_s_0_350=8.42e-11 mcm5m2d_cf_w_1_120_s_0_350=5.23e-12
+  mcm5m2d_ca_w_1_120_s_0_420=2.84e-05 mcm5m2d_cc_w_1_120_s_0_420=7.45e-11 mcm5m2d_cf_w_1_120_s_0_420=6.17e-12
+  mcm5m2d_ca_w_1_120_s_0_560=2.84e-05 mcm5m2d_cc_w_1_120_s_0_560=6.11e-11 mcm5m2d_cf_w_1_120_s_0_560=8.02e-12
+  mcm5m2d_ca_w_1_120_s_0_840=2.84e-05 mcm5m2d_cc_w_1_120_s_0_840=4.47e-11 mcm5m2d_cf_w_1_120_s_0_840=1.15e-11
+  mcm5m2d_ca_w_1_120_s_1_540=2.84e-05 mcm5m2d_cc_w_1_120_s_1_540=2.54e-11 mcm5m2d_cf_w_1_120_s_1_540=1.90e-11
+  mcm5m2d_ca_w_1_120_s_3_500=2.84e-05 mcm5m2d_cc_w_1_120_s_3_500=7.44e-12 mcm5m2d_cf_w_1_120_s_3_500=3.11e-11
+  mcm5m2p1_ca_w_0_140_s_0_140=3.09e-05 mcm5m2p1_cc_w_0_140_s_0_140=9.12e-11 mcm5m2p1_cf_w_0_140_s_0_140=2.48e-12
+  mcm5m2p1_ca_w_0_140_s_0_175=3.09e-05 mcm5m2p1_cc_w_0_140_s_0_175=9.07e-11 mcm5m2p1_cf_w_0_140_s_0_175=3.01e-12
+  mcm5m2p1_ca_w_0_140_s_0_210=3.09e-05 mcm5m2p1_cc_w_0_140_s_0_210=8.62e-11 mcm5m2p1_cf_w_0_140_s_0_210=3.57e-12
+  mcm5m2p1_ca_w_0_140_s_0_280=3.09e-05 mcm5m2p1_cc_w_0_140_s_0_280=7.76e-11 mcm5m2p1_cf_w_0_140_s_0_280=4.62e-12
+  mcm5m2p1_ca_w_0_140_s_0_350=3.09e-05 mcm5m2p1_cc_w_0_140_s_0_350=6.82e-11 mcm5m2p1_cf_w_0_140_s_0_350=5.64e-12
+  mcm5m2p1_ca_w_0_140_s_0_420=3.09e-05 mcm5m2p1_cc_w_0_140_s_0_420=6.00e-11 mcm5m2p1_cf_w_0_140_s_0_420=6.72e-12
+  mcm5m2p1_ca_w_0_140_s_0_560=3.09e-05 mcm5m2p1_cc_w_0_140_s_0_560=4.87e-11 mcm5m2p1_cf_w_0_140_s_0_560=8.68e-12
+  mcm5m2p1_ca_w_0_140_s_0_840=3.09e-05 mcm5m2p1_cc_w_0_140_s_0_840=3.54e-11 mcm5m2p1_cf_w_0_140_s_0_840=1.23e-11
+  mcm5m2p1_ca_w_0_140_s_1_540=3.09e-05 mcm5m2p1_cc_w_0_140_s_1_540=1.94e-11 mcm5m2p1_cf_w_0_140_s_1_540=1.98e-11
+  mcm5m2p1_ca_w_0_140_s_3_500=3.09e-05 mcm5m2p1_cc_w_0_140_s_3_500=5.12e-12 mcm5m2p1_cf_w_0_140_s_3_500=3.04e-11
+  mcm5m2p1_ca_w_1_120_s_0_140=3.09e-05 mcm5m2p1_cc_w_1_120_s_0_140=1.14e-10 mcm5m2p1_cf_w_1_120_s_0_140=2.52e-12
+  mcm5m2p1_ca_w_1_120_s_0_175=3.09e-05 mcm5m2p1_cc_w_1_120_s_0_175=1.10e-10 mcm5m2p1_cf_w_1_120_s_0_175=3.07e-12
+  mcm5m2p1_ca_w_1_120_s_0_210=3.09e-05 mcm5m2p1_cc_w_1_120_s_0_210=1.06e-10 mcm5m2p1_cf_w_1_120_s_0_210=3.59e-12
+  mcm5m2p1_ca_w_1_120_s_0_280=3.09e-05 mcm5m2p1_cc_w_1_120_s_0_280=9.43e-11 mcm5m2p1_cf_w_1_120_s_0_280=4.66e-12
+  mcm5m2p1_ca_w_1_120_s_0_350=3.09e-05 mcm5m2p1_cc_w_1_120_s_0_350=8.28e-11 mcm5m2p1_cf_w_1_120_s_0_350=5.70e-12
+  mcm5m2p1_ca_w_1_120_s_0_420=3.09e-05 mcm5m2p1_cc_w_1_120_s_0_420=7.36e-11 mcm5m2p1_cf_w_1_120_s_0_420=6.73e-12
+  mcm5m2p1_ca_w_1_120_s_0_560=3.09e-05 mcm5m2p1_cc_w_1_120_s_0_560=5.99e-11 mcm5m2p1_cf_w_1_120_s_0_560=8.73e-12
+  mcm5m2p1_ca_w_1_120_s_0_840=3.09e-05 mcm5m2p1_cc_w_1_120_s_0_840=4.33e-11 mcm5m2p1_cf_w_1_120_s_0_840=1.25e-11
+  mcm5m2p1_ca_w_1_120_s_1_540=3.09e-05 mcm5m2p1_cc_w_1_120_s_1_540=2.42e-11 mcm5m2p1_cf_w_1_120_s_1_540=2.04e-11
+  mcm5m2p1_ca_w_1_120_s_3_500=3.09e-05 mcm5m2p1_cc_w_1_120_s_3_500=6.66e-12 mcm5m2p1_cf_w_1_120_s_3_500=3.27e-11
+  mcm5m2l1_ca_w_0_140_s_0_140=4.14e-05 mcm5m2l1_cc_w_0_140_s_0_140=9.00e-11 mcm5m2l1_cf_w_0_140_s_0_140=3.29e-12
+  mcm5m2l1_ca_w_0_140_s_0_175=4.14e-05 mcm5m2l1_cc_w_0_140_s_0_175=8.94e-11 mcm5m2l1_cf_w_0_140_s_0_175=4.00e-12
+  mcm5m2l1_ca_w_0_140_s_0_210=4.14e-05 mcm5m2l1_cc_w_0_140_s_0_210=8.47e-11 mcm5m2l1_cf_w_0_140_s_0_210=4.74e-12
+  mcm5m2l1_ca_w_0_140_s_0_280=4.14e-05 mcm5m2l1_cc_w_0_140_s_0_280=7.58e-11 mcm5m2l1_cf_w_0_140_s_0_280=6.13e-12
+  mcm5m2l1_ca_w_0_140_s_0_350=4.14e-05 mcm5m2l1_cc_w_0_140_s_0_350=6.63e-11 mcm5m2l1_cf_w_0_140_s_0_350=7.49e-12
+  mcm5m2l1_ca_w_0_140_s_0_420=4.14e-05 mcm5m2l1_cc_w_0_140_s_0_420=5.76e-11 mcm5m2l1_cf_w_0_140_s_0_420=8.89e-12
+  mcm5m2l1_ca_w_0_140_s_0_560=4.14e-05 mcm5m2l1_cc_w_0_140_s_0_560=4.63e-11 mcm5m2l1_cf_w_0_140_s_0_560=1.14e-11
+  mcm5m2l1_ca_w_0_140_s_0_840=4.14e-05 mcm5m2l1_cc_w_0_140_s_0_840=3.24e-11 mcm5m2l1_cf_w_0_140_s_0_840=1.60e-11
+  mcm5m2l1_ca_w_0_140_s_1_540=4.14e-05 mcm5m2l1_cc_w_0_140_s_1_540=1.64e-11 mcm5m2l1_cf_w_0_140_s_1_540=2.49e-11
+  mcm5m2l1_ca_w_0_140_s_3_500=4.14e-05 mcm5m2l1_cc_w_0_140_s_3_500=3.49e-12 mcm5m2l1_cf_w_0_140_s_3_500=3.53e-11
+  mcm5m2l1_ca_w_1_120_s_0_140=4.14e-05 mcm5m2l1_cc_w_1_120_s_0_140=1.10e-10 mcm5m2l1_cf_w_1_120_s_0_140=3.32e-12
+  mcm5m2l1_ca_w_1_120_s_0_175=4.14e-05 mcm5m2l1_cc_w_1_120_s_0_175=1.07e-10 mcm5m2l1_cf_w_1_120_s_0_175=4.04e-12
+  mcm5m2l1_ca_w_1_120_s_0_210=4.14e-05 mcm5m2l1_cc_w_1_120_s_0_210=1.02e-10 mcm5m2l1_cf_w_1_120_s_0_210=4.74e-12
+  mcm5m2l1_ca_w_1_120_s_0_280=4.14e-05 mcm5m2l1_cc_w_1_120_s_0_280=9.04e-11 mcm5m2l1_cf_w_1_120_s_0_280=6.16e-12
+  mcm5m2l1_ca_w_1_120_s_0_350=4.14e-05 mcm5m2l1_cc_w_1_120_s_0_350=7.91e-11 mcm5m2l1_cf_w_1_120_s_0_350=7.53e-12
+  mcm5m2l1_ca_w_1_120_s_0_420=4.14e-05 mcm5m2l1_cc_w_1_120_s_0_420=6.96e-11 mcm5m2l1_cf_w_1_120_s_0_420=8.88e-12
+  mcm5m2l1_ca_w_1_120_s_0_560=4.14e-05 mcm5m2l1_cc_w_1_120_s_0_560=5.57e-11 mcm5m2l1_cf_w_1_120_s_0_560=1.15e-11
+  mcm5m2l1_ca_w_1_120_s_0_840=4.14e-05 mcm5m2l1_cc_w_1_120_s_0_840=3.93e-11 mcm5m2l1_cf_w_1_120_s_0_840=1.62e-11
+  mcm5m2l1_ca_w_1_120_s_1_540=4.14e-05 mcm5m2l1_cc_w_1_120_s_1_540=2.03e-11 mcm5m2l1_cf_w_1_120_s_1_540=2.56e-11
+  mcm5m2l1_ca_w_1_120_s_3_500=4.14e-05 mcm5m2l1_cc_w_1_120_s_3_500=4.66e-12 mcm5m2l1_cf_w_1_120_s_3_500=3.78e-11
+  mcm5m2m1_ca_w_0_140_s_0_140=1.01e-04 mcm5m2m1_cc_w_0_140_s_0_140=8.34e-11 mcm5m2m1_cf_w_0_140_s_0_140=7.66e-12
+  mcm5m2m1_ca_w_0_140_s_0_175=1.01e-04 mcm5m2m1_cc_w_0_140_s_0_175=8.18e-11 mcm5m2m1_cf_w_0_140_s_0_175=9.40e-12
+  mcm5m2m1_ca_w_0_140_s_0_210=1.01e-04 mcm5m2m1_cc_w_0_140_s_0_210=7.76e-11 mcm5m2m1_cf_w_0_140_s_0_210=1.11e-11
+  mcm5m2m1_ca_w_0_140_s_0_280=1.01e-04 mcm5m2m1_cc_w_0_140_s_0_280=6.83e-11 mcm5m2m1_cf_w_0_140_s_0_280=1.43e-11
+  mcm5m2m1_ca_w_0_140_s_0_350=1.01e-04 mcm5m2m1_cc_w_0_140_s_0_350=5.79e-11 mcm5m2m1_cf_w_0_140_s_0_350=1.73e-11
+  mcm5m2m1_ca_w_0_140_s_0_420=1.01e-04 mcm5m2m1_cc_w_0_140_s_0_420=4.92e-11 mcm5m2m1_cf_w_0_140_s_0_420=2.02e-11
+  mcm5m2m1_ca_w_0_140_s_0_560=1.01e-04 mcm5m2m1_cc_w_0_140_s_0_560=3.70e-11 mcm5m2m1_cf_w_0_140_s_0_560=2.53e-11
+  mcm5m2m1_ca_w_0_140_s_0_840=1.01e-04 mcm5m2m1_cc_w_0_140_s_0_840=2.33e-11 mcm5m2m1_cf_w_0_140_s_0_840=3.32e-11
+  mcm5m2m1_ca_w_0_140_s_1_540=1.01e-04 mcm5m2m1_cc_w_0_140_s_1_540=9.12e-12 mcm5m2m1_cf_w_0_140_s_1_540=4.44e-11
+  mcm5m2m1_ca_w_0_140_s_3_500=1.01e-04 mcm5m2m1_cc_w_0_140_s_3_500=1.30e-12 mcm5m2m1_cf_w_0_140_s_3_500=5.18e-11
+  mcm5m2m1_ca_w_1_120_s_0_140=1.01e-04 mcm5m2m1_cc_w_1_120_s_0_140=9.84e-11 mcm5m2m1_cf_w_1_120_s_0_140=7.67e-12
+  mcm5m2m1_ca_w_1_120_s_0_175=1.01e-04 mcm5m2m1_cc_w_1_120_s_0_175=9.49e-11 mcm5m2m1_cf_w_1_120_s_0_175=9.42e-12
+  mcm5m2m1_ca_w_1_120_s_0_210=1.01e-04 mcm5m2m1_cc_w_1_120_s_0_210=9.08e-11 mcm5m2m1_cf_w_1_120_s_0_210=1.11e-11
+  mcm5m2m1_ca_w_1_120_s_0_280=1.01e-04 mcm5m2m1_cc_w_1_120_s_0_280=7.86e-11 mcm5m2m1_cf_w_1_120_s_0_280=1.43e-11
+  mcm5m2m1_ca_w_1_120_s_0_350=1.01e-04 mcm5m2m1_cc_w_1_120_s_0_350=6.74e-11 mcm5m2m1_cf_w_1_120_s_0_350=1.74e-11
+  mcm5m2m1_ca_w_1_120_s_0_420=1.01e-04 mcm5m2m1_cc_w_1_120_s_0_420=5.79e-11 mcm5m2m1_cf_w_1_120_s_0_420=2.01e-11
+  mcm5m2m1_ca_w_1_120_s_0_560=1.01e-04 mcm5m2m1_cc_w_1_120_s_0_560=4.45e-11 mcm5m2m1_cf_w_1_120_s_0_560=2.53e-11
+  mcm5m2m1_ca_w_1_120_s_0_840=1.01e-04 mcm5m2m1_cc_w_1_120_s_0_840=2.89e-11 mcm5m2m1_cf_w_1_120_s_0_840=3.35e-11
+  mcm5m2m1_ca_w_1_120_s_1_540=1.01e-04 mcm5m2m1_cc_w_1_120_s_1_540=1.25e-11 mcm5m2m1_cf_w_1_120_s_1_540=4.57e-11
+  mcm5m2m1_ca_w_1_120_s_3_500=1.01e-04 mcm5m2m1_cc_w_1_120_s_3_500=2.07e-12 mcm5m2m1_cf_w_1_120_s_3_500=5.54e-11
+  mcrdlm2f_ca_w_0_140_s_0_140=1.77e-05 mcrdlm2f_cc_w_0_140_s_0_140=9.27e-11 mcrdlm2f_cf_w_0_140_s_0_140=1.42e-12
+  mcrdlm2f_ca_w_0_140_s_0_175=1.77e-05 mcrdlm2f_cc_w_0_140_s_0_175=9.13e-11 mcrdlm2f_cf_w_0_140_s_0_175=1.73e-12
+  mcrdlm2f_ca_w_0_140_s_0_210=1.77e-05 mcrdlm2f_cc_w_0_140_s_0_210=8.76e-11 mcrdlm2f_cf_w_0_140_s_0_210=2.05e-12
+  mcrdlm2f_ca_w_0_140_s_0_280=1.77e-05 mcrdlm2f_cc_w_0_140_s_0_280=7.93e-11 mcrdlm2f_cf_w_0_140_s_0_280=2.65e-12
+  mcrdlm2f_ca_w_0_140_s_0_350=1.77e-05 mcrdlm2f_cc_w_0_140_s_0_350=7.09e-11 mcrdlm2f_cf_w_0_140_s_0_350=3.25e-12
+  mcrdlm2f_ca_w_0_140_s_0_420=1.77e-05 mcrdlm2f_cc_w_0_140_s_0_420=6.24e-11 mcrdlm2f_cf_w_0_140_s_0_420=3.88e-12
+  mcrdlm2f_ca_w_0_140_s_0_560=1.77e-05 mcrdlm2f_cc_w_0_140_s_0_560=5.23e-11 mcrdlm2f_cf_w_0_140_s_0_560=5.04e-12
+  mcrdlm2f_ca_w_0_140_s_0_840=1.77e-05 mcrdlm2f_cc_w_0_140_s_0_840=4.02e-11 mcrdlm2f_cf_w_0_140_s_0_840=7.24e-12
+  mcrdlm2f_ca_w_0_140_s_1_540=1.77e-05 mcrdlm2f_cc_w_0_140_s_1_540=2.57e-11 mcrdlm2f_cf_w_0_140_s_1_540=1.22e-11
+  mcrdlm2f_ca_w_0_140_s_3_500=1.77e-05 mcrdlm2f_cc_w_0_140_s_3_500=1.11e-11 mcrdlm2f_cf_w_0_140_s_3_500=2.13e-11
+  mcrdlm2f_ca_w_1_120_s_0_140=1.77e-05 mcrdlm2f_cc_w_1_120_s_0_140=1.20e-10 mcrdlm2f_cf_w_1_120_s_0_140=1.45e-12
+  mcrdlm2f_ca_w_1_120_s_0_175=1.77e-05 mcrdlm2f_cc_w_1_120_s_0_175=1.17e-10 mcrdlm2f_cf_w_1_120_s_0_175=1.76e-12
+  mcrdlm2f_ca_w_1_120_s_0_210=1.77e-05 mcrdlm2f_cc_w_1_120_s_0_210=1.13e-10 mcrdlm2f_cf_w_1_120_s_0_210=2.06e-12
+  mcrdlm2f_ca_w_1_120_s_0_280=1.77e-05 mcrdlm2f_cc_w_1_120_s_0_280=1.01e-10 mcrdlm2f_cf_w_1_120_s_0_280=2.67e-12
+  mcrdlm2f_ca_w_1_120_s_0_350=1.77e-05 mcrdlm2f_cc_w_1_120_s_0_350=9.03e-11 mcrdlm2f_cf_w_1_120_s_0_350=3.28e-12
+  mcrdlm2f_ca_w_1_120_s_0_420=1.77e-05 mcrdlm2f_cc_w_1_120_s_0_420=8.12e-11 mcrdlm2f_cf_w_1_120_s_0_420=3.88e-12
+  mcrdlm2f_ca_w_1_120_s_0_560=1.77e-05 mcrdlm2f_cc_w_1_120_s_0_560=6.77e-11 mcrdlm2f_cf_w_1_120_s_0_560=5.05e-12
+  mcrdlm2f_ca_w_1_120_s_0_840=1.77e-05 mcrdlm2f_cc_w_1_120_s_0_840=5.22e-11 mcrdlm2f_cf_w_1_120_s_0_840=7.33e-12
+  mcrdlm2f_ca_w_1_120_s_1_540=1.77e-05 mcrdlm2f_cc_w_1_120_s_1_540=3.39e-11 mcrdlm2f_cf_w_1_120_s_1_540=1.24e-11
+  mcrdlm2f_ca_w_1_120_s_3_500=1.77e-05 mcrdlm2f_cc_w_1_120_s_3_500=1.52e-11 mcrdlm2f_cf_w_1_120_s_3_500=2.27e-11
+  mcrdlm2d_ca_w_0_140_s_0_140=2.07e-05 mcrdlm2d_cc_w_0_140_s_0_140=9.24e-11 mcrdlm2d_cf_w_0_140_s_0_140=1.66e-12
+  mcrdlm2d_ca_w_0_140_s_0_175=2.07e-05 mcrdlm2d_cc_w_0_140_s_0_175=9.11e-11 mcrdlm2d_cf_w_0_140_s_0_175=2.02e-12
+  mcrdlm2d_ca_w_0_140_s_0_210=2.07e-05 mcrdlm2d_cc_w_0_140_s_0_210=8.71e-11 mcrdlm2d_cf_w_0_140_s_0_210=2.39e-12
+  mcrdlm2d_ca_w_0_140_s_0_280=2.07e-05 mcrdlm2d_cc_w_0_140_s_0_280=7.87e-11 mcrdlm2d_cf_w_0_140_s_0_280=3.09e-12
+  mcrdlm2d_ca_w_0_140_s_0_350=2.07e-05 mcrdlm2d_cc_w_0_140_s_0_350=6.98e-11 mcrdlm2d_cf_w_0_140_s_0_350=3.78e-12
+  mcrdlm2d_ca_w_0_140_s_0_420=2.07e-05 mcrdlm2d_cc_w_0_140_s_0_420=6.22e-11 mcrdlm2d_cf_w_0_140_s_0_420=4.50e-12
+  mcrdlm2d_ca_w_0_140_s_0_560=2.07e-05 mcrdlm2d_cc_w_0_140_s_0_560=5.15e-11 mcrdlm2d_cf_w_0_140_s_0_560=5.85e-12
+  mcrdlm2d_ca_w_0_140_s_0_840=2.07e-05 mcrdlm2d_cc_w_0_140_s_0_840=3.91e-11 mcrdlm2d_cf_w_0_140_s_0_840=8.37e-12
+  mcrdlm2d_ca_w_0_140_s_1_540=2.07e-05 mcrdlm2d_cc_w_0_140_s_1_540=2.44e-11 mcrdlm2d_cf_w_0_140_s_1_540=1.39e-11
+  mcrdlm2d_ca_w_0_140_s_3_500=2.07e-05 mcrdlm2d_cc_w_0_140_s_3_500=9.83e-12 mcrdlm2d_cf_w_0_140_s_3_500=2.36e-11
+  mcrdlm2d_ca_w_1_120_s_0_140=2.07e-05 mcrdlm2d_cc_w_1_120_s_0_140=1.19e-10 mcrdlm2d_cf_w_1_120_s_0_140=1.69e-12
+  mcrdlm2d_ca_w_1_120_s_0_175=2.07e-05 mcrdlm2d_cc_w_1_120_s_0_175=1.16e-10 mcrdlm2d_cf_w_1_120_s_0_175=2.05e-12
+  mcrdlm2d_ca_w_1_120_s_0_210=2.07e-05 mcrdlm2d_cc_w_1_120_s_0_210=1.12e-10 mcrdlm2d_cf_w_1_120_s_0_210=2.41e-12
+  mcrdlm2d_ca_w_1_120_s_0_280=2.07e-05 mcrdlm2d_cc_w_1_120_s_0_280=9.99e-11 mcrdlm2d_cf_w_1_120_s_0_280=3.12e-12
+  mcrdlm2d_ca_w_1_120_s_0_350=2.07e-05 mcrdlm2d_cc_w_1_120_s_0_350=8.88e-11 mcrdlm2d_cf_w_1_120_s_0_350=3.83e-12
+  mcrdlm2d_ca_w_1_120_s_0_420=2.07e-05 mcrdlm2d_cc_w_1_120_s_0_420=7.96e-11 mcrdlm2d_cf_w_1_120_s_0_420=4.52e-12
+  mcrdlm2d_ca_w_1_120_s_0_560=2.07e-05 mcrdlm2d_cc_w_1_120_s_0_560=6.61e-11 mcrdlm2d_cf_w_1_120_s_0_560=5.88e-12
+  mcrdlm2d_ca_w_1_120_s_0_840=2.07e-05 mcrdlm2d_cc_w_1_120_s_0_840=5.05e-11 mcrdlm2d_cf_w_1_120_s_0_840=8.48e-12
+  mcrdlm2d_ca_w_1_120_s_1_540=2.07e-05 mcrdlm2d_cc_w_1_120_s_1_540=3.21e-11 mcrdlm2d_cf_w_1_120_s_1_540=1.43e-11
+  mcrdlm2d_ca_w_1_120_s_3_500=2.07e-05 mcrdlm2d_cc_w_1_120_s_3_500=1.37e-11 mcrdlm2d_cf_w_1_120_s_3_500=2.52e-11
+  mcrdlm2p1_ca_w_0_140_s_0_140=2.32e-05 mcrdlm2p1_cc_w_0_140_s_0_140=9.21e-11 mcrdlm2p1_cf_w_0_140_s_0_140=1.86e-12
+  mcrdlm2p1_ca_w_0_140_s_0_175=2.32e-05 mcrdlm2p1_cc_w_0_140_s_0_175=9.06e-11 mcrdlm2p1_cf_w_0_140_s_0_175=2.27e-12
+  mcrdlm2p1_ca_w_0_140_s_0_210=2.32e-05 mcrdlm2p1_cc_w_0_140_s_0_210=8.68e-11 mcrdlm2p1_cf_w_0_140_s_0_210=2.68e-12
+  mcrdlm2p1_ca_w_0_140_s_0_280=2.32e-05 mcrdlm2p1_cc_w_0_140_s_0_280=7.82e-11 mcrdlm2p1_cf_w_0_140_s_0_280=3.46e-12
+  mcrdlm2p1_ca_w_0_140_s_0_350=2.32e-05 mcrdlm2p1_cc_w_0_140_s_0_350=6.93e-11 mcrdlm2p1_cf_w_0_140_s_0_350=4.24e-12
+  mcrdlm2p1_ca_w_0_140_s_0_420=2.32e-05 mcrdlm2p1_cc_w_0_140_s_0_420=6.13e-11 mcrdlm2p1_cf_w_0_140_s_0_420=5.06e-12
+  mcrdlm2p1_ca_w_0_140_s_0_560=2.32e-05 mcrdlm2p1_cc_w_0_140_s_0_560=5.08e-11 mcrdlm2p1_cf_w_0_140_s_0_560=6.53e-12
+  mcrdlm2p1_ca_w_0_140_s_0_840=2.32e-05 mcrdlm2p1_cc_w_0_140_s_0_840=3.83e-11 mcrdlm2p1_cf_w_0_140_s_0_840=9.34e-12
+  mcrdlm2p1_ca_w_0_140_s_1_540=2.32e-05 mcrdlm2p1_cc_w_0_140_s_1_540=2.34e-11 mcrdlm2p1_cf_w_0_140_s_1_540=1.54e-11
+  mcrdlm2p1_ca_w_0_140_s_3_500=2.32e-05 mcrdlm2p1_cc_w_0_140_s_3_500=8.97e-12 mcrdlm2p1_cf_w_0_140_s_3_500=2.54e-11
+  mcrdlm2p1_ca_w_1_120_s_0_140=2.32e-05 mcrdlm2p1_cc_w_1_120_s_0_140=1.18e-10 mcrdlm2p1_cf_w_1_120_s_0_140=1.92e-12
+  mcrdlm2p1_ca_w_1_120_s_0_175=2.32e-05 mcrdlm2p1_cc_w_1_120_s_0_175=1.15e-10 mcrdlm2p1_cf_w_1_120_s_0_175=2.32e-12
+  mcrdlm2p1_ca_w_1_120_s_0_210=2.32e-05 mcrdlm2p1_cc_w_1_120_s_0_210=1.10e-10 mcrdlm2p1_cf_w_1_120_s_0_210=2.72e-12
+  mcrdlm2p1_ca_w_1_120_s_0_280=2.32e-05 mcrdlm2p1_cc_w_1_120_s_0_280=9.88e-11 mcrdlm2p1_cf_w_1_120_s_0_280=3.52e-12
+  mcrdlm2p1_ca_w_1_120_s_0_350=2.32e-05 mcrdlm2p1_cc_w_1_120_s_0_350=8.74e-11 mcrdlm2p1_cf_w_1_120_s_0_350=4.31e-12
+  mcrdlm2p1_ca_w_1_120_s_0_420=2.32e-05 mcrdlm2p1_cc_w_1_120_s_0_420=7.84e-11 mcrdlm2p1_cf_w_1_120_s_0_420=5.08e-12
+  mcrdlm2p1_ca_w_1_120_s_0_560=2.32e-05 mcrdlm2p1_cc_w_1_120_s_0_560=6.48e-11 mcrdlm2p1_cf_w_1_120_s_0_560=6.59e-12
+  mcrdlm2p1_ca_w_1_120_s_0_840=2.32e-05 mcrdlm2p1_cc_w_1_120_s_0_840=4.92e-11 mcrdlm2p1_cf_w_1_120_s_0_840=9.47e-12
+  mcrdlm2p1_ca_w_1_120_s_1_540=2.32e-05 mcrdlm2p1_cc_w_1_120_s_1_540=3.09e-11 mcrdlm2p1_cf_w_1_120_s_1_540=1.58e-11
+  mcrdlm2p1_ca_w_1_120_s_3_500=2.32e-05 mcrdlm2p1_cc_w_1_120_s_3_500=1.27e-11 mcrdlm2p1_cf_w_1_120_s_3_500=2.72e-11
+  mcrdlm2l1_ca_w_0_140_s_0_140=3.37e-05 mcrdlm2l1_cc_w_0_140_s_0_140=9.09e-11 mcrdlm2l1_cf_w_0_140_s_0_140=2.67e-12
+  mcrdlm2l1_ca_w_0_140_s_0_175=3.37e-05 mcrdlm2l1_cc_w_0_140_s_0_175=8.95e-11 mcrdlm2l1_cf_w_0_140_s_0_175=3.26e-12
+  mcrdlm2l1_ca_w_0_140_s_0_210=3.37e-05 mcrdlm2l1_cc_w_0_140_s_0_210=8.53e-11 mcrdlm2l1_cf_w_0_140_s_0_210=3.85e-12
+  mcrdlm2l1_ca_w_0_140_s_0_280=3.37e-05 mcrdlm2l1_cc_w_0_140_s_0_280=7.69e-11 mcrdlm2l1_cf_w_0_140_s_0_280=5.00e-12
+  mcrdlm2l1_ca_w_0_140_s_0_350=3.37e-05 mcrdlm2l1_cc_w_0_140_s_0_350=6.74e-11 mcrdlm2l1_cf_w_0_140_s_0_350=6.09e-12
+  mcrdlm2l1_ca_w_0_140_s_0_420=3.37e-05 mcrdlm2l1_cc_w_0_140_s_0_420=5.93e-11 mcrdlm2l1_cf_w_0_140_s_0_420=7.21e-12
+  mcrdlm2l1_ca_w_0_140_s_0_560=3.37e-05 mcrdlm2l1_cc_w_0_140_s_0_560=4.84e-11 mcrdlm2l1_cf_w_0_140_s_0_560=9.30e-12
+  mcrdlm2l1_ca_w_0_140_s_0_840=3.37e-05 mcrdlm2l1_cc_w_0_140_s_0_840=3.53e-11 mcrdlm2l1_cf_w_0_140_s_0_840=1.31e-11
+  mcrdlm2l1_ca_w_0_140_s_1_540=3.37e-05 mcrdlm2l1_cc_w_0_140_s_1_540=2.00e-11 mcrdlm2l1_cf_w_0_140_s_1_540=2.08e-11
+  mcrdlm2l1_ca_w_0_140_s_3_500=3.37e-05 mcrdlm2l1_cc_w_0_140_s_3_500=6.54e-12 mcrdlm2l1_cf_w_0_140_s_3_500=3.14e-11
+  mcrdlm2l1_ca_w_1_120_s_0_140=3.37e-05 mcrdlm2l1_cc_w_1_120_s_0_140=1.14e-10 mcrdlm2l1_cf_w_1_120_s_0_140=2.70e-12
+  mcrdlm2l1_ca_w_1_120_s_0_175=3.37e-05 mcrdlm2l1_cc_w_1_120_s_0_175=1.11e-10 mcrdlm2l1_cf_w_1_120_s_0_175=3.29e-12
+  mcrdlm2l1_ca_w_1_120_s_0_210=3.37e-05 mcrdlm2l1_cc_w_1_120_s_0_210=1.06e-10 mcrdlm2l1_cf_w_1_120_s_0_210=3.87e-12
+  mcrdlm2l1_ca_w_1_120_s_0_280=3.37e-05 mcrdlm2l1_cc_w_1_120_s_0_280=9.47e-11 mcrdlm2l1_cf_w_1_120_s_0_280=5.02e-12
+  mcrdlm2l1_ca_w_1_120_s_0_350=3.37e-05 mcrdlm2l1_cc_w_1_120_s_0_350=8.36e-11 mcrdlm2l1_cf_w_1_120_s_0_350=6.14e-12
+  mcrdlm2l1_ca_w_1_120_s_0_420=3.37e-05 mcrdlm2l1_cc_w_1_120_s_0_420=7.43e-11 mcrdlm2l1_cf_w_1_120_s_0_420=7.24e-12
+  mcrdlm2l1_ca_w_1_120_s_0_560=3.37e-05 mcrdlm2l1_cc_w_1_120_s_0_560=6.08e-11 mcrdlm2l1_cf_w_1_120_s_0_560=9.36e-12
+  mcrdlm2l1_ca_w_1_120_s_0_840=3.37e-05 mcrdlm2l1_cc_w_1_120_s_0_840=4.50e-11 mcrdlm2l1_cf_w_1_120_s_0_840=1.33e-11
+  mcrdlm2l1_ca_w_1_120_s_1_540=3.37e-05 mcrdlm2l1_cc_w_1_120_s_1_540=2.67e-11 mcrdlm2l1_cf_w_1_120_s_1_540=2.14e-11
+  mcrdlm2l1_ca_w_1_120_s_3_500=3.37e-05 mcrdlm2l1_cc_w_1_120_s_3_500=9.80e-12 mcrdlm2l1_cf_w_1_120_s_3_500=3.37e-11
+  mcrdlm2m1_ca_w_0_140_s_0_140=9.32e-05 mcrdlm2m1_cc_w_0_140_s_0_140=8.47e-11 mcrdlm2m1_cf_w_0_140_s_0_140=7.05e-12
+  mcrdlm2m1_ca_w_0_140_s_0_175=9.32e-05 mcrdlm2m1_cc_w_0_140_s_0_175=8.34e-11 mcrdlm2m1_cf_w_0_140_s_0_175=8.65e-12
+  mcrdlm2m1_ca_w_0_140_s_0_210=9.32e-05 mcrdlm2m1_cc_w_0_140_s_0_210=7.89e-11 mcrdlm2m1_cf_w_0_140_s_0_210=1.02e-11
+  mcrdlm2m1_ca_w_0_140_s_0_280=9.32e-05 mcrdlm2m1_cc_w_0_140_s_0_280=6.96e-11 mcrdlm2m1_cf_w_0_140_s_0_280=1.32e-11
+  mcrdlm2m1_ca_w_0_140_s_0_350=9.32e-05 mcrdlm2m1_cc_w_0_140_s_0_350=5.94e-11 mcrdlm2m1_cf_w_0_140_s_0_350=1.59e-11
+  mcrdlm2m1_ca_w_0_140_s_0_420=9.32e-05 mcrdlm2m1_cc_w_0_140_s_0_420=5.07e-11 mcrdlm2m1_cf_w_0_140_s_0_420=1.85e-11
+  mcrdlm2m1_ca_w_0_140_s_0_560=9.32e-05 mcrdlm2m1_cc_w_0_140_s_0_560=3.91e-11 mcrdlm2m1_cf_w_0_140_s_0_560=2.32e-11
+  mcrdlm2m1_ca_w_0_140_s_0_840=9.32e-05 mcrdlm2m1_cc_w_0_140_s_0_840=2.58e-11 mcrdlm2m1_cf_w_0_140_s_0_840=3.06e-11
+  mcrdlm2m1_ca_w_0_140_s_1_540=9.32e-05 mcrdlm2m1_cc_w_0_140_s_1_540=1.18e-11 mcrdlm2m1_cf_w_0_140_s_1_540=4.16e-11
+  mcrdlm2m1_ca_w_0_140_s_3_500=9.32e-05 mcrdlm2m1_cc_w_0_140_s_3_500=2.89e-12 mcrdlm2m1_cf_w_0_140_s_3_500=5.01e-11
+  mcrdlm2m1_ca_w_1_120_s_0_140=9.32e-05 mcrdlm2m1_cc_w_1_120_s_0_140=1.02e-10 mcrdlm2m1_cf_w_1_120_s_0_140=7.08e-12
+  mcrdlm2m1_ca_w_1_120_s_0_175=9.32e-05 mcrdlm2m1_cc_w_1_120_s_0_175=9.95e-11 mcrdlm2m1_cf_w_1_120_s_0_175=8.68e-12
+  mcrdlm2m1_ca_w_1_120_s_0_210=9.32e-05 mcrdlm2m1_cc_w_1_120_s_0_210=9.48e-11 mcrdlm2m1_cf_w_1_120_s_0_210=1.02e-11
+  mcrdlm2m1_ca_w_1_120_s_0_280=9.32e-05 mcrdlm2m1_cc_w_1_120_s_0_280=8.30e-11 mcrdlm2m1_cf_w_1_120_s_0_280=1.32e-11
+  mcrdlm2m1_ca_w_1_120_s_0_350=9.32e-05 mcrdlm2m1_cc_w_1_120_s_0_350=7.22e-11 mcrdlm2m1_cf_w_1_120_s_0_350=1.59e-11
+  mcrdlm2m1_ca_w_1_120_s_0_420=9.32e-05 mcrdlm2m1_cc_w_1_120_s_0_420=6.28e-11 mcrdlm2m1_cf_w_1_120_s_0_420=1.86e-11
+  mcrdlm2m1_ca_w_1_120_s_0_560=9.32e-05 mcrdlm2m1_cc_w_1_120_s_0_560=4.95e-11 mcrdlm2m1_cf_w_1_120_s_0_560=2.32e-11
+  mcrdlm2m1_ca_w_1_120_s_0_840=9.32e-05 mcrdlm2m1_cc_w_1_120_s_0_840=3.44e-11 mcrdlm2m1_cf_w_1_120_s_0_840=3.09e-11
+  mcrdlm2m1_ca_w_1_120_s_1_540=9.32e-05 mcrdlm2m1_cc_w_1_120_s_1_540=1.79e-11 mcrdlm2m1_cf_w_1_120_s_1_540=4.26e-11
+  mcrdlm2m1_ca_w_1_120_s_3_500=9.32e-05 mcrdlm2m1_cc_w_1_120_s_3_500=5.41e-12 mcrdlm2m1_cf_w_1_120_s_3_500=5.39e-11
+  mcm4m3f_ca_w_0_300_s_0_300=7.52e-05 mcm4m3f_cc_w_0_300_s_0_300=8.31e-11 mcm4m3f_cf_w_0_300_s_0_300=1.09e-11
+  mcm4m3f_ca_w_0_300_s_0_360=7.52e-05 mcm4m3f_cc_w_0_300_s_0_360=7.61e-11 mcm4m3f_cf_w_0_300_s_0_360=1.27e-11
+  mcm4m3f_ca_w_0_300_s_0_450=7.52e-05 mcm4m3f_cc_w_0_300_s_0_450=6.76e-11 mcm4m3f_cf_w_0_300_s_0_450=1.54e-11
+  mcm4m3f_ca_w_0_300_s_0_600=7.52e-05 mcm4m3f_cc_w_0_300_s_0_600=5.53e-11 mcm4m3f_cf_w_0_300_s_0_600=1.95e-11
+  mcm4m3f_ca_w_0_300_s_0_800=7.52e-05 mcm4m3f_cc_w_0_300_s_0_800=4.35e-11 mcm4m3f_cf_w_0_300_s_0_800=2.43e-11
+  mcm4m3f_ca_w_0_300_s_1_000=7.52e-05 mcm4m3f_cc_w_0_300_s_1_000=3.45e-11 mcm4m3f_cf_w_0_300_s_1_000=2.86e-11
+  mcm4m3f_ca_w_0_300_s_1_200=7.52e-05 mcm4m3f_cc_w_0_300_s_1_200=2.78e-11 mcm4m3f_cf_w_0_300_s_1_200=3.22e-11
+  mcm4m3f_ca_w_0_300_s_2_100=7.52e-05 mcm4m3f_cc_w_0_300_s_2_100=1.18e-11 mcm4m3f_cf_w_0_300_s_2_100=4.31e-11
+  mcm4m3f_ca_w_0_300_s_3_300=7.52e-05 mcm4m3f_cc_w_0_300_s_3_300=4.49e-12 mcm4m3f_cf_w_0_300_s_3_300=4.95e-11
+  mcm4m3f_ca_w_0_300_s_9_000=7.52e-05 mcm4m3f_cc_w_0_300_s_9_000=1.05e-13 mcm4m3f_cf_w_0_300_s_9_000=5.38e-11
+  mcm4m3f_ca_w_2_400_s_0_300=7.52e-05 mcm4m3f_cc_w_2_400_s_0_300=9.23e-11 mcm4m3f_cf_w_2_400_s_0_300=1.10e-11
+  mcm4m3f_ca_w_2_400_s_0_360=7.52e-05 mcm4m3f_cc_w_2_400_s_0_360=8.49e-11 mcm4m3f_cf_w_2_400_s_0_360=1.28e-11
+  mcm4m3f_ca_w_2_400_s_0_450=7.52e-05 mcm4m3f_cc_w_2_400_s_0_450=7.53e-11 mcm4m3f_cf_w_2_400_s_0_450=1.55e-11
+  mcm4m3f_ca_w_2_400_s_0_600=7.52e-05 mcm4m3f_cc_w_2_400_s_0_600=6.22e-11 mcm4m3f_cf_w_2_400_s_0_600=1.96e-11
+  mcm4m3f_ca_w_2_400_s_0_800=7.52e-05 mcm4m3f_cc_w_2_400_s_0_800=4.89e-11 mcm4m3f_cf_w_2_400_s_0_800=2.45e-11
+  mcm4m3f_ca_w_2_400_s_1_000=7.52e-05 mcm4m3f_cc_w_2_400_s_1_000=3.92e-11 mcm4m3f_cf_w_2_400_s_1_000=2.88e-11
+  mcm4m3f_ca_w_2_400_s_1_200=7.52e-05 mcm4m3f_cc_w_2_400_s_1_200=3.17e-11 mcm4m3f_cf_w_2_400_s_1_200=3.25e-11
+  mcm4m3f_ca_w_2_400_s_2_100=7.52e-05 mcm4m3f_cc_w_2_400_s_2_100=1.42e-11 mcm4m3f_cf_w_2_400_s_2_100=4.41e-11
+  mcm4m3f_ca_w_2_400_s_3_300=7.52e-05 mcm4m3f_cc_w_2_400_s_3_300=5.71e-12 mcm4m3f_cf_w_2_400_s_3_300=5.14e-11
+  mcm4m3f_ca_w_2_400_s_9_000=7.52e-05 mcm4m3f_cc_w_2_400_s_9_000=1.35e-13 mcm4m3f_cf_w_2_400_s_9_000=5.67e-11
+  mcm4m3d_ca_w_0_300_s_0_300=7.67e-05 mcm4m3d_cc_w_0_300_s_0_300=8.27e-11 mcm4m3d_cf_w_0_300_s_0_300=1.11e-11
+  mcm4m3d_ca_w_0_300_s_0_360=7.67e-05 mcm4m3d_cc_w_0_300_s_0_360=7.60e-11 mcm4m3d_cf_w_0_300_s_0_360=1.30e-11
+  mcm4m3d_ca_w_0_300_s_0_450=7.67e-05 mcm4m3d_cc_w_0_300_s_0_450=6.71e-11 mcm4m3d_cf_w_0_300_s_0_450=1.57e-11
+  mcm4m3d_ca_w_0_300_s_0_600=7.67e-05 mcm4m3d_cc_w_0_300_s_0_600=5.49e-11 mcm4m3d_cf_w_0_300_s_0_600=1.99e-11
+  mcm4m3d_ca_w_0_300_s_0_800=7.67e-05 mcm4m3d_cc_w_0_300_s_0_800=4.28e-11 mcm4m3d_cf_w_0_300_s_0_800=2.48e-11
+  mcm4m3d_ca_w_0_300_s_1_000=7.67e-05 mcm4m3d_cc_w_0_300_s_1_000=3.38e-11 mcm4m3d_cf_w_0_300_s_1_000=2.92e-11
+  mcm4m3d_ca_w_0_300_s_1_200=7.67e-05 mcm4m3d_cc_w_0_300_s_1_200=2.70e-11 mcm4m3d_cf_w_0_300_s_1_200=3.29e-11
+  mcm4m3d_ca_w_0_300_s_2_100=7.67e-05 mcm4m3d_cc_w_0_300_s_2_100=1.12e-11 mcm4m3d_cf_w_0_300_s_2_100=4.40e-11
+  mcm4m3d_ca_w_0_300_s_3_300=7.67e-05 mcm4m3d_cc_w_0_300_s_3_300=3.99e-12 mcm4m3d_cf_w_0_300_s_3_300=5.02e-11
+  mcm4m3d_ca_w_0_300_s_9_000=7.67e-05 mcm4m3d_cc_w_0_300_s_9_000=5.50e-14 mcm4m3d_cf_w_0_300_s_9_000=5.41e-11
+  mcm4m3d_ca_w_2_400_s_0_300=7.67e-05 mcm4m3d_cc_w_2_400_s_0_300=9.11e-11 mcm4m3d_cf_w_2_400_s_0_300=1.12e-11
+  mcm4m3d_ca_w_2_400_s_0_360=7.67e-05 mcm4m3d_cc_w_2_400_s_0_360=8.37e-11 mcm4m3d_cf_w_2_400_s_0_360=1.31e-11
+  mcm4m3d_ca_w_2_400_s_0_450=7.67e-05 mcm4m3d_cc_w_2_400_s_0_450=7.42e-11 mcm4m3d_cf_w_2_400_s_0_450=1.58e-11
+  mcm4m3d_ca_w_2_400_s_0_600=7.67e-05 mcm4m3d_cc_w_2_400_s_0_600=6.10e-11 mcm4m3d_cf_w_2_400_s_0_600=2.00e-11
+  mcm4m3d_ca_w_2_400_s_0_800=7.67e-05 mcm4m3d_cc_w_2_400_s_0_800=4.77e-11 mcm4m3d_cf_w_2_400_s_0_800=2.50e-11
+  mcm4m3d_ca_w_2_400_s_1_000=7.67e-05 mcm4m3d_cc_w_2_400_s_1_000=3.79e-11 mcm4m3d_cf_w_2_400_s_1_000=2.94e-11
+  mcm4m3d_ca_w_2_400_s_1_200=7.67e-05 mcm4m3d_cc_w_2_400_s_1_200=3.05e-11 mcm4m3d_cf_w_2_400_s_1_200=3.33e-11
+  mcm4m3d_ca_w_2_400_s_2_100=7.67e-05 mcm4m3d_cc_w_2_400_s_2_100=1.32e-11 mcm4m3d_cf_w_2_400_s_2_100=4.49e-11
+  mcm4m3d_ca_w_2_400_s_3_300=7.67e-05 mcm4m3d_cc_w_2_400_s_3_300=4.92e-12 mcm4m3d_cf_w_2_400_s_3_300=5.20e-11
+  mcm4m3d_ca_w_2_400_s_9_000=7.67e-05 mcm4m3d_cc_w_2_400_s_9_000=1.05e-13 mcm4m3d_cf_w_2_400_s_9_000=5.67e-11
+  mcm4m3p1_ca_w_0_300_s_0_300=7.78e-05 mcm4m3p1_cc_w_0_300_s_0_300=8.24e-11 mcm4m3p1_cf_w_0_300_s_0_300=1.13e-11
+  mcm4m3p1_ca_w_0_300_s_0_360=7.78e-05 mcm4m3p1_cc_w_0_300_s_0_360=7.56e-11 mcm4m3p1_cf_w_0_300_s_0_360=1.32e-11
+  mcm4m3p1_ca_w_0_300_s_0_450=7.78e-05 mcm4m3p1_cc_w_0_300_s_0_450=6.68e-11 mcm4m3p1_cf_w_0_300_s_0_450=1.60e-11
+  mcm4m3p1_ca_w_0_300_s_0_600=7.78e-05 mcm4m3p1_cc_w_0_300_s_0_600=5.45e-11 mcm4m3p1_cf_w_0_300_s_0_600=2.02e-11
+  mcm4m3p1_ca_w_0_300_s_0_800=7.78e-05 mcm4m3p1_cc_w_0_300_s_0_800=4.24e-11 mcm4m3p1_cf_w_0_300_s_0_800=2.53e-11
+  mcm4m3p1_ca_w_0_300_s_1_000=7.78e-05 mcm4m3p1_cc_w_0_300_s_1_000=3.33e-11 mcm4m3p1_cf_w_0_300_s_1_000=2.96e-11
+  mcm4m3p1_ca_w_0_300_s_1_200=7.78e-05 mcm4m3p1_cc_w_0_300_s_1_200=2.65e-11 mcm4m3p1_cf_w_0_300_s_1_200=3.35e-11
+  mcm4m3p1_ca_w_0_300_s_2_100=7.78e-05 mcm4m3p1_cc_w_0_300_s_2_100=1.07e-11 mcm4m3p1_cf_w_0_300_s_2_100=4.46e-11
+  mcm4m3p1_ca_w_0_300_s_3_300=7.78e-05 mcm4m3p1_cc_w_0_300_s_3_300=3.72e-12 mcm4m3p1_cf_w_0_300_s_3_300=5.07e-11
+  mcm4m3p1_ca_w_0_300_s_9_000=7.78e-05 mcm4m3p1_cc_w_0_300_s_9_000=8.50e-14 mcm4m3p1_cf_w_0_300_s_9_000=5.43e-11
+  mcm4m3p1_ca_w_2_400_s_0_300=7.78e-05 mcm4m3p1_cc_w_2_400_s_0_300=9.03e-11 mcm4m3p1_cf_w_2_400_s_0_300=1.14e-11
+  mcm4m3p1_ca_w_2_400_s_0_360=7.78e-05 mcm4m3p1_cc_w_2_400_s_0_360=8.28e-11 mcm4m3p1_cf_w_2_400_s_0_360=1.33e-11
+  mcm4m3p1_ca_w_2_400_s_0_450=7.78e-05 mcm4m3p1_cc_w_2_400_s_0_450=7.32e-11 mcm4m3p1_cf_w_2_400_s_0_450=1.61e-11
+  mcm4m3p1_ca_w_2_400_s_0_600=7.78e-05 mcm4m3p1_cc_w_2_400_s_0_600=6.01e-11 mcm4m3p1_cf_w_2_400_s_0_600=2.04e-11
+  mcm4m3p1_ca_w_2_400_s_0_800=7.78e-05 mcm4m3p1_cc_w_2_400_s_0_800=4.68e-11 mcm4m3p1_cf_w_2_400_s_0_800=2.55e-11
+  mcm4m3p1_ca_w_2_400_s_1_000=7.78e-05 mcm4m3p1_cc_w_2_400_s_1_000=3.70e-11 mcm4m3p1_cf_w_2_400_s_1_000=3.00e-11
+  mcm4m3p1_ca_w_2_400_s_1_200=7.78e-05 mcm4m3p1_cc_w_2_400_s_1_200=2.96e-11 mcm4m3p1_cf_w_2_400_s_1_200=3.38e-11
+  mcm4m3p1_ca_w_2_400_s_2_100=7.78e-05 mcm4m3p1_cc_w_2_400_s_2_100=1.25e-11 mcm4m3p1_cf_w_2_400_s_2_100=4.55e-11
+  mcm4m3p1_ca_w_2_400_s_3_300=7.78e-05 mcm4m3p1_cc_w_2_400_s_3_300=4.44e-12 mcm4m3p1_cf_w_2_400_s_3_300=5.25e-11
+  mcm4m3p1_ca_w_2_400_s_9_000=7.78e-05 mcm4m3p1_cc_w_2_400_s_9_000=8.00e-14 mcm4m3p1_cf_w_2_400_s_9_000=5.68e-11
+  mcm4m3l1_ca_w_0_300_s_0_300=8.17e-05 mcm4m3l1_cc_w_0_300_s_0_300=8.11e-11 mcm4m3l1_cf_w_0_300_s_0_300=1.19e-11
+  mcm4m3l1_ca_w_0_300_s_0_360=8.17e-05 mcm4m3l1_cc_w_0_300_s_0_360=7.46e-11 mcm4m3l1_cf_w_0_300_s_0_360=1.39e-11
+  mcm4m3l1_ca_w_0_300_s_0_450=8.17e-05 mcm4m3l1_cc_w_0_300_s_0_450=6.57e-11 mcm4m3l1_cf_w_0_300_s_0_450=1.68e-11
+  mcm4m3l1_ca_w_0_300_s_0_600=8.17e-05 mcm4m3l1_cc_w_0_300_s_0_600=5.32e-11 mcm4m3l1_cf_w_0_300_s_0_600=2.13e-11
+  mcm4m3l1_ca_w_0_300_s_0_800=8.17e-05 mcm4m3l1_cc_w_0_300_s_0_800=4.09e-11 mcm4m3l1_cf_w_0_300_s_0_800=2.67e-11
+  mcm4m3l1_ca_w_0_300_s_1_000=8.17e-05 mcm4m3l1_cc_w_0_300_s_1_000=3.18e-11 mcm4m3l1_cf_w_0_300_s_1_000=3.12e-11
+  mcm4m3l1_ca_w_0_300_s_1_200=8.17e-05 mcm4m3l1_cc_w_0_300_s_1_200=2.49e-11 mcm4m3l1_cf_w_0_300_s_1_200=3.53e-11
+  mcm4m3l1_ca_w_0_300_s_2_100=8.17e-05 mcm4m3l1_cc_w_0_300_s_2_100=9.38e-12 mcm4m3l1_cf_w_0_300_s_2_100=4.65e-11
+  mcm4m3l1_ca_w_0_300_s_3_300=8.17e-05 mcm4m3l1_cc_w_0_300_s_3_300=2.84e-12 mcm4m3l1_cf_w_0_300_s_3_300=5.23e-11
+  mcm4m3l1_ca_w_0_300_s_9_000=8.17e-05 mcm4m3l1_cc_w_0_300_s_9_000=6.50e-14 mcm4m3l1_cf_w_0_300_s_9_000=5.51e-11
+  mcm4m3l1_ca_w_2_400_s_0_300=8.17e-05 mcm4m3l1_cc_w_2_400_s_0_300=8.76e-11 mcm4m3l1_cf_w_2_400_s_0_300=1.20e-11
+  mcm4m3l1_ca_w_2_400_s_0_360=8.17e-05 mcm4m3l1_cc_w_2_400_s_0_360=8.03e-11 mcm4m3l1_cf_w_2_400_s_0_360=1.40e-11
+  mcm4m3l1_ca_w_2_400_s_0_450=8.17e-05 mcm4m3l1_cc_w_2_400_s_0_450=7.06e-11 mcm4m3l1_cf_w_2_400_s_0_450=1.70e-11
+  mcm4m3l1_ca_w_2_400_s_0_600=8.17e-05 mcm4m3l1_cc_w_2_400_s_0_600=5.74e-11 mcm4m3l1_cf_w_2_400_s_0_600=2.15e-11
+  mcm4m3l1_ca_w_2_400_s_0_800=8.17e-05 mcm4m3l1_cc_w_2_400_s_0_800=4.41e-11 mcm4m3l1_cf_w_2_400_s_0_800=2.69e-11
+  mcm4m3l1_ca_w_2_400_s_1_000=8.17e-05 mcm4m3l1_cc_w_2_400_s_1_000=3.44e-11 mcm4m3l1_cf_w_2_400_s_1_000=3.16e-11
+  mcm4m3l1_ca_w_2_400_s_1_200=8.17e-05 mcm4m3l1_cc_w_2_400_s_1_200=2.71e-11 mcm4m3l1_cf_w_2_400_s_1_200=3.56e-11
+  mcm4m3l1_ca_w_2_400_s_2_100=8.17e-05 mcm4m3l1_cc_w_2_400_s_2_100=1.04e-11 mcm4m3l1_cf_w_2_400_s_2_100=4.74e-11
+  mcm4m3l1_ca_w_2_400_s_3_300=8.17e-05 mcm4m3l1_cc_w_2_400_s_3_300=3.23e-12 mcm4m3l1_cf_w_2_400_s_3_300=5.39e-11
+  mcm4m3l1_ca_w_2_400_s_9_000=8.17e-05 mcm4m3l1_cc_w_2_400_s_9_000=5.50e-14 mcm4m3l1_cf_w_2_400_s_9_000=5.71e-11
+  mcm4m3m1_ca_w_0_300_s_0_300=9.19e-05 mcm4m3m1_cc_w_0_300_s_0_300=7.91e-11 mcm4m3m1_cf_w_0_300_s_0_300=1.35e-11
+  mcm4m3m1_ca_w_0_300_s_0_360=9.19e-05 mcm4m3m1_cc_w_0_300_s_0_360=7.21e-11 mcm4m3m1_cf_w_0_300_s_0_360=1.58e-11
+  mcm4m3m1_ca_w_0_300_s_0_450=9.19e-05 mcm4m3m1_cc_w_0_300_s_0_450=6.30e-11 mcm4m3m1_cf_w_0_300_s_0_450=1.91e-11
+  mcm4m3m1_ca_w_0_300_s_0_600=9.19e-05 mcm4m3m1_cc_w_0_300_s_0_600=5.02e-11 mcm4m3m1_cf_w_0_300_s_0_600=2.41e-11
+  mcm4m3m1_ca_w_0_300_s_0_800=9.19e-05 mcm4m3m1_cc_w_0_300_s_0_800=3.77e-11 mcm4m3m1_cf_w_0_300_s_0_800=3.01e-11
+  mcm4m3m1_ca_w_0_300_s_1_000=9.19e-05 mcm4m3m1_cc_w_0_300_s_1_000=2.84e-11 mcm4m3m1_cf_w_0_300_s_1_000=3.53e-11
+  mcm4m3m1_ca_w_0_300_s_1_200=9.19e-05 mcm4m3m1_cc_w_0_300_s_1_200=2.16e-11 mcm4m3m1_cf_w_0_300_s_1_200=3.95e-11
+  mcm4m3m1_ca_w_0_300_s_2_100=9.19e-05 mcm4m3m1_cc_w_0_300_s_2_100=6.82e-12 mcm4m3m1_cf_w_0_300_s_2_100=5.09e-11
+  mcm4m3m1_ca_w_0_300_s_3_300=9.19e-05 mcm4m3m1_cc_w_0_300_s_3_300=1.60e-12 mcm4m3m1_cf_w_0_300_s_3_300=5.59e-11
+  mcm4m3m1_ca_w_0_300_s_9_000=9.19e-05 mcm4m3m1_cc_w_0_300_s_9_000=3.00e-14 mcm4m3m1_cf_w_0_300_s_9_000=5.75e-11
+  mcm4m3m1_ca_w_2_400_s_0_300=9.19e-05 mcm4m3m1_cc_w_2_400_s_0_300=8.27e-11 mcm4m3m1_cf_w_2_400_s_0_300=1.36e-11
+  mcm4m3m1_ca_w_2_400_s_0_360=9.19e-05 mcm4m3m1_cc_w_2_400_s_0_360=7.54e-11 mcm4m3m1_cf_w_2_400_s_0_360=1.59e-11
+  mcm4m3m1_ca_w_2_400_s_0_450=9.19e-05 mcm4m3m1_cc_w_2_400_s_0_450=6.58e-11 mcm4m3m1_cf_w_2_400_s_0_450=1.92e-11
+  mcm4m3m1_ca_w_2_400_s_0_600=9.19e-05 mcm4m3m1_cc_w_2_400_s_0_600=5.26e-11 mcm4m3m1_cf_w_2_400_s_0_600=2.43e-11
+  mcm4m3m1_ca_w_2_400_s_0_800=9.19e-05 mcm4m3m1_cc_w_2_400_s_0_800=3.93e-11 mcm4m3m1_cf_w_2_400_s_0_800=3.04e-11
+  mcm4m3m1_ca_w_2_400_s_1_000=9.19e-05 mcm4m3m1_cc_w_2_400_s_1_000=2.96e-11 mcm4m3m1_cf_w_2_400_s_1_000=3.56e-11
+  mcm4m3m1_ca_w_2_400_s_1_200=9.19e-05 mcm4m3m1_cc_w_2_400_s_1_200=2.26e-11 mcm4m3m1_cf_w_2_400_s_1_200=3.99e-11
+  mcm4m3m1_ca_w_2_400_s_2_100=9.19e-05 mcm4m3m1_cc_w_2_400_s_2_100=7.25e-12 mcm4m3m1_cf_w_2_400_s_2_100=5.18e-11
+  mcm4m3m1_ca_w_2_400_s_3_300=9.19e-05 mcm4m3m1_cc_w_2_400_s_3_300=1.70e-12 mcm4m3m1_cf_w_2_400_s_3_300=5.70e-11
+  mcm4m3m1_ca_w_2_400_s_9_000=9.19e-05 mcm4m3m1_cc_w_2_400_s_9_000=0.00e+00 mcm4m3m1_cf_w_2_400_s_9_000=5.87e-11
+  mcm4m3m2_ca_w_0_300_s_0_300=1.29e-04 mcm4m3m2_cc_w_0_300_s_0_300=7.22e-11 mcm4m3m2_cf_w_0_300_s_0_300=1.90e-11
+  mcm4m3m2_ca_w_0_300_s_0_360=1.29e-04 mcm4m3m2_cc_w_0_300_s_0_360=6.52e-11 mcm4m3m2_cf_w_0_300_s_0_360=2.20e-11
+  mcm4m3m2_ca_w_0_300_s_0_450=1.29e-04 mcm4m3m2_cc_w_0_300_s_0_450=5.59e-11 mcm4m3m2_cf_w_0_300_s_0_450=2.64e-11
+  mcm4m3m2_ca_w_0_300_s_0_600=1.29e-04 mcm4m3m2_cc_w_0_300_s_0_600=4.30e-11 mcm4m3m2_cf_w_0_300_s_0_600=3.30e-11
+  mcm4m3m2_ca_w_0_300_s_0_800=1.29e-04 mcm4m3m2_cc_w_0_300_s_0_800=3.04e-11 mcm4m3m2_cf_w_0_300_s_0_800=4.06e-11
+  mcm4m3m2_ca_w_0_300_s_1_000=1.29e-04 mcm4m3m2_cc_w_0_300_s_1_000=2.14e-11 mcm4m3m2_cf_w_0_300_s_1_000=4.67e-11
+  mcm4m3m2_ca_w_0_300_s_1_200=1.29e-04 mcm4m3m2_cc_w_0_300_s_1_200=1.50e-11 mcm4m3m2_cf_w_0_300_s_1_200=5.15e-11
+  mcm4m3m2_ca_w_0_300_s_2_100=1.29e-04 mcm4m3m2_cc_w_0_300_s_2_100=3.27e-12 mcm4m3m2_cf_w_0_300_s_2_100=6.18e-11
+  mcm4m3m2_ca_w_0_300_s_3_300=1.29e-04 mcm4m3m2_cc_w_0_300_s_3_300=5.00e-13 mcm4m3m2_cf_w_0_300_s_3_300=6.46e-11
+  mcm4m3m2_ca_w_0_300_s_9_000=1.29e-04 mcm4m3m2_cc_w_0_300_s_9_000=3.50e-14 mcm4m3m2_cf_w_0_300_s_9_000=6.51e-11
+  mcm4m3m2_ca_w_2_400_s_0_300=1.29e-04 mcm4m3m2_cc_w_2_400_s_0_300=7.34e-11 mcm4m3m2_cf_w_2_400_s_0_300=1.90e-11
+  mcm4m3m2_ca_w_2_400_s_0_360=1.29e-04 mcm4m3m2_cc_w_2_400_s_0_360=6.62e-11 mcm4m3m2_cf_w_2_400_s_0_360=2.21e-11
+  mcm4m3m2_ca_w_2_400_s_0_450=1.29e-04 mcm4m3m2_cc_w_2_400_s_0_450=5.66e-11 mcm4m3m2_cf_w_2_400_s_0_450=2.66e-11
+  mcm4m3m2_ca_w_2_400_s_0_600=1.29e-04 mcm4m3m2_cc_w_2_400_s_0_600=4.37e-11 mcm4m3m2_cf_w_2_400_s_0_600=3.32e-11
+  mcm4m3m2_ca_w_2_400_s_0_800=1.29e-04 mcm4m3m2_cc_w_2_400_s_0_800=3.08e-11 mcm4m3m2_cf_w_2_400_s_0_800=4.08e-11
+  mcm4m3m2_ca_w_2_400_s_1_000=1.29e-04 mcm4m3m2_cc_w_2_400_s_1_000=2.18e-11 mcm4m3m2_cf_w_2_400_s_1_000=4.71e-11
+  mcm4m3m2_ca_w_2_400_s_1_200=1.29e-04 mcm4m3m2_cc_w_2_400_s_1_200=1.53e-11 mcm4m3m2_cf_w_2_400_s_1_200=5.19e-11
+  mcm4m3m2_ca_w_2_400_s_2_100=1.29e-04 mcm4m3m2_cc_w_2_400_s_2_100=3.30e-12 mcm4m3m2_cf_w_2_400_s_2_100=6.25e-11
+  mcm4m3m2_ca_w_2_400_s_3_300=1.29e-04 mcm4m3m2_cc_w_2_400_s_3_300=4.50e-13 mcm4m3m2_cf_w_2_400_s_3_300=6.53e-11
+  mcm4m3m2_ca_w_2_400_s_9_000=1.29e-04 mcm4m3m2_cc_w_2_400_s_9_000=0.00e+00 mcm4m3m2_cf_w_2_400_s_9_000=6.59e-11
+  mcm5m3f_ca_w_0_300_s_0_300=2.83e-05 mcm5m3f_cc_w_0_300_s_0_300=9.12e-11 mcm5m3f_cf_w_0_300_s_0_300=4.56e-12
+  mcm5m3f_ca_w_0_300_s_0_360=2.83e-05 mcm5m3f_cc_w_0_300_s_0_360=8.50e-11 mcm5m3f_cf_w_0_300_s_0_360=5.37e-12
+  mcm5m3f_ca_w_0_300_s_0_450=2.83e-05 mcm5m3f_cc_w_0_300_s_0_450=7.66e-11 mcm5m3f_cf_w_0_300_s_0_450=6.61e-12
+  mcm5m3f_ca_w_0_300_s_0_600=2.83e-05 mcm5m3f_cc_w_0_300_s_0_600=6.53e-11 mcm5m3f_cf_w_0_300_s_0_600=8.59e-12
+  mcm5m3f_ca_w_0_300_s_0_800=2.83e-05 mcm5m3f_cc_w_0_300_s_0_800=5.39e-11 mcm5m3f_cf_w_0_300_s_0_800=1.10e-11
+  mcm5m3f_ca_w_0_300_s_1_000=2.83e-05 mcm5m3f_cc_w_0_300_s_1_000=4.51e-11 mcm5m3f_cf_w_0_300_s_1_000=1.34e-11
+  mcm5m3f_ca_w_0_300_s_1_200=2.83e-05 mcm5m3f_cc_w_0_300_s_1_200=3.80e-11 mcm5m3f_cf_w_0_300_s_1_200=1.56e-11
+  mcm5m3f_ca_w_0_300_s_2_100=2.83e-05 mcm5m3f_cc_w_0_300_s_2_100=2.05e-11 mcm5m3f_cf_w_0_300_s_2_100=2.40e-11
+  mcm5m3f_ca_w_0_300_s_3_300=2.83e-05 mcm5m3f_cc_w_0_300_s_3_300=1.01e-11 mcm5m3f_cf_w_0_300_s_3_300=3.12e-11
+  mcm5m3f_ca_w_0_300_s_9_000=2.83e-05 mcm5m3f_cc_w_0_300_s_9_000=5.05e-13 mcm5m3f_cf_w_0_300_s_9_000=3.97e-11
+  mcm5m3f_ca_w_2_400_s_0_300=2.83e-05 mcm5m3f_cc_w_2_400_s_0_300=1.06e-10 mcm5m3f_cf_w_2_400_s_0_300=4.61e-12
+  mcm5m3f_ca_w_2_400_s_0_360=2.83e-05 mcm5m3f_cc_w_2_400_s_0_360=9.88e-11 mcm5m3f_cf_w_2_400_s_0_360=5.42e-12
+  mcm5m3f_ca_w_2_400_s_0_450=2.83e-05 mcm5m3f_cc_w_2_400_s_0_450=8.90e-11 mcm5m3f_cf_w_2_400_s_0_450=6.61e-12
+  mcm5m3f_ca_w_2_400_s_0_600=2.83e-05 mcm5m3f_cc_w_2_400_s_0_600=7.57e-11 mcm5m3f_cf_w_2_400_s_0_600=8.57e-12
+  mcm5m3f_ca_w_2_400_s_0_800=2.83e-05 mcm5m3f_cc_w_2_400_s_0_800=6.22e-11 mcm5m3f_cf_w_2_400_s_0_800=1.11e-11
+  mcm5m3f_ca_w_2_400_s_1_000=2.83e-05 mcm5m3f_cc_w_2_400_s_1_000=5.20e-11 mcm5m3f_cf_w_2_400_s_1_000=1.35e-11
+  mcm5m3f_ca_w_2_400_s_1_200=2.83e-05 mcm5m3f_cc_w_2_400_s_1_200=4.41e-11 mcm5m3f_cf_w_2_400_s_1_200=1.58e-11
+  mcm5m3f_ca_w_2_400_s_2_100=2.83e-05 mcm5m3f_cc_w_2_400_s_2_100=2.41e-11 mcm5m3f_cf_w_2_400_s_2_100=2.46e-11
+  mcm5m3f_ca_w_2_400_s_3_300=2.83e-05 mcm5m3f_cc_w_2_400_s_3_300=1.21e-11 mcm5m3f_cf_w_2_400_s_3_300=3.26e-11
+  mcm5m3f_ca_w_2_400_s_9_000=2.83e-05 mcm5m3f_cc_w_2_400_s_9_000=5.90e-13 mcm5m3f_cf_w_2_400_s_9_000=4.28e-11
+  mcm5m3d_ca_w_0_300_s_0_300=2.98e-05 mcm5m3d_cc_w_0_300_s_0_300=9.08e-11 mcm5m3d_cf_w_0_300_s_0_300=4.80e-12
+  mcm5m3d_ca_w_0_300_s_0_360=2.98e-05 mcm5m3d_cc_w_0_300_s_0_360=8.46e-11 mcm5m3d_cf_w_0_300_s_0_360=5.66e-12
+  mcm5m3d_ca_w_0_300_s_0_450=2.98e-05 mcm5m3d_cc_w_0_300_s_0_450=7.61e-11 mcm5m3d_cf_w_0_300_s_0_450=6.95e-12
+  mcm5m3d_ca_w_0_300_s_0_600=2.98e-05 mcm5m3d_cc_w_0_300_s_0_600=6.48e-11 mcm5m3d_cf_w_0_300_s_0_600=9.03e-12
+  mcm5m3d_ca_w_0_300_s_0_800=2.98e-05 mcm5m3d_cc_w_0_300_s_0_800=5.33e-11 mcm5m3d_cf_w_0_300_s_0_800=1.16e-11
+  mcm5m3d_ca_w_0_300_s_1_000=2.98e-05 mcm5m3d_cc_w_0_300_s_1_000=4.43e-11 mcm5m3d_cf_w_0_300_s_1_000=1.40e-11
+  mcm5m3d_ca_w_0_300_s_1_200=2.98e-05 mcm5m3d_cc_w_0_300_s_1_200=3.74e-11 mcm5m3d_cf_w_0_300_s_1_200=1.64e-11
+  mcm5m3d_ca_w_0_300_s_2_100=2.98e-05 mcm5m3d_cc_w_0_300_s_2_100=1.97e-11 mcm5m3d_cf_w_0_300_s_2_100=2.51e-11
+  mcm5m3d_ca_w_0_300_s_3_300=2.98e-05 mcm5m3d_cc_w_0_300_s_3_300=9.43e-12 mcm5m3d_cf_w_0_300_s_3_300=3.23e-11
+  mcm5m3d_ca_w_0_300_s_9_000=2.98e-05 mcm5m3d_cc_w_0_300_s_9_000=3.95e-13 mcm5m3d_cf_w_0_300_s_9_000=4.04e-11
+  mcm5m3d_ca_w_2_400_s_0_300=2.98e-05 mcm5m3d_cc_w_2_400_s_0_300=1.05e-10 mcm5m3d_cf_w_2_400_s_0_300=4.85e-12
+  mcm5m3d_ca_w_2_400_s_0_360=2.98e-05 mcm5m3d_cc_w_2_400_s_0_360=9.77e-11 mcm5m3d_cf_w_2_400_s_0_360=5.70e-12
+  mcm5m3d_ca_w_2_400_s_0_450=2.98e-05 mcm5m3d_cc_w_2_400_s_0_450=8.78e-11 mcm5m3d_cf_w_2_400_s_0_450=6.97e-12
+  mcm5m3d_ca_w_2_400_s_0_600=2.98e-05 mcm5m3d_cc_w_2_400_s_0_600=7.45e-11 mcm5m3d_cf_w_2_400_s_0_600=9.02e-12
+  mcm5m3d_ca_w_2_400_s_0_800=2.98e-05 mcm5m3d_cc_w_2_400_s_0_800=6.10e-11 mcm5m3d_cf_w_2_400_s_0_800=1.17e-11
+  mcm5m3d_ca_w_2_400_s_1_000=2.98e-05 mcm5m3d_cc_w_2_400_s_1_000=5.07e-11 mcm5m3d_cf_w_2_400_s_1_000=1.42e-11
+  mcm5m3d_ca_w_2_400_s_1_200=2.98e-05 mcm5m3d_cc_w_2_400_s_1_200=4.28e-11 mcm5m3d_cf_w_2_400_s_1_200=1.66e-11
+  mcm5m3d_ca_w_2_400_s_2_100=2.98e-05 mcm5m3d_cc_w_2_400_s_2_100=2.29e-11 mcm5m3d_cf_w_2_400_s_2_100=2.57e-11
+  mcm5m3d_ca_w_2_400_s_3_300=2.98e-05 mcm5m3d_cc_w_2_400_s_3_300=1.11e-11 mcm5m3d_cf_w_2_400_s_3_300=3.38e-11
+  mcm5m3d_ca_w_2_400_s_9_000=2.98e-05 mcm5m3d_cc_w_2_400_s_9_000=4.50e-13 mcm5m3d_cf_w_2_400_s_9_000=4.33e-11
+  mcm5m3p1_ca_w_0_300_s_0_300=3.10e-05 mcm5m3p1_cc_w_0_300_s_0_300=9.05e-11 mcm5m3p1_cf_w_0_300_s_0_300=4.99e-12
+  mcm5m3p1_ca_w_0_300_s_0_360=3.10e-05 mcm5m3p1_cc_w_0_300_s_0_360=8.43e-11 mcm5m3p1_cf_w_0_300_s_0_360=5.88e-12
+  mcm5m3p1_ca_w_0_300_s_0_450=3.10e-05 mcm5m3p1_cc_w_0_300_s_0_450=7.61e-11 mcm5m3p1_cf_w_0_300_s_0_450=7.22e-12
+  mcm5m3p1_ca_w_0_300_s_0_600=3.10e-05 mcm5m3p1_cc_w_0_300_s_0_600=6.44e-11 mcm5m3p1_cf_w_0_300_s_0_600=9.38e-12
+  mcm5m3p1_ca_w_0_300_s_0_800=3.10e-05 mcm5m3p1_cc_w_0_300_s_0_800=5.27e-11 mcm5m3p1_cf_w_0_300_s_0_800=1.20e-11
+  mcm5m3p1_ca_w_0_300_s_1_000=3.10e-05 mcm5m3p1_cc_w_0_300_s_1_000=4.39e-11 mcm5m3p1_cf_w_0_300_s_1_000=1.46e-11
+  mcm5m3p1_ca_w_0_300_s_1_200=3.10e-05 mcm5m3p1_cc_w_0_300_s_1_200=3.68e-11 mcm5m3p1_cf_w_0_300_s_1_200=1.69e-11
+  mcm5m3p1_ca_w_0_300_s_2_100=3.10e-05 mcm5m3p1_cc_w_0_300_s_2_100=1.91e-11 mcm5m3p1_cf_w_0_300_s_2_100=2.58e-11
+  mcm5m3p1_ca_w_0_300_s_3_300=3.10e-05 mcm5m3p1_cc_w_0_300_s_3_300=8.93e-12 mcm5m3p1_cf_w_0_300_s_3_300=3.32e-11
+  mcm5m3p1_ca_w_0_300_s_9_000=3.10e-05 mcm5m3p1_cc_w_0_300_s_9_000=3.40e-13 mcm5m3p1_cf_w_0_300_s_9_000=4.09e-11
+  mcm5m3p1_ca_w_2_400_s_0_300=3.10e-05 mcm5m3p1_cc_w_2_400_s_0_300=1.04e-10 mcm5m3p1_cf_w_2_400_s_0_300=5.06e-12
+  mcm5m3p1_ca_w_2_400_s_0_360=3.10e-05 mcm5m3p1_cc_w_2_400_s_0_360=9.66e-11 mcm5m3p1_cf_w_2_400_s_0_360=5.96e-12
+  mcm5m3p1_ca_w_2_400_s_0_450=3.10e-05 mcm5m3p1_cc_w_2_400_s_0_450=8.70e-11 mcm5m3p1_cf_w_2_400_s_0_450=7.26e-12
+  mcm5m3p1_ca_w_2_400_s_0_600=3.10e-05 mcm5m3p1_cc_w_2_400_s_0_600=7.36e-11 mcm5m3p1_cf_w_2_400_s_0_600=9.38e-12
+  mcm5m3p1_ca_w_2_400_s_0_800=3.10e-05 mcm5m3p1_cc_w_2_400_s_0_800=6.01e-11 mcm5m3p1_cf_w_2_400_s_0_800=1.21e-11
+  mcm5m3p1_ca_w_2_400_s_1_000=3.10e-05 mcm5m3p1_cc_w_2_400_s_1_000=4.98e-11 mcm5m3p1_cf_w_2_400_s_1_000=1.48e-11
+  mcm5m3p1_ca_w_2_400_s_1_200=3.10e-05 mcm5m3p1_cc_w_2_400_s_1_200=4.20e-11 mcm5m3p1_cf_w_2_400_s_1_200=1.72e-11
+  mcm5m3p1_ca_w_2_400_s_2_100=3.10e-05 mcm5m3p1_cc_w_2_400_s_2_100=2.20e-11 mcm5m3p1_cf_w_2_400_s_2_100=2.65e-11
+  mcm5m3p1_ca_w_2_400_s_3_300=3.10e-05 mcm5m3p1_cc_w_2_400_s_3_300=1.04e-11 mcm5m3p1_cf_w_2_400_s_3_300=3.47e-11
+  mcm5m3p1_ca_w_2_400_s_9_000=3.10e-05 mcm5m3p1_cc_w_2_400_s_9_000=3.90e-13 mcm5m3p1_cf_w_2_400_s_9_000=4.37e-11
+  mcm5m3l1_ca_w_0_300_s_0_300=3.48e-05 mcm5m3l1_cc_w_0_300_s_0_300=8.96e-11 mcm5m3l1_cf_w_0_300_s_0_300=5.60e-12
+  mcm5m3l1_ca_w_0_300_s_0_360=3.48e-05 mcm5m3l1_cc_w_0_300_s_0_360=8.33e-11 mcm5m3l1_cf_w_0_300_s_0_360=6.60e-12
+  mcm5m3l1_ca_w_0_300_s_0_450=3.48e-05 mcm5m3l1_cc_w_0_300_s_0_450=7.50e-11 mcm5m3l1_cf_w_0_300_s_0_450=8.09e-12
+  mcm5m3l1_ca_w_0_300_s_0_600=3.48e-05 mcm5m3l1_cc_w_0_300_s_0_600=6.31e-11 mcm5m3l1_cf_w_0_300_s_0_600=1.05e-11
+  mcm5m3l1_ca_w_0_300_s_0_800=3.48e-05 mcm5m3l1_cc_w_0_300_s_0_800=5.13e-11 mcm5m3l1_cf_w_0_300_s_0_800=1.34e-11
+  mcm5m3l1_ca_w_0_300_s_1_000=3.48e-05 mcm5m3l1_cc_w_0_300_s_1_000=4.21e-11 mcm5m3l1_cf_w_0_300_s_1_000=1.62e-11
+  mcm5m3l1_ca_w_0_300_s_1_200=3.48e-05 mcm5m3l1_cc_w_0_300_s_1_200=3.51e-11 mcm5m3l1_cf_w_0_300_s_1_200=1.88e-11
+  mcm5m3l1_ca_w_0_300_s_2_100=3.48e-05 mcm5m3l1_cc_w_0_300_s_2_100=1.74e-11 mcm5m3l1_cf_w_0_300_s_2_100=2.83e-11
+  mcm5m3l1_ca_w_0_300_s_3_300=3.48e-05 mcm5m3l1_cc_w_0_300_s_3_300=7.56e-12 mcm5m3l1_cf_w_0_300_s_3_300=3.57e-11
+  mcm5m3l1_ca_w_0_300_s_9_000=3.48e-05 mcm5m3l1_cc_w_0_300_s_9_000=2.10e-13 mcm5m3l1_cf_w_0_300_s_9_000=4.25e-11
+  mcm5m3l1_ca_w_2_400_s_0_300=3.48e-05 mcm5m3l1_cc_w_2_400_s_0_300=1.02e-10 mcm5m3l1_cf_w_2_400_s_0_300=5.66e-12
+  mcm5m3l1_ca_w_2_400_s_0_360=3.48e-05 mcm5m3l1_cc_w_2_400_s_0_360=9.42e-11 mcm5m3l1_cf_w_2_400_s_0_360=6.64e-12
+  mcm5m3l1_ca_w_2_400_s_0_450=3.48e-05 mcm5m3l1_cc_w_2_400_s_0_450=8.43e-11 mcm5m3l1_cf_w_2_400_s_0_450=8.11e-12
+  mcm5m3l1_ca_w_2_400_s_0_600=3.48e-05 mcm5m3l1_cc_w_2_400_s_0_600=7.09e-11 mcm5m3l1_cf_w_2_400_s_0_600=1.05e-11
+  mcm5m3l1_ca_w_2_400_s_0_800=3.48e-05 mcm5m3l1_cc_w_2_400_s_0_800=5.75e-11 mcm5m3l1_cf_w_2_400_s_0_800=1.35e-11
+  mcm5m3l1_ca_w_2_400_s_1_000=3.48e-05 mcm5m3l1_cc_w_2_400_s_1_000=4.72e-11 mcm5m3l1_cf_w_2_400_s_1_000=1.64e-11
+  mcm5m3l1_ca_w_2_400_s_1_200=3.48e-05 mcm5m3l1_cc_w_2_400_s_1_200=3.94e-11 mcm5m3l1_cf_w_2_400_s_1_200=1.92e-11
+  mcm5m3l1_ca_w_2_400_s_2_100=3.48e-05 mcm5m3l1_cc_w_2_400_s_2_100=1.97e-11 mcm5m3l1_cf_w_2_400_s_2_100=2.91e-11
+  mcm5m3l1_ca_w_2_400_s_3_300=3.48e-05 mcm5m3l1_cc_w_2_400_s_3_300=8.65e-12 mcm5m3l1_cf_w_2_400_s_3_300=3.72e-11
+  mcm5m3l1_ca_w_2_400_s_9_000=3.48e-05 mcm5m3l1_cc_w_2_400_s_9_000=2.50e-13 mcm5m3l1_cf_w_2_400_s_9_000=4.50e-11
+  mcm5m3m1_ca_w_0_300_s_0_300=4.50e-05 mcm5m3m1_cc_w_0_300_s_0_300=8.72e-11 mcm5m3m1_cf_w_0_300_s_0_300=7.19e-12
+  mcm5m3m1_ca_w_0_300_s_0_360=4.50e-05 mcm5m3m1_cc_w_0_300_s_0_360=8.07e-11 mcm5m3m1_cf_w_0_300_s_0_360=8.44e-12
+  mcm5m3m1_ca_w_0_300_s_0_450=4.50e-05 mcm5m3m1_cc_w_0_300_s_0_450=7.20e-11 mcm5m3m1_cf_w_0_300_s_0_450=1.03e-11
+  mcm5m3m1_ca_w_0_300_s_0_600=4.50e-05 mcm5m3m1_cc_w_0_300_s_0_600=6.01e-11 mcm5m3m1_cf_w_0_300_s_0_600=1.33e-11
+  mcm5m3m1_ca_w_0_300_s_0_800=4.50e-05 mcm5m3m1_cc_w_0_300_s_0_800=4.80e-11 mcm5m3m1_cf_w_0_300_s_0_800=1.69e-11
+  mcm5m3m1_ca_w_0_300_s_1_000=4.50e-05 mcm5m3m1_cc_w_0_300_s_1_000=3.87e-11 mcm5m3m1_cf_w_0_300_s_1_000=2.03e-11
+  mcm5m3m1_ca_w_0_300_s_1_200=4.50e-05 mcm5m3m1_cc_w_0_300_s_1_200=3.15e-11 mcm5m3m1_cf_w_0_300_s_1_200=2.34e-11
+  mcm5m3m1_ca_w_0_300_s_2_100=4.50e-05 mcm5m3m1_cc_w_0_300_s_2_100=1.42e-11 mcm5m3m1_cf_w_0_300_s_2_100=3.39e-11
+  mcm5m3m1_ca_w_0_300_s_3_300=4.50e-05 mcm5m3m1_cc_w_0_300_s_3_300=5.33e-12 mcm5m3m1_cf_w_0_300_s_3_300=4.12e-11
+  mcm5m3m1_ca_w_0_300_s_9_000=4.50e-05 mcm5m3m1_cc_w_0_300_s_9_000=8.50e-14 mcm5m3m1_cf_w_0_300_s_9_000=4.62e-11
+  mcm5m3m1_ca_w_2_400_s_0_300=4.50e-05 mcm5m3m1_cc_w_2_400_s_0_300=9.67e-11 mcm5m3m1_cf_w_2_400_s_0_300=7.22e-12
+  mcm5m3m1_ca_w_2_400_s_0_360=4.50e-05 mcm5m3m1_cc_w_2_400_s_0_360=8.93e-11 mcm5m3m1_cf_w_2_400_s_0_360=8.47e-12
+  mcm5m3m1_ca_w_2_400_s_0_450=4.50e-05 mcm5m3m1_cc_w_2_400_s_0_450=7.93e-11 mcm5m3m1_cf_w_2_400_s_0_450=1.03e-11
+  mcm5m3m1_ca_w_2_400_s_0_600=4.50e-05 mcm5m3m1_cc_w_2_400_s_0_600=6.59e-11 mcm5m3m1_cf_w_2_400_s_0_600=1.33e-11
+  mcm5m3m1_ca_w_2_400_s_0_800=4.50e-05 mcm5m3m1_cc_w_2_400_s_0_800=5.25e-11 mcm5m3m1_cf_w_2_400_s_0_800=1.70e-11
+  mcm5m3m1_ca_w_2_400_s_1_000=4.50e-05 mcm5m3m1_cc_w_2_400_s_1_000=4.25e-11 mcm5m3m1_cf_w_2_400_s_1_000=2.06e-11
+  mcm5m3m1_ca_w_2_400_s_1_200=4.50e-05 mcm5m3m1_cc_w_2_400_s_1_200=3.47e-11 mcm5m3m1_cf_w_2_400_s_1_200=2.38e-11
+  mcm5m3m1_ca_w_2_400_s_2_100=4.50e-05 mcm5m3m1_cc_w_2_400_s_2_100=1.58e-11 mcm5m3m1_cf_w_2_400_s_2_100=3.48e-11
+  mcm5m3m1_ca_w_2_400_s_3_300=4.50e-05 mcm5m3m1_cc_w_2_400_s_3_300=6.00e-12 mcm5m3m1_cf_w_2_400_s_3_300=4.27e-11
+  mcm5m3m1_ca_w_2_400_s_9_000=4.50e-05 mcm5m3m1_cc_w_2_400_s_9_000=1.40e-13 mcm5m3m1_cf_w_2_400_s_9_000=4.83e-11
+  mcm5m3m2_ca_w_0_300_s_0_300=8.23e-05 mcm5m3m2_cc_w_0_300_s_0_300=8.05e-11 mcm5m3m2_cf_w_0_300_s_0_300=1.26e-11
+  mcm5m3m2_ca_w_0_300_s_0_360=8.23e-05 mcm5m3m2_cc_w_0_300_s_0_360=7.39e-11 mcm5m3m2_cf_w_0_300_s_0_360=1.47e-11
+  mcm5m3m2_ca_w_0_300_s_0_450=8.23e-05 mcm5m3m2_cc_w_0_300_s_0_450=6.49e-11 mcm5m3m2_cf_w_0_300_s_0_450=1.77e-11
+  mcm5m3m2_ca_w_0_300_s_0_600=8.23e-05 mcm5m3m2_cc_w_0_300_s_0_600=5.28e-11 mcm5m3m2_cf_w_0_300_s_0_600=2.23e-11
+  mcm5m3m2_ca_w_0_300_s_0_800=8.23e-05 mcm5m3m2_cc_w_0_300_s_0_800=4.06e-11 mcm5m3m2_cf_w_0_300_s_0_800=2.76e-11
+  mcm5m3m2_ca_w_0_300_s_1_000=8.23e-05 mcm5m3m2_cc_w_0_300_s_1_000=3.15e-11 mcm5m3m2_cf_w_0_300_s_1_000=3.23e-11
+  mcm5m3m2_ca_w_0_300_s_1_200=8.23e-05 mcm5m3m2_cc_w_0_300_s_1_200=2.46e-11 mcm5m3m2_cf_w_0_300_s_1_200=3.64e-11
+  mcm5m3m2_ca_w_0_300_s_2_100=8.23e-05 mcm5m3m2_cc_w_0_300_s_2_100=9.11e-12 mcm5m3m2_cf_w_0_300_s_2_100=4.77e-11
+  mcm5m3m2_ca_w_0_300_s_3_300=8.23e-05 mcm5m3m2_cc_w_0_300_s_3_300=2.76e-12 mcm5m3m2_cf_w_0_300_s_3_300=5.35e-11
+  mcm5m3m2_ca_w_0_300_s_9_000=8.23e-05 mcm5m3m2_cc_w_0_300_s_9_000=5.50e-14 mcm5m3m2_cf_w_0_300_s_9_000=5.62e-11
+  mcm5m3m2_ca_w_2_400_s_0_300=8.23e-05 mcm5m3m2_cc_w_2_400_s_0_300=8.72e-11 mcm5m3m2_cf_w_2_400_s_0_300=1.27e-11
+  mcm5m3m2_ca_w_2_400_s_0_360=8.23e-05 mcm5m3m2_cc_w_2_400_s_0_360=8.00e-11 mcm5m3m2_cf_w_2_400_s_0_360=1.47e-11
+  mcm5m3m2_ca_w_2_400_s_0_450=8.23e-05 mcm5m3m2_cc_w_2_400_s_0_450=7.03e-11 mcm5m3m2_cf_w_2_400_s_0_450=1.77e-11
+  mcm5m3m2_ca_w_2_400_s_0_600=8.23e-05 mcm5m3m2_cc_w_2_400_s_0_600=5.70e-11 mcm5m3m2_cf_w_2_400_s_0_600=2.23e-11
+  mcm5m3m2_ca_w_2_400_s_0_800=8.23e-05 mcm5m3m2_cc_w_2_400_s_0_800=4.39e-11 mcm5m3m2_cf_w_2_400_s_0_800=2.78e-11
+  mcm5m3m2_ca_w_2_400_s_1_000=8.23e-05 mcm5m3m2_cc_w_2_400_s_1_000=3.42e-11 mcm5m3m2_cf_w_2_400_s_1_000=3.25e-11
+  mcm5m3m2_ca_w_2_400_s_1_200=8.23e-05 mcm5m3m2_cc_w_2_400_s_1_200=2.69e-11 mcm5m3m2_cf_w_2_400_s_1_200=3.66e-11
+  mcm5m3m2_ca_w_2_400_s_2_100=8.23e-05 mcm5m3m2_cc_w_2_400_s_2_100=1.03e-11 mcm5m3m2_cf_w_2_400_s_2_100=4.86e-11
+  mcm5m3m2_ca_w_2_400_s_3_300=8.23e-05 mcm5m3m2_cc_w_2_400_s_3_300=3.17e-12 mcm5m3m2_cf_w_2_400_s_3_300=5.50e-11
+  mcm5m3m2_ca_w_2_400_s_9_000=8.23e-05 mcm5m3m2_cc_w_2_400_s_9_000=1.00e-14 mcm5m3m2_cf_w_2_400_s_9_000=5.80e-11
+  mcrdlm3f_ca_w_0_300_s_0_300=1.39e-05 mcrdlm3f_cc_w_0_300_s_0_300=9.49e-11 mcrdlm3f_cf_w_0_300_s_0_300=2.29e-12
+  mcrdlm3f_ca_w_0_300_s_0_360=1.39e-05 mcrdlm3f_cc_w_0_300_s_0_360=8.92e-11 mcrdlm3f_cf_w_0_300_s_0_360=2.70e-12
+  mcrdlm3f_ca_w_0_300_s_0_450=1.39e-05 mcrdlm3f_cc_w_0_300_s_0_450=8.10e-11 mcrdlm3f_cf_w_0_300_s_0_450=3.33e-12
+  mcrdlm3f_ca_w_0_300_s_0_600=1.39e-05 mcrdlm3f_cc_w_0_300_s_0_600=7.02e-11 mcrdlm3f_cf_w_0_300_s_0_600=4.36e-12
+  mcrdlm3f_ca_w_0_300_s_0_800=1.39e-05 mcrdlm3f_cc_w_0_300_s_0_800=5.99e-11 mcrdlm3f_cf_w_0_300_s_0_800=5.58e-12
+  mcrdlm3f_ca_w_0_300_s_1_000=1.39e-05 mcrdlm3f_cc_w_0_300_s_1_000=5.17e-11 mcrdlm3f_cf_w_0_300_s_1_000=6.84e-12
+  mcrdlm3f_ca_w_0_300_s_1_200=1.39e-05 mcrdlm3f_cc_w_0_300_s_1_200=4.55e-11 mcrdlm3f_cf_w_0_300_s_1_200=8.07e-12
+  mcrdlm3f_ca_w_0_300_s_2_100=1.39e-05 mcrdlm3f_cc_w_0_300_s_2_100=2.93e-11 mcrdlm3f_cf_w_0_300_s_2_100=1.33e-11
+  mcrdlm3f_ca_w_0_300_s_3_300=1.39e-05 mcrdlm3f_cc_w_0_300_s_3_300=1.91e-11 mcrdlm3f_cf_w_0_300_s_3_300=1.84e-11
+  mcrdlm3f_ca_w_0_300_s_9_000=1.39e-05 mcrdlm3f_cc_w_0_300_s_9_000=3.81e-12 mcrdlm3f_cf_w_0_300_s_9_000=2.99e-11
+  mcrdlm3f_ca_w_2_400_s_0_300=1.39e-05 mcrdlm3f_cc_w_2_400_s_0_300=1.18e-10 mcrdlm3f_cf_w_2_400_s_0_300=2.32e-12
+  mcrdlm3f_ca_w_2_400_s_0_360=1.39e-05 mcrdlm3f_cc_w_2_400_s_0_360=1.11e-10 mcrdlm3f_cf_w_2_400_s_0_360=2.73e-12
+  mcrdlm3f_ca_w_2_400_s_0_450=1.39e-05 mcrdlm3f_cc_w_2_400_s_0_450=1.02e-10 mcrdlm3f_cf_w_2_400_s_0_450=3.33e-12
+  mcrdlm3f_ca_w_2_400_s_0_600=1.39e-05 mcrdlm3f_cc_w_2_400_s_0_600=8.85e-11 mcrdlm3f_cf_w_2_400_s_0_600=4.33e-12
+  mcrdlm3f_ca_w_2_400_s_0_800=1.39e-05 mcrdlm3f_cc_w_2_400_s_0_800=7.55e-11 mcrdlm3f_cf_w_2_400_s_0_800=5.64e-12
+  mcrdlm3f_ca_w_2_400_s_1_000=1.39e-05 mcrdlm3f_cc_w_2_400_s_1_000=6.55e-11 mcrdlm3f_cf_w_2_400_s_1_000=6.92e-12
+  mcrdlm3f_ca_w_2_400_s_1_200=1.39e-05 mcrdlm3f_cc_w_2_400_s_1_200=5.79e-11 mcrdlm3f_cf_w_2_400_s_1_200=8.16e-12
+  mcrdlm3f_ca_w_2_400_s_2_100=1.39e-05 mcrdlm3f_cc_w_2_400_s_2_100=3.80e-11 mcrdlm3f_cf_w_2_400_s_2_100=1.33e-11
+  mcrdlm3f_ca_w_2_400_s_3_300=1.39e-05 mcrdlm3f_cc_w_2_400_s_3_300=2.50e-11 mcrdlm3f_cf_w_2_400_s_3_300=1.91e-11
+  mcrdlm3f_ca_w_2_400_s_9_000=1.39e-05 mcrdlm3f_cc_w_2_400_s_9_000=5.35e-12 mcrdlm3f_cf_w_2_400_s_9_000=3.30e-11
+  mcrdlm3d_ca_w_0_300_s_0_300=1.54e-05 mcrdlm3d_cc_w_0_300_s_0_300=9.47e-11 mcrdlm3d_cf_w_0_300_s_0_300=2.53e-12
+  mcrdlm3d_ca_w_0_300_s_0_360=1.54e-05 mcrdlm3d_cc_w_0_300_s_0_360=8.88e-11 mcrdlm3d_cf_w_0_300_s_0_360=2.98e-12
+  mcrdlm3d_ca_w_0_300_s_0_450=1.54e-05 mcrdlm3d_cc_w_0_300_s_0_450=8.06e-11 mcrdlm3d_cf_w_0_300_s_0_450=3.68e-12
+  mcrdlm3d_ca_w_0_300_s_0_600=1.54e-05 mcrdlm3d_cc_w_0_300_s_0_600=6.97e-11 mcrdlm3d_cf_w_0_300_s_0_600=4.80e-12
+  mcrdlm3d_ca_w_0_300_s_0_800=1.54e-05 mcrdlm3d_cc_w_0_300_s_0_800=5.93e-11 mcrdlm3d_cf_w_0_300_s_0_800=6.15e-12
+  mcrdlm3d_ca_w_0_300_s_1_000=1.54e-05 mcrdlm3d_cc_w_0_300_s_1_000=5.10e-11 mcrdlm3d_cf_w_0_300_s_1_000=7.52e-12
+  mcrdlm3d_ca_w_0_300_s_1_200=1.54e-05 mcrdlm3d_cc_w_0_300_s_1_200=4.47e-11 mcrdlm3d_cf_w_0_300_s_1_200=8.86e-12
+  mcrdlm3d_ca_w_0_300_s_2_100=1.54e-05 mcrdlm3d_cc_w_0_300_s_2_100=2.83e-11 mcrdlm3d_cf_w_0_300_s_2_100=1.45e-11
+  mcrdlm3d_ca_w_0_300_s_3_300=1.54e-05 mcrdlm3d_cc_w_0_300_s_3_300=1.82e-11 mcrdlm3d_cf_w_0_300_s_3_300=1.99e-11
+  mcrdlm3d_ca_w_0_300_s_9_000=1.54e-05 mcrdlm3d_cc_w_0_300_s_9_000=3.37e-12 mcrdlm3d_cf_w_0_300_s_9_000=3.13e-11
+  mcrdlm3d_ca_w_2_400_s_0_300=1.54e-05 mcrdlm3d_cc_w_2_400_s_0_300=1.17e-10 mcrdlm3d_cf_w_2_400_s_0_300=2.57e-12
+  mcrdlm3d_ca_w_2_400_s_0_360=1.54e-05 mcrdlm3d_cc_w_2_400_s_0_360=1.10e-10 mcrdlm3d_cf_w_2_400_s_0_360=3.02e-12
+  mcrdlm3d_ca_w_2_400_s_0_450=1.54e-05 mcrdlm3d_cc_w_2_400_s_0_450=1.01e-10 mcrdlm3d_cf_w_2_400_s_0_450=3.69e-12
+  mcrdlm3d_ca_w_2_400_s_0_600=1.54e-05 mcrdlm3d_cc_w_2_400_s_0_600=8.73e-11 mcrdlm3d_cf_w_2_400_s_0_600=4.78e-12
+  mcrdlm3d_ca_w_2_400_s_0_800=1.54e-05 mcrdlm3d_cc_w_2_400_s_0_800=7.42e-11 mcrdlm3d_cf_w_2_400_s_0_800=6.22e-12
+  mcrdlm3d_ca_w_2_400_s_1_000=1.54e-05 mcrdlm3d_cc_w_2_400_s_1_000=6.42e-11 mcrdlm3d_cf_w_2_400_s_1_000=7.61e-12
+  mcrdlm3d_ca_w_2_400_s_1_200=1.54e-05 mcrdlm3d_cc_w_2_400_s_1_200=5.66e-11 mcrdlm3d_cf_w_2_400_s_1_200=8.97e-12
+  mcrdlm3d_ca_w_2_400_s_2_100=1.54e-05 mcrdlm3d_cc_w_2_400_s_2_100=3.66e-11 mcrdlm3d_cf_w_2_400_s_2_100=1.45e-11
+  mcrdlm3d_ca_w_2_400_s_3_300=1.54e-05 mcrdlm3d_cc_w_2_400_s_3_300=2.38e-11 mcrdlm3d_cf_w_2_400_s_3_300=2.06e-11
+  mcrdlm3d_ca_w_2_400_s_9_000=1.54e-05 mcrdlm3d_cc_w_2_400_s_9_000=4.79e-12 mcrdlm3d_cf_w_2_400_s_9_000=3.46e-11
+  mcrdlm3p1_ca_w_0_300_s_0_300=1.65e-05 mcrdlm3p1_cc_w_0_300_s_0_300=9.44e-11 mcrdlm3p1_cf_w_0_300_s_0_300=2.72e-12
+  mcrdlm3p1_ca_w_0_300_s_0_360=1.65e-05 mcrdlm3p1_cc_w_0_300_s_0_360=8.84e-11 mcrdlm3p1_cf_w_0_300_s_0_360=3.20e-12
+  mcrdlm3p1_ca_w_0_300_s_0_450=1.65e-05 mcrdlm3p1_cc_w_0_300_s_0_450=8.02e-11 mcrdlm3p1_cf_w_0_300_s_0_450=3.94e-12
+  mcrdlm3p1_ca_w_0_300_s_0_600=1.65e-05 mcrdlm3p1_cc_w_0_300_s_0_600=6.93e-11 mcrdlm3p1_cf_w_0_300_s_0_600=5.15e-12
+  mcrdlm3p1_ca_w_0_300_s_0_800=1.65e-05 mcrdlm3p1_cc_w_0_300_s_0_800=5.87e-11 mcrdlm3p1_cf_w_0_300_s_0_800=6.58e-12
+  mcrdlm3p1_ca_w_0_300_s_1_000=1.65e-05 mcrdlm3p1_cc_w_0_300_s_1_000=5.05e-11 mcrdlm3p1_cf_w_0_300_s_1_000=8.06e-12
+  mcrdlm3p1_ca_w_0_300_s_1_200=1.65e-05 mcrdlm3p1_cc_w_0_300_s_1_200=4.42e-11 mcrdlm3p1_cf_w_0_300_s_1_200=9.47e-12
+  mcrdlm3p1_ca_w_0_300_s_2_100=1.65e-05 mcrdlm3p1_cc_w_0_300_s_2_100=2.76e-11 mcrdlm3p1_cf_w_0_300_s_2_100=1.54e-11
+  mcrdlm3p1_ca_w_0_300_s_3_300=1.65e-05 mcrdlm3p1_cc_w_0_300_s_3_300=1.75e-11 mcrdlm3p1_cf_w_0_300_s_3_300=2.10e-11
+  mcrdlm3p1_ca_w_0_300_s_9_000=1.65e-05 mcrdlm3p1_cc_w_0_300_s_9_000=3.09e-12 mcrdlm3p1_cf_w_0_300_s_9_000=3.23e-11
+  mcrdlm3p1_ca_w_2_400_s_0_300=1.65e-05 mcrdlm3p1_cc_w_2_400_s_0_300=1.16e-10 mcrdlm3p1_cf_w_2_400_s_0_300=2.79e-12
+  mcrdlm3p1_ca_w_2_400_s_0_360=1.65e-05 mcrdlm3p1_cc_w_2_400_s_0_360=1.09e-10 mcrdlm3p1_cf_w_2_400_s_0_360=3.26e-12
+  mcrdlm3p1_ca_w_2_400_s_0_450=1.65e-05 mcrdlm3p1_cc_w_2_400_s_0_450=9.97e-11 mcrdlm3p1_cf_w_2_400_s_0_450=3.98e-12
+  mcrdlm3p1_ca_w_2_400_s_0_600=1.65e-05 mcrdlm3p1_cc_w_2_400_s_0_600=8.64e-11 mcrdlm3p1_cf_w_2_400_s_0_600=5.15e-12
+  mcrdlm3p1_ca_w_2_400_s_0_800=1.65e-05 mcrdlm3p1_cc_w_2_400_s_0_800=7.33e-11 mcrdlm3p1_cf_w_2_400_s_0_800=6.68e-12
+  mcrdlm3p1_ca_w_2_400_s_1_000=1.65e-05 mcrdlm3p1_cc_w_2_400_s_1_000=6.33e-11 mcrdlm3p1_cf_w_2_400_s_1_000=8.17e-12
+  mcrdlm3p1_ca_w_2_400_s_1_200=1.65e-05 mcrdlm3p1_cc_w_2_400_s_1_200=5.57e-11 mcrdlm3p1_cf_w_2_400_s_1_200=9.61e-12
+  mcrdlm3p1_ca_w_2_400_s_2_100=1.65e-05 mcrdlm3p1_cc_w_2_400_s_2_100=3.57e-11 mcrdlm3p1_cf_w_2_400_s_2_100=1.55e-11
+  mcrdlm3p1_ca_w_2_400_s_3_300=1.65e-05 mcrdlm3p1_cc_w_2_400_s_3_300=2.29e-11 mcrdlm3p1_cf_w_2_400_s_3_300=2.18e-11
+  mcrdlm3p1_ca_w_2_400_s_9_000=1.65e-05 mcrdlm3p1_cc_w_2_400_s_9_000=4.43e-12 mcrdlm3p1_cf_w_2_400_s_9_000=3.57e-11
+  mcrdlm3l1_ca_w_0_300_s_0_300=2.04e-05 mcrdlm3l1_cc_w_0_300_s_0_300=9.34e-11 mcrdlm3l1_cf_w_0_300_s_0_300=3.33e-12
+  mcrdlm3l1_ca_w_0_300_s_0_360=2.04e-05 mcrdlm3l1_cc_w_0_300_s_0_360=8.75e-11 mcrdlm3l1_cf_w_0_300_s_0_360=3.92e-12
+  mcrdlm3l1_ca_w_0_300_s_0_450=2.04e-05 mcrdlm3l1_cc_w_0_300_s_0_450=7.91e-11 mcrdlm3l1_cf_w_0_300_s_0_450=4.82e-12
+  mcrdlm3l1_ca_w_0_300_s_0_600=2.04e-05 mcrdlm3l1_cc_w_0_300_s_0_600=6.81e-11 mcrdlm3l1_cf_w_0_300_s_0_600=6.27e-12
+  mcrdlm3l1_ca_w_0_300_s_0_800=2.04e-05 mcrdlm3l1_cc_w_0_300_s_0_800=5.73e-11 mcrdlm3l1_cf_w_0_300_s_0_800=8.01e-12
+  mcrdlm3l1_ca_w_0_300_s_1_000=2.04e-05 mcrdlm3l1_cc_w_0_300_s_1_000=4.88e-11 mcrdlm3l1_cf_w_0_300_s_1_000=9.73e-12
+  mcrdlm3l1_ca_w_0_300_s_1_200=2.04e-05 mcrdlm3l1_cc_w_0_300_s_1_200=4.24e-11 mcrdlm3l1_cf_w_0_300_s_1_200=1.14e-11
+  mcrdlm3l1_ca_w_0_300_s_2_100=2.04e-05 mcrdlm3l1_cc_w_0_300_s_2_100=2.57e-11 mcrdlm3l1_cf_w_0_300_s_2_100=1.82e-11
+  mcrdlm3l1_ca_w_0_300_s_3_300=2.04e-05 mcrdlm3l1_cc_w_0_300_s_3_300=1.56e-11 mcrdlm3l1_cf_w_0_300_s_3_300=2.43e-11
+  mcrdlm3l1_ca_w_0_300_s_9_000=2.04e-05 mcrdlm3l1_cc_w_0_300_s_9_000=2.42e-12 mcrdlm3l1_cf_w_0_300_s_9_000=3.52e-11
+  mcrdlm3l1_ca_w_2_400_s_0_300=2.04e-05 mcrdlm3l1_cc_w_2_400_s_0_300=1.14e-10 mcrdlm3l1_cf_w_2_400_s_0_300=3.37e-12
+  mcrdlm3l1_ca_w_2_400_s_0_360=2.04e-05 mcrdlm3l1_cc_w_2_400_s_0_360=1.06e-10 mcrdlm3l1_cf_w_2_400_s_0_360=3.96e-12
+  mcrdlm3l1_ca_w_2_400_s_0_450=2.04e-05 mcrdlm3l1_cc_w_2_400_s_0_450=9.68e-11 mcrdlm3l1_cf_w_2_400_s_0_450=4.83e-12
+  mcrdlm3l1_ca_w_2_400_s_0_600=2.04e-05 mcrdlm3l1_cc_w_2_400_s_0_600=8.37e-11 mcrdlm3l1_cf_w_2_400_s_0_600=6.24e-12
+  mcrdlm3l1_ca_w_2_400_s_0_800=2.04e-05 mcrdlm3l1_cc_w_2_400_s_0_800=7.06e-11 mcrdlm3l1_cf_w_2_400_s_0_800=8.09e-12
+  mcrdlm3l1_ca_w_2_400_s_1_000=2.04e-05 mcrdlm3l1_cc_w_2_400_s_1_000=6.06e-11 mcrdlm3l1_cf_w_2_400_s_1_000=9.87e-12
+  mcrdlm3l1_ca_w_2_400_s_1_200=2.04e-05 mcrdlm3l1_cc_w_2_400_s_1_200=5.31e-11 mcrdlm3l1_cf_w_2_400_s_1_200=1.16e-11
+  mcrdlm3l1_ca_w_2_400_s_2_100=2.04e-05 mcrdlm3l1_cc_w_2_400_s_2_100=3.33e-11 mcrdlm3l1_cf_w_2_400_s_2_100=1.84e-11
+  mcrdlm3l1_ca_w_2_400_s_3_300=2.04e-05 mcrdlm3l1_cc_w_2_400_s_3_300=2.07e-11 mcrdlm3l1_cf_w_2_400_s_3_300=2.53e-11
+  mcrdlm3l1_ca_w_2_400_s_9_000=2.04e-05 mcrdlm3l1_cc_w_2_400_s_9_000=3.61e-12 mcrdlm3l1_cf_w_2_400_s_9_000=3.89e-11
+  mcrdlm3m1_ca_w_0_300_s_0_300=3.06e-05 mcrdlm3m1_cc_w_0_300_s_0_300=9.11e-11 mcrdlm3m1_cf_w_0_300_s_0_300=4.91e-12
+  mcrdlm3m1_ca_w_0_300_s_0_360=3.06e-05 mcrdlm3m1_cc_w_0_300_s_0_360=8.50e-11 mcrdlm3m1_cf_w_0_300_s_0_360=5.76e-12
+  mcrdlm3m1_ca_w_0_300_s_0_450=3.06e-05 mcrdlm3m1_cc_w_0_300_s_0_450=7.64e-11 mcrdlm3m1_cf_w_0_300_s_0_450=7.03e-12
+  mcrdlm3m1_ca_w_0_300_s_0_600=3.06e-05 mcrdlm3m1_cc_w_0_300_s_0_600=6.50e-11 mcrdlm3m1_cf_w_0_300_s_0_600=9.08e-12
+  mcrdlm3m1_ca_w_0_300_s_0_800=3.06e-05 mcrdlm3m1_cc_w_0_300_s_0_800=5.39e-11 mcrdlm3m1_cf_w_0_300_s_0_800=1.15e-11
+  mcrdlm3m1_ca_w_0_300_s_1_000=3.06e-05 mcrdlm3m1_cc_w_0_300_s_1_000=4.53e-11 mcrdlm3m1_cf_w_0_300_s_1_000=1.39e-11
+  mcrdlm3m1_ca_w_0_300_s_1_200=3.06e-05 mcrdlm3m1_cc_w_0_300_s_1_200=3.87e-11 mcrdlm3m1_cf_w_0_300_s_1_200=1.61e-11
+  mcrdlm3m1_ca_w_0_300_s_2_100=3.06e-05 mcrdlm3m1_cc_w_0_300_s_2_100=2.18e-11 mcrdlm3m1_cf_w_0_300_s_2_100=2.46e-11
+  mcrdlm3m1_ca_w_0_300_s_3_300=3.06e-05 mcrdlm3m1_cc_w_0_300_s_3_300=1.23e-11 mcrdlm3m1_cf_w_0_300_s_3_300=3.13e-11
+  mcrdlm3m1_ca_w_0_300_s_9_000=3.06e-05 mcrdlm3m1_cc_w_0_300_s_9_000=1.59e-12 mcrdlm3m1_cf_w_0_300_s_9_000=4.09e-11
+  mcrdlm3m1_ca_w_2_400_s_0_300=3.06e-05 mcrdlm3m1_cc_w_2_400_s_0_300=1.09e-10 mcrdlm3m1_cf_w_2_400_s_0_300=4.94e-12
+  mcrdlm3m1_ca_w_2_400_s_0_360=3.06e-05 mcrdlm3m1_cc_w_2_400_s_0_360=1.02e-10 mcrdlm3m1_cf_w_2_400_s_0_360=5.78e-12
+  mcrdlm3m1_ca_w_2_400_s_0_450=3.06e-05 mcrdlm3m1_cc_w_2_400_s_0_450=9.19e-11 mcrdlm3m1_cf_w_2_400_s_0_450=7.04e-12
+  mcrdlm3m1_ca_w_2_400_s_0_600=3.06e-05 mcrdlm3m1_cc_w_2_400_s_0_600=7.88e-11 mcrdlm3m1_cf_w_2_400_s_0_600=9.05e-12
+  mcrdlm3m1_ca_w_2_400_s_0_800=3.06e-05 mcrdlm3m1_cc_w_2_400_s_0_800=6.57e-11 mcrdlm3m1_cf_w_2_400_s_0_800=1.16e-11
+  mcrdlm3m1_ca_w_2_400_s_1_000=3.06e-05 mcrdlm3m1_cc_w_2_400_s_1_000=5.58e-11 mcrdlm3m1_cf_w_2_400_s_1_000=1.41e-11
+  mcrdlm3m1_ca_w_2_400_s_1_200=3.06e-05 mcrdlm3m1_cc_w_2_400_s_1_200=4.82e-11 mcrdlm3m1_cf_w_2_400_s_1_200=1.63e-11
+  mcrdlm3m1_ca_w_2_400_s_2_100=3.06e-05 mcrdlm3m1_cc_w_2_400_s_2_100=2.88e-11 mcrdlm3m1_cf_w_2_400_s_2_100=2.48e-11
+  mcrdlm3m1_ca_w_2_400_s_3_300=3.06e-05 mcrdlm3m1_cc_w_2_400_s_3_300=1.70e-11 mcrdlm3m1_cf_w_2_400_s_3_300=3.26e-11
+  mcrdlm3m1_ca_w_2_400_s_9_000=3.06e-05 mcrdlm3m1_cc_w_2_400_s_9_000=2.50e-12 mcrdlm3m1_cf_w_2_400_s_9_000=4.49e-11
+  mcrdlm3m2_ca_w_0_300_s_0_300=6.79e-05 mcrdlm3m2_cc_w_0_300_s_0_300=8.45e-11 mcrdlm3m2_cf_w_0_300_s_0_300=1.03e-11
+  mcrdlm3m2_ca_w_0_300_s_0_360=6.79e-05 mcrdlm3m2_cc_w_0_300_s_0_360=7.77e-11 mcrdlm3m2_cf_w_0_300_s_0_360=1.20e-11
+  mcrdlm3m2_ca_w_0_300_s_0_450=6.79e-05 mcrdlm3m2_cc_w_0_300_s_0_450=6.93e-11 mcrdlm3m2_cf_w_0_300_s_0_450=1.44e-11
+  mcrdlm3m2_ca_w_0_300_s_0_600=6.79e-05 mcrdlm3m2_cc_w_0_300_s_0_600=5.76e-11 mcrdlm3m2_cf_w_0_300_s_0_600=1.81e-11
+  mcrdlm3m2_ca_w_0_300_s_0_800=6.79e-05 mcrdlm3m2_cc_w_0_300_s_0_800=4.63e-11 mcrdlm3m2_cf_w_0_300_s_0_800=2.24e-11
+  mcrdlm3m2_ca_w_0_300_s_1_000=6.79e-05 mcrdlm3m2_cc_w_0_300_s_1_000=3.78e-11 mcrdlm3m2_cf_w_0_300_s_1_000=2.62e-11
+  mcrdlm3m2_ca_w_0_300_s_1_200=6.79e-05 mcrdlm3m2_cc_w_0_300_s_1_200=3.14e-11 mcrdlm3m2_cf_w_0_300_s_1_200=2.94e-11
+  mcrdlm3m2_ca_w_0_300_s_2_100=6.79e-05 mcrdlm3m2_cc_w_0_300_s_2_100=1.55e-11 mcrdlm3m2_cf_w_0_300_s_2_100=4.01e-11
+  mcrdlm3m2_ca_w_0_300_s_3_300=6.79e-05 mcrdlm3m2_cc_w_0_300_s_3_300=7.93e-12 mcrdlm3m2_cf_w_0_300_s_3_300=4.65e-11
+  mcrdlm3m2_ca_w_0_300_s_9_000=6.79e-05 mcrdlm3m2_cc_w_0_300_s_9_000=8.39e-13 mcrdlm3m2_cf_w_0_300_s_9_000=5.32e-11
+  mcrdlm3m2_ca_w_2_400_s_0_300=6.79e-05 mcrdlm3m2_cc_w_2_400_s_0_300=9.92e-11 mcrdlm3m2_cf_w_2_400_s_0_300=1.04e-11
+  mcrdlm3m2_ca_w_2_400_s_0_360=6.79e-05 mcrdlm3m2_cc_w_2_400_s_0_360=9.22e-11 mcrdlm3m2_cf_w_2_400_s_0_360=1.20e-11
+  mcrdlm3m2_ca_w_2_400_s_0_450=6.79e-05 mcrdlm3m2_cc_w_2_400_s_0_450=8.28e-11 mcrdlm3m2_cf_w_2_400_s_0_450=1.44e-11
+  mcrdlm3m2_ca_w_2_400_s_0_600=6.79e-05 mcrdlm3m2_cc_w_2_400_s_0_600=6.99e-11 mcrdlm3m2_cf_w_2_400_s_0_600=1.81e-11
+  mcrdlm3m2_ca_w_2_400_s_0_800=6.79e-05 mcrdlm3m2_cc_w_2_400_s_0_800=5.70e-11 mcrdlm3m2_cf_w_2_400_s_0_800=2.24e-11
+  mcrdlm3m2_ca_w_2_400_s_1_000=6.79e-05 mcrdlm3m2_cc_w_2_400_s_1_000=4.75e-11 mcrdlm3m2_cf_w_2_400_s_1_000=2.63e-11
+  mcrdlm3m2_ca_w_2_400_s_1_200=6.79e-05 mcrdlm3m2_cc_w_2_400_s_1_200=4.01e-11 mcrdlm3m2_cf_w_2_400_s_1_200=2.96e-11
+  mcrdlm3m2_ca_w_2_400_s_2_100=6.79e-05 mcrdlm3m2_cc_w_2_400_s_2_100=2.24e-11 mcrdlm3m2_cf_w_2_400_s_2_100=4.04e-11
+  mcrdlm3m2_ca_w_2_400_s_3_300=6.79e-05 mcrdlm3m2_cc_w_2_400_s_3_300=1.23e-11 mcrdlm3m2_cf_w_2_400_s_3_300=4.84e-11
+  mcrdlm3m2_ca_w_2_400_s_9_000=6.79e-05 mcrdlm3m2_cc_w_2_400_s_9_000=1.55e-12 mcrdlm3m2_cf_w_2_400_s_9_000=5.83e-11
+  mcm5m4f_ca_w_0_300_s_0_300=6.06e-05 mcm5m4f_cc_w_0_300_s_0_300=8.52e-11 mcm5m4f_cf_w_0_300_s_0_300=8.98e-12
+  mcm5m4f_ca_w_0_300_s_0_360=6.06e-05 mcm5m4f_cc_w_0_300_s_0_360=7.87e-11 mcm5m4f_cf_w_0_300_s_0_360=1.05e-11
+  mcm5m4f_ca_w_0_300_s_0_450=6.06e-05 mcm5m4f_cc_w_0_300_s_0_450=7.01e-11 mcm5m4f_cf_w_0_300_s_0_450=1.27e-11
+  mcm5m4f_ca_w_0_300_s_0_600=6.06e-05 mcm5m4f_cc_w_0_300_s_0_600=5.82e-11 mcm5m4f_cf_w_0_300_s_0_600=1.62e-11
+  mcm5m4f_ca_w_0_300_s_0_800=6.06e-05 mcm5m4f_cc_w_0_300_s_0_800=4.64e-11 mcm5m4f_cf_w_0_300_s_0_800=2.04e-11
+  mcm5m4f_ca_w_0_300_s_1_000=6.06e-05 mcm5m4f_cc_w_0_300_s_1_000=3.77e-11 mcm5m4f_cf_w_0_300_s_1_000=2.41e-11
+  mcm5m4f_ca_w_0_300_s_1_200=6.06e-05 mcm5m4f_cc_w_0_300_s_1_200=3.08e-11 mcm5m4f_cf_w_0_300_s_1_200=2.74e-11
+  mcm5m4f_ca_w_0_300_s_2_100=6.06e-05 mcm5m4f_cc_w_0_300_s_2_100=1.44e-11 mcm5m4f_cf_w_0_300_s_2_100=3.80e-11
+  mcm5m4f_ca_w_0_300_s_3_300=6.06e-05 mcm5m4f_cc_w_0_300_s_3_300=6.29e-12 mcm5m4f_cf_w_0_300_s_3_300=4.48e-11
+  mcm5m4f_ca_w_0_300_s_9_000=6.06e-05 mcm5m4f_cc_w_0_300_s_9_000=2.95e-13 mcm5m4f_cf_w_0_300_s_9_000=5.04e-11
+  mcm5m4f_ca_w_2_400_s_0_300=6.06e-05 mcm5m4f_cc_w_2_400_s_0_300=9.70e-11 mcm5m4f_cf_w_2_400_s_0_300=9.06e-12
+  mcm5m4f_ca_w_2_400_s_0_360=6.06e-05 mcm5m4f_cc_w_2_400_s_0_360=8.97e-11 mcm5m4f_cf_w_2_400_s_0_360=1.06e-11
+  mcm5m4f_ca_w_2_400_s_0_450=6.06e-05 mcm5m4f_cc_w_2_400_s_0_450=8.00e-11 mcm5m4f_cf_w_2_400_s_0_450=1.28e-11
+  mcm5m4f_ca_w_2_400_s_0_600=6.06e-05 mcm5m4f_cc_w_2_400_s_0_600=6.70e-11 mcm5m4f_cf_w_2_400_s_0_600=1.63e-11
+  mcm5m4f_ca_w_2_400_s_0_800=6.06e-05 mcm5m4f_cc_w_2_400_s_0_800=5.37e-11 mcm5m4f_cf_w_2_400_s_0_800=2.06e-11
+  mcm5m4f_ca_w_2_400_s_1_000=6.06e-05 mcm5m4f_cc_w_2_400_s_1_000=4.38e-11 mcm5m4f_cf_w_2_400_s_1_000=2.44e-11
+  mcm5m4f_ca_w_2_400_s_1_200=6.06e-05 mcm5m4f_cc_w_2_400_s_1_200=3.64e-11 mcm5m4f_cf_w_2_400_s_1_200=2.77e-11
+  mcm5m4f_ca_w_2_400_s_2_100=6.06e-05 mcm5m4f_cc_w_2_400_s_2_100=1.81e-11 mcm5m4f_cf_w_2_400_s_2_100=3.87e-11
+  mcm5m4f_ca_w_2_400_s_3_300=6.06e-05 mcm5m4f_cc_w_2_400_s_3_300=8.37e-12 mcm5m4f_cf_w_2_400_s_3_300=4.65e-11
+  mcm5m4f_ca_w_2_400_s_9_000=6.06e-05 mcm5m4f_cc_w_2_400_s_9_000=3.65e-13 mcm5m4f_cf_w_2_400_s_9_000=5.40e-11
+  mcm5m4d_ca_w_0_300_s_0_300=6.13e-05 mcm5m4d_cc_w_0_300_s_0_300=8.51e-11 mcm5m4d_cf_w_0_300_s_0_300=9.09e-12
+  mcm5m4d_ca_w_0_300_s_0_360=6.13e-05 mcm5m4d_cc_w_0_300_s_0_360=7.85e-11 mcm5m4d_cf_w_0_300_s_0_360=1.06e-11
+  mcm5m4d_ca_w_0_300_s_0_450=6.13e-05 mcm5m4d_cc_w_0_300_s_0_450=6.99e-11 mcm5m4d_cf_w_0_300_s_0_450=1.29e-11
+  mcm5m4d_ca_w_0_300_s_0_600=6.13e-05 mcm5m4d_cc_w_0_300_s_0_600=5.79e-11 mcm5m4d_cf_w_0_300_s_0_600=1.65e-11
+  mcm5m4d_ca_w_0_300_s_0_800=6.13e-05 mcm5m4d_cc_w_0_300_s_0_800=4.60e-11 mcm5m4d_cf_w_0_300_s_0_800=2.06e-11
+  mcm5m4d_ca_w_0_300_s_1_000=6.13e-05 mcm5m4d_cc_w_0_300_s_1_000=3.73e-11 mcm5m4d_cf_w_0_300_s_1_000=2.44e-11
+  mcm5m4d_ca_w_0_300_s_1_200=6.13e-05 mcm5m4d_cc_w_0_300_s_1_200=3.05e-11 mcm5m4d_cf_w_0_300_s_1_200=2.78e-11
+  mcm5m4d_ca_w_0_300_s_2_100=6.13e-05 mcm5m4d_cc_w_0_300_s_2_100=1.40e-11 mcm5m4d_cf_w_0_300_s_2_100=3.84e-11
+  mcm5m4d_ca_w_0_300_s_3_300=6.13e-05 mcm5m4d_cc_w_0_300_s_3_300=5.99e-12 mcm5m4d_cf_w_0_300_s_3_300=4.52e-11
+  mcm5m4d_ca_w_0_300_s_9_000=6.13e-05 mcm5m4d_cc_w_0_300_s_9_000=2.30e-13 mcm5m4d_cf_w_0_300_s_9_000=5.05e-11
+  mcm5m4d_ca_w_2_400_s_0_300=6.13e-05 mcm5m4d_cc_w_2_400_s_0_300=9.63e-11 mcm5m4d_cf_w_2_400_s_0_300=9.18e-12
+  mcm5m4d_ca_w_2_400_s_0_360=6.13e-05 mcm5m4d_cc_w_2_400_s_0_360=8.91e-11 mcm5m4d_cf_w_2_400_s_0_360=1.07e-11
+  mcm5m4d_ca_w_2_400_s_0_450=6.13e-05 mcm5m4d_cc_w_2_400_s_0_450=7.93e-11 mcm5m4d_cf_w_2_400_s_0_450=1.30e-11
+  mcm5m4d_ca_w_2_400_s_0_600=6.13e-05 mcm5m4d_cc_w_2_400_s_0_600=6.62e-11 mcm5m4d_cf_w_2_400_s_0_600=1.65e-11
+  mcm5m4d_ca_w_2_400_s_0_800=6.13e-05 mcm5m4d_cc_w_2_400_s_0_800=5.29e-11 mcm5m4d_cf_w_2_400_s_0_800=2.08e-11
+  mcm5m4d_ca_w_2_400_s_1_000=6.13e-05 mcm5m4d_cc_w_2_400_s_1_000=4.32e-11 mcm5m4d_cf_w_2_400_s_1_000=2.47e-11
+  mcm5m4d_ca_w_2_400_s_1_200=6.13e-05 mcm5m4d_cc_w_2_400_s_1_200=3.56e-11 mcm5m4d_cf_w_2_400_s_1_200=2.81e-11
+  mcm5m4d_ca_w_2_400_s_2_100=6.13e-05 mcm5m4d_cc_w_2_400_s_2_100=1.74e-11 mcm5m4d_cf_w_2_400_s_2_100=3.92e-11
+  mcm5m4d_ca_w_2_400_s_3_300=6.13e-05 mcm5m4d_cc_w_2_400_s_3_300=7.79e-12 mcm5m4d_cf_w_2_400_s_3_300=4.69e-11
+  mcm5m4d_ca_w_2_400_s_9_000=6.13e-05 mcm5m4d_cc_w_2_400_s_9_000=3.15e-13 mcm5m4d_cf_w_2_400_s_9_000=5.40e-11
+  mcm5m4p1_ca_w_0_300_s_0_300=6.19e-05 mcm5m4p1_cc_w_0_300_s_0_300=8.49e-11 mcm5m4p1_cf_w_0_300_s_0_300=9.18e-12
+  mcm5m4p1_ca_w_0_300_s_0_360=6.19e-05 mcm5m4p1_cc_w_0_300_s_0_360=7.84e-11 mcm5m4p1_cf_w_0_300_s_0_360=1.07e-11
+  mcm5m4p1_ca_w_0_300_s_0_450=6.19e-05 mcm5m4p1_cc_w_0_300_s_0_450=6.97e-11 mcm5m4p1_cf_w_0_300_s_0_450=1.30e-11
+  mcm5m4p1_ca_w_0_300_s_0_600=6.19e-05 mcm5m4p1_cc_w_0_300_s_0_600=5.77e-11 mcm5m4p1_cf_w_0_300_s_0_600=1.66e-11
+  mcm5m4p1_ca_w_0_300_s_0_800=6.19e-05 mcm5m4p1_cc_w_0_300_s_0_800=4.58e-11 mcm5m4p1_cf_w_0_300_s_0_800=2.08e-11
+  mcm5m4p1_ca_w_0_300_s_1_000=6.19e-05 mcm5m4p1_cc_w_0_300_s_1_000=3.71e-11 mcm5m4p1_cf_w_0_300_s_1_000=2.47e-11
+  mcm5m4p1_ca_w_0_300_s_1_200=6.19e-05 mcm5m4p1_cc_w_0_300_s_1_200=3.02e-11 mcm5m4p1_cf_w_0_300_s_1_200=2.80e-11
+  mcm5m4p1_ca_w_0_300_s_2_100=6.19e-05 mcm5m4p1_cc_w_0_300_s_2_100=1.38e-11 mcm5m4p1_cf_w_0_300_s_2_100=3.87e-11
+  mcm5m4p1_ca_w_0_300_s_3_300=6.19e-05 mcm5m4p1_cc_w_0_300_s_3_300=5.74e-12 mcm5m4p1_cf_w_0_300_s_3_300=4.55e-11
+  mcm5m4p1_ca_w_0_300_s_9_000=6.19e-05 mcm5m4p1_cc_w_0_300_s_9_000=1.95e-13 mcm5m4p1_cf_w_0_300_s_9_000=5.07e-11
+  mcm5m4p1_ca_w_2_400_s_0_300=6.19e-05 mcm5m4p1_cc_w_2_400_s_0_300=9.58e-11 mcm5m4p1_cf_w_2_400_s_0_300=9.27e-12
+  mcm5m4p1_ca_w_2_400_s_0_360=6.19e-05 mcm5m4p1_cc_w_2_400_s_0_360=8.85e-11 mcm5m4p1_cf_w_2_400_s_0_360=1.08e-11
+  mcm5m4p1_ca_w_2_400_s_0_450=6.19e-05 mcm5m4p1_cc_w_2_400_s_0_450=7.89e-11 mcm5m4p1_cf_w_2_400_s_0_450=1.31e-11
+  mcm5m4p1_ca_w_2_400_s_0_600=6.19e-05 mcm5m4p1_cc_w_2_400_s_0_600=6.58e-11 mcm5m4p1_cf_w_2_400_s_0_600=1.67e-11
+  mcm5m4p1_ca_w_2_400_s_0_800=6.19e-05 mcm5m4p1_cc_w_2_400_s_0_800=5.24e-11 mcm5m4p1_cf_w_2_400_s_0_800=2.10e-11
+  mcm5m4p1_ca_w_2_400_s_1_000=6.19e-05 mcm5m4p1_cc_w_2_400_s_1_000=4.26e-11 mcm5m4p1_cf_w_2_400_s_1_000=2.49e-11
+  mcm5m4p1_ca_w_2_400_s_1_200=6.19e-05 mcm5m4p1_cc_w_2_400_s_1_200=3.51e-11 mcm5m4p1_cf_w_2_400_s_1_200=2.83e-11
+  mcm5m4p1_ca_w_2_400_s_2_100=6.19e-05 mcm5m4p1_cc_w_2_400_s_2_100=1.69e-11 mcm5m4p1_cf_w_2_400_s_2_100=3.95e-11
+  mcm5m4p1_ca_w_2_400_s_3_300=6.19e-05 mcm5m4p1_cc_w_2_400_s_3_300=7.41e-12 mcm5m4p1_cf_w_2_400_s_3_300=4.72e-11
+  mcm5m4p1_ca_w_2_400_s_9_000=6.19e-05 mcm5m4p1_cc_w_2_400_s_9_000=2.55e-13 mcm5m4p1_cf_w_2_400_s_9_000=5.40e-11
+  mcm5m4l1_ca_w_0_300_s_0_300=6.34e-05 mcm5m4l1_cc_w_0_300_s_0_300=8.46e-11 mcm5m4l1_cf_w_0_300_s_0_300=9.42e-12
+  mcm5m4l1_ca_w_0_300_s_0_360=6.34e-05 mcm5m4l1_cc_w_0_300_s_0_360=7.80e-11 mcm5m4l1_cf_w_0_300_s_0_360=1.10e-11
+  mcm5m4l1_ca_w_0_300_s_0_450=6.34e-05 mcm5m4l1_cc_w_0_300_s_0_450=6.93e-11 mcm5m4l1_cf_w_0_300_s_0_450=1.34e-11
+  mcm5m4l1_ca_w_0_300_s_0_600=6.34e-05 mcm5m4l1_cc_w_0_300_s_0_600=5.72e-11 mcm5m4l1_cf_w_0_300_s_0_600=1.71e-11
+  mcm5m4l1_ca_w_0_300_s_0_800=6.34e-05 mcm5m4l1_cc_w_0_300_s_0_800=4.52e-11 mcm5m4l1_cf_w_0_300_s_0_800=2.14e-11
+  mcm5m4l1_ca_w_0_300_s_1_000=6.34e-05 mcm5m4l1_cc_w_0_300_s_1_000=3.63e-11 mcm5m4l1_cf_w_0_300_s_1_000=2.53e-11
+  mcm5m4l1_ca_w_0_300_s_1_200=6.34e-05 mcm5m4l1_cc_w_0_300_s_1_200=2.95e-11 mcm5m4l1_cf_w_0_300_s_1_200=2.88e-11
+  mcm5m4l1_ca_w_0_300_s_2_100=6.34e-05 mcm5m4l1_cc_w_0_300_s_2_100=1.30e-11 mcm5m4l1_cf_w_0_300_s_2_100=3.96e-11
+  mcm5m4l1_ca_w_0_300_s_3_300=6.34e-05 mcm5m4l1_cc_w_0_300_s_3_300=5.16e-12 mcm5m4l1_cf_w_0_300_s_3_300=4.63e-11
+  mcm5m4l1_ca_w_0_300_s_9_000=6.34e-05 mcm5m4l1_cc_w_0_300_s_9_000=1.50e-13 mcm5m4l1_cf_w_0_300_s_9_000=5.11e-11
+  mcm5m4l1_ca_w_2_400_s_0_300=6.34e-05 mcm5m4l1_cc_w_2_400_s_0_300=9.45e-11 mcm5m4l1_cf_w_2_400_s_0_300=9.51e-12
+  mcm5m4l1_ca_w_2_400_s_0_360=6.34e-05 mcm5m4l1_cc_w_2_400_s_0_360=8.72e-11 mcm5m4l1_cf_w_2_400_s_0_360=1.11e-11
+  mcm5m4l1_ca_w_2_400_s_0_450=6.34e-05 mcm5m4l1_cc_w_2_400_s_0_450=7.75e-11 mcm5m4l1_cf_w_2_400_s_0_450=1.34e-11
+  mcm5m4l1_ca_w_2_400_s_0_600=6.34e-05 mcm5m4l1_cc_w_2_400_s_0_600=6.44e-11 mcm5m4l1_cf_w_2_400_s_0_600=1.71e-11
+  mcm5m4l1_ca_w_2_400_s_0_800=6.34e-05 mcm5m4l1_cc_w_2_400_s_0_800=5.11e-11 mcm5m4l1_cf_w_2_400_s_0_800=2.16e-11
+  mcm5m4l1_ca_w_2_400_s_1_000=6.34e-05 mcm5m4l1_cc_w_2_400_s_1_000=4.12e-11 mcm5m4l1_cf_w_2_400_s_1_000=2.56e-11
+  mcm5m4l1_ca_w_2_400_s_1_200=6.34e-05 mcm5m4l1_cc_w_2_400_s_1_200=3.37e-11 mcm5m4l1_cf_w_2_400_s_1_200=2.91e-11
+  mcm5m4l1_ca_w_2_400_s_2_100=6.34e-05 mcm5m4l1_cc_w_2_400_s_2_100=1.57e-11 mcm5m4l1_cf_w_2_400_s_2_100=4.04e-11
+  mcm5m4l1_ca_w_2_400_s_3_300=6.34e-05 mcm5m4l1_cc_w_2_400_s_3_300=6.47e-12 mcm5m4l1_cf_w_2_400_s_3_300=4.80e-11
+  mcm5m4l1_ca_w_2_400_s_9_000=6.34e-05 mcm5m4l1_cc_w_2_400_s_9_000=1.85e-13 mcm5m4l1_cf_w_2_400_s_9_000=5.40e-11
+  mcm5m4m1_ca_w_0_300_s_0_300=6.64e-05 mcm5m4m1_cc_w_0_300_s_0_300=8.38e-11 mcm5m4m1_cf_w_0_300_s_0_300=9.90e-12
+  mcm5m4m1_ca_w_0_300_s_0_360=6.64e-05 mcm5m4m1_cc_w_0_300_s_0_360=7.72e-11 mcm5m4m1_cf_w_0_300_s_0_360=1.16e-11
+  mcm5m4m1_ca_w_0_300_s_0_450=6.64e-05 mcm5m4m1_cc_w_0_300_s_0_450=6.84e-11 mcm5m4m1_cf_w_0_300_s_0_450=1.40e-11
+  mcm5m4m1_ca_w_0_300_s_0_600=6.64e-05 mcm5m4m1_cc_w_0_300_s_0_600=5.63e-11 mcm5m4m1_cf_w_0_300_s_0_600=1.79e-11
+  mcm5m4m1_ca_w_0_300_s_0_800=6.64e-05 mcm5m4m1_cc_w_0_300_s_0_800=4.41e-11 mcm5m4m1_cf_w_0_300_s_0_800=2.25e-11
+  mcm5m4m1_ca_w_0_300_s_1_000=6.64e-05 mcm5m4m1_cc_w_0_300_s_1_000=3.50e-11 mcm5m4m1_cf_w_0_300_s_1_000=2.66e-11
+  mcm5m4m1_ca_w_0_300_s_1_200=6.64e-05 mcm5m4m1_cc_w_0_300_s_1_200=2.81e-11 mcm5m4m1_cf_w_0_300_s_1_200=3.02e-11
+  mcm5m4m1_ca_w_0_300_s_2_100=6.64e-05 mcm5m4m1_cc_w_0_300_s_2_100=1.18e-11 mcm5m4m1_cf_w_0_300_s_2_100=4.12e-11
+  mcm5m4m1_ca_w_0_300_s_3_300=6.64e-05 mcm5m4m1_cc_w_0_300_s_3_300=4.23e-12 mcm5m4m1_cf_w_0_300_s_3_300=4.78e-11
+  mcm5m4m1_ca_w_0_300_s_9_000=6.64e-05 mcm5m4m1_cc_w_0_300_s_9_000=8.00e-14 mcm5m4m1_cf_w_0_300_s_9_000=5.17e-11
+  mcm5m4m1_ca_w_2_400_s_0_300=6.64e-05 mcm5m4m1_cc_w_2_400_s_0_300=9.21e-11 mcm5m4m1_cf_w_2_400_s_0_300=9.98e-12
+  mcm5m4m1_ca_w_2_400_s_0_360=6.64e-05 mcm5m4m1_cc_w_2_400_s_0_360=8.49e-11 mcm5m4m1_cf_w_2_400_s_0_360=1.17e-11
+  mcm5m4m1_ca_w_2_400_s_0_450=6.64e-05 mcm5m4m1_cc_w_2_400_s_0_450=7.52e-11 mcm5m4m1_cf_w_2_400_s_0_450=1.41e-11
+  mcm5m4m1_ca_w_2_400_s_0_600=6.64e-05 mcm5m4m1_cc_w_2_400_s_0_600=6.20e-11 mcm5m4m1_cf_w_2_400_s_0_600=1.80e-11
+  mcm5m4m1_ca_w_2_400_s_0_800=6.64e-05 mcm5m4m1_cc_w_2_400_s_0_800=4.87e-11 mcm5m4m1_cf_w_2_400_s_0_800=2.27e-11
+  mcm5m4m1_ca_w_2_400_s_1_000=6.64e-05 mcm5m4m1_cc_w_2_400_s_1_000=3.88e-11 mcm5m4m1_cf_w_2_400_s_1_000=2.69e-11
+  mcm5m4m1_ca_w_2_400_s_1_200=6.64e-05 mcm5m4m1_cc_w_2_400_s_1_200=3.14e-11 mcm5m4m1_cf_w_2_400_s_1_200=3.06e-11
+  mcm5m4m1_ca_w_2_400_s_2_100=6.64e-05 mcm5m4m1_cc_w_2_400_s_2_100=1.36e-11 mcm5m4m1_cf_w_2_400_s_2_100=4.22e-11
+  mcm5m4m1_ca_w_2_400_s_3_300=6.64e-05 mcm5m4m1_cc_w_2_400_s_3_300=4.97e-12 mcm5m4m1_cf_w_2_400_s_3_300=4.94e-11
+  mcm5m4m1_ca_w_2_400_s_9_000=6.64e-05 mcm5m4m1_cc_w_2_400_s_9_000=9.50e-14 mcm5m4m1_cf_w_2_400_s_9_000=5.42e-11
+  mcm5m4m2_ca_w_0_300_s_0_300=7.15e-05 mcm5m4m2_cc_w_0_300_s_0_300=8.25e-11 mcm5m4m2_cf_w_0_300_s_0_300=1.07e-11
+  mcm5m4m2_ca_w_0_300_s_0_360=7.15e-05 mcm5m4m2_cc_w_0_300_s_0_360=7.58e-11 mcm5m4m2_cf_w_0_300_s_0_360=1.26e-11
+  mcm5m4m2_ca_w_0_300_s_0_450=7.15e-05 mcm5m4m2_cc_w_0_300_s_0_450=6.69e-11 mcm5m4m2_cf_w_0_300_s_0_450=1.52e-11
+  mcm5m4m2_ca_w_0_300_s_0_600=7.15e-05 mcm5m4m2_cc_w_0_300_s_0_600=5.45e-11 mcm5m4m2_cf_w_0_300_s_0_600=1.94e-11
+  mcm5m4m2_ca_w_0_300_s_0_800=7.15e-05 mcm5m4m2_cc_w_0_300_s_0_800=4.22e-11 mcm5m4m2_cf_w_0_300_s_0_800=2.43e-11
+  mcm5m4m2_ca_w_0_300_s_1_000=7.15e-05 mcm5m4m2_cc_w_0_300_s_1_000=3.29e-11 mcm5m4m2_cf_w_0_300_s_1_000=2.88e-11
+  mcm5m4m2_ca_w_0_300_s_1_200=7.15e-05 mcm5m4m2_cc_w_0_300_s_1_200=2.60e-11 mcm5m4m2_cf_w_0_300_s_1_200=3.26e-11
+  mcm5m4m2_ca_w_0_300_s_2_100=7.15e-05 mcm5m4m2_cc_w_0_300_s_2_100=9.92e-12 mcm5m4m2_cf_w_0_300_s_2_100=4.39e-11
+  mcm5m4m2_ca_w_0_300_s_3_300=7.15e-05 mcm5m4m2_cc_w_0_300_s_3_300=3.04e-12 mcm5m4m2_cf_w_0_300_s_3_300=5.01e-11
+  mcm5m4m2_ca_w_0_300_s_9_000=7.15e-05 mcm5m4m2_cc_w_0_300_s_9_000=3.50e-14 mcm5m4m2_cf_w_0_300_s_9_000=5.30e-11
+  mcm5m4m2_ca_w_2_400_s_0_300=7.15e-05 mcm5m4m2_cc_w_2_400_s_0_300=8.88e-11 mcm5m4m2_cf_w_2_400_s_0_300=1.08e-11
+  mcm5m4m2_ca_w_2_400_s_0_360=7.15e-05 mcm5m4m2_cc_w_2_400_s_0_360=8.16e-11 mcm5m4m2_cf_w_2_400_s_0_360=1.26e-11
+  mcm5m4m2_ca_w_2_400_s_0_450=7.15e-05 mcm5m4m2_cc_w_2_400_s_0_450=7.18e-11 mcm5m4m2_cf_w_2_400_s_0_450=1.53e-11
+  mcm5m4m2_ca_w_2_400_s_0_600=7.15e-05 mcm5m4m2_cc_w_2_400_s_0_600=5.87e-11 mcm5m4m2_cf_w_2_400_s_0_600=1.95e-11
+  mcm5m4m2_ca_w_2_400_s_0_800=7.15e-05 mcm5m4m2_cc_w_2_400_s_0_800=4.55e-11 mcm5m4m2_cf_w_2_400_s_0_800=2.46e-11
+  mcm5m4m2_ca_w_2_400_s_1_000=7.15e-05 mcm5m4m2_cc_w_2_400_s_1_000=3.55e-11 mcm5m4m2_cf_w_2_400_s_1_000=2.91e-11
+  mcm5m4m2_ca_w_2_400_s_1_200=7.15e-05 mcm5m4m2_cc_w_2_400_s_1_200=2.81e-11 mcm5m4m2_cf_w_2_400_s_1_200=3.30e-11
+  mcm5m4m2_ca_w_2_400_s_2_100=7.15e-05 mcm5m4m2_cc_w_2_400_s_2_100=1.09e-11 mcm5m4m2_cf_w_2_400_s_2_100=4.49e-11
+  mcm5m4m2_ca_w_2_400_s_3_300=7.15e-05 mcm5m4m2_cc_w_2_400_s_3_300=3.38e-12 mcm5m4m2_cf_w_2_400_s_3_300=5.15e-11
+  mcm5m4m2_ca_w_2_400_s_9_000=7.15e-05 mcm5m4m2_cc_w_2_400_s_9_000=5.00e-14 mcm5m4m2_cf_w_2_400_s_9_000=5.48e-11
+  mcm5m4m3_ca_w_0_300_s_0_300=1.17e-04 mcm5m4m3_cc_w_0_300_s_0_300=7.39e-11 mcm5m4m3_cf_w_0_300_s_0_300=1.75e-11
+  mcm5m4m3_ca_w_0_300_s_0_360=1.17e-04 mcm5m4m3_cc_w_0_300_s_0_360=6.69e-11 mcm5m4m3_cf_w_0_300_s_0_360=2.03e-11
+  mcm5m4m3_ca_w_0_300_s_0_450=1.17e-04 mcm5m4m3_cc_w_0_300_s_0_450=5.75e-11 mcm5m4m3_cf_w_0_300_s_0_450=2.44e-11
+  mcm5m4m3_ca_w_0_300_s_0_600=1.17e-04 mcm5m4m3_cc_w_0_300_s_0_600=4.48e-11 mcm5m4m3_cf_w_0_300_s_0_600=3.07e-11
+  mcm5m4m3_ca_w_0_300_s_0_800=1.17e-04 mcm5m4m3_cc_w_0_300_s_0_800=3.21e-11 mcm5m4m3_cf_w_0_300_s_0_800=3.78e-11
+  mcm5m4m3_ca_w_0_300_s_1_000=1.17e-04 mcm5m4m3_cc_w_0_300_s_1_000=2.30e-11 mcm5m4m3_cf_w_0_300_s_1_000=4.38e-11
+  mcm5m4m3_ca_w_0_300_s_1_200=1.17e-04 mcm5m4m3_cc_w_0_300_s_1_200=1.65e-11 mcm5m4m3_cf_w_0_300_s_1_200=4.84e-11
+  mcm5m4m3_ca_w_0_300_s_2_100=1.17e-04 mcm5m4m3_cc_w_0_300_s_2_100=3.93e-12 mcm5m4m3_cf_w_0_300_s_2_100=5.92e-11
+  mcm5m4m3_ca_w_0_300_s_3_300=1.17e-04 mcm5m4m3_cc_w_0_300_s_3_300=6.25e-13 mcm5m4m3_cf_w_0_300_s_3_300=6.25e-11
+  mcm5m4m3_ca_w_0_300_s_9_000=1.17e-04 mcm5m4m3_cc_w_0_300_s_9_000=0.00e+00 mcm5m4m3_cf_w_0_300_s_9_000=6.31e-11
+  mcm5m4m3_ca_w_2_400_s_0_300=1.17e-04 mcm5m4m3_cc_w_2_400_s_0_300=7.56e-11 mcm5m4m3_cf_w_2_400_s_0_300=1.76e-11
+  mcm5m4m3_ca_w_2_400_s_0_360=1.17e-04 mcm5m4m3_cc_w_2_400_s_0_360=6.84e-11 mcm5m4m3_cf_w_2_400_s_0_360=2.05e-11
+  mcm5m4m3_ca_w_2_400_s_0_450=1.17e-04 mcm5m4m3_cc_w_2_400_s_0_450=5.87e-11 mcm5m4m3_cf_w_2_400_s_0_450=2.46e-11
+  mcm5m4m3_ca_w_2_400_s_0_600=1.17e-04 mcm5m4m3_cc_w_2_400_s_0_600=4.57e-11 mcm5m4m3_cf_w_2_400_s_0_600=3.08e-11
+  mcm5m4m3_ca_w_2_400_s_0_800=1.17e-04 mcm5m4m3_cc_w_2_400_s_0_800=3.27e-11 mcm5m4m3_cf_w_2_400_s_0_800=3.80e-11
+  mcm5m4m3_ca_w_2_400_s_1_000=1.17e-04 mcm5m4m3_cc_w_2_400_s_1_000=2.35e-11 mcm5m4m3_cf_w_2_400_s_1_000=4.41e-11
+  mcm5m4m3_ca_w_2_400_s_1_200=1.17e-04 mcm5m4m3_cc_w_2_400_s_1_200=1.69e-11 mcm5m4m3_cf_w_2_400_s_1_200=4.88e-11
+  mcm5m4m3_ca_w_2_400_s_2_100=1.17e-04 mcm5m4m3_cc_w_2_400_s_2_100=4.00e-12 mcm5m4m3_cf_w_2_400_s_2_100=5.98e-11
+  mcm5m4m3_ca_w_2_400_s_3_300=1.17e-04 mcm5m4m3_cc_w_2_400_s_3_300=7.00e-13 mcm5m4m3_cf_w_2_400_s_3_300=6.31e-11
+  mcm5m4m3_ca_w_2_400_s_9_000=1.17e-04 mcm5m4m3_cc_w_2_400_s_9_000=5.00e-14 mcm5m4m3_cf_w_2_400_s_9_000=6.38e-11
+  mcrdlm4f_ca_w_0_300_s_0_300=1.11e-05 mcrdlm4f_cc_w_0_300_s_0_300=9.59e-11 mcrdlm4f_cf_w_0_300_s_0_300=1.83e-12
+  mcrdlm4f_ca_w_0_300_s_0_360=1.11e-05 mcrdlm4f_cc_w_0_300_s_0_360=9.01e-11 mcrdlm4f_cf_w_0_300_s_0_360=2.16e-12
+  mcrdlm4f_ca_w_0_300_s_0_450=1.11e-05 mcrdlm4f_cc_w_0_300_s_0_450=8.21e-11 mcrdlm4f_cf_w_0_300_s_0_450=2.68e-12
+  mcrdlm4f_ca_w_0_300_s_0_600=1.11e-05 mcrdlm4f_cc_w_0_300_s_0_600=7.16e-11 mcrdlm4f_cf_w_0_300_s_0_600=3.52e-12
+  mcrdlm4f_ca_w_0_300_s_0_800=1.11e-05 mcrdlm4f_cc_w_0_300_s_0_800=6.14e-11 mcrdlm4f_cf_w_0_300_s_0_800=4.50e-12
+  mcrdlm4f_ca_w_0_300_s_1_000=1.11e-05 mcrdlm4f_cc_w_0_300_s_1_000=5.34e-11 mcrdlm4f_cf_w_0_300_s_1_000=5.52e-12
+  mcrdlm4f_ca_w_0_300_s_1_200=1.11e-05 mcrdlm4f_cc_w_0_300_s_1_200=4.75e-11 mcrdlm4f_cf_w_0_300_s_1_200=6.55e-12
+  mcrdlm4f_ca_w_0_300_s_2_100=1.11e-05 mcrdlm4f_cc_w_0_300_s_2_100=3.15e-11 mcrdlm4f_cf_w_0_300_s_2_100=1.10e-11
+  mcrdlm4f_ca_w_0_300_s_3_300=1.11e-05 mcrdlm4f_cc_w_0_300_s_3_300=2.12e-11 mcrdlm4f_cf_w_0_300_s_3_300=1.54e-11
+  mcrdlm4f_ca_w_0_300_s_9_000=1.11e-05 mcrdlm4f_cc_w_0_300_s_9_000=4.68e-12 mcrdlm4f_cf_w_0_300_s_9_000=2.70e-11
+  mcrdlm4f_ca_w_2_400_s_0_300=1.11e-05 mcrdlm4f_cc_w_2_400_s_0_300=1.21e-10 mcrdlm4f_cf_w_2_400_s_0_300=1.86e-12
+  mcrdlm4f_ca_w_2_400_s_0_360=1.11e-05 mcrdlm4f_cc_w_2_400_s_0_360=1.14e-10 mcrdlm4f_cf_w_2_400_s_0_360=2.19e-12
+  mcrdlm4f_ca_w_2_400_s_0_450=1.11e-05 mcrdlm4f_cc_w_2_400_s_0_450=1.05e-10 mcrdlm4f_cf_w_2_400_s_0_450=2.67e-12
+  mcrdlm4f_ca_w_2_400_s_0_600=1.11e-05 mcrdlm4f_cc_w_2_400_s_0_600=9.17e-11 mcrdlm4f_cf_w_2_400_s_0_600=3.48e-12
+  mcrdlm4f_ca_w_2_400_s_0_800=1.11e-05 mcrdlm4f_cc_w_2_400_s_0_800=7.85e-11 mcrdlm4f_cf_w_2_400_s_0_800=4.54e-12
+  mcrdlm4f_ca_w_2_400_s_1_000=1.11e-05 mcrdlm4f_cc_w_2_400_s_1_000=6.87e-11 mcrdlm4f_cf_w_2_400_s_1_000=5.59e-12
+  mcrdlm4f_ca_w_2_400_s_1_200=1.11e-05 mcrdlm4f_cc_w_2_400_s_1_200=6.10e-11 mcrdlm4f_cf_w_2_400_s_1_200=6.61e-12
+  mcrdlm4f_ca_w_2_400_s_2_100=1.11e-05 mcrdlm4f_cc_w_2_400_s_2_100=4.08e-11 mcrdlm4f_cf_w_2_400_s_2_100=1.09e-11
+  mcrdlm4f_ca_w_2_400_s_3_300=1.11e-05 mcrdlm4f_cc_w_2_400_s_3_300=2.74e-11 mcrdlm4f_cf_w_2_400_s_3_300=1.60e-11
+  mcrdlm4f_ca_w_2_400_s_9_000=1.11e-05 mcrdlm4f_cc_w_2_400_s_9_000=6.29e-12 mcrdlm4f_cf_w_2_400_s_9_000=2.97e-11
+  mcrdlm4d_ca_w_0_300_s_0_300=1.18e-05 mcrdlm4d_cc_w_0_300_s_0_300=9.57e-11 mcrdlm4d_cf_w_0_300_s_0_300=1.95e-12
+  mcrdlm4d_ca_w_0_300_s_0_360=1.18e-05 mcrdlm4d_cc_w_0_300_s_0_360=8.98e-11 mcrdlm4d_cf_w_0_300_s_0_360=2.30e-12
+  mcrdlm4d_ca_w_0_300_s_0_450=1.18e-05 mcrdlm4d_cc_w_0_300_s_0_450=8.19e-11 mcrdlm4d_cf_w_0_300_s_0_450=2.85e-12
+  mcrdlm4d_ca_w_0_300_s_0_600=1.18e-05 mcrdlm4d_cc_w_0_300_s_0_600=7.13e-11 mcrdlm4d_cf_w_0_300_s_0_600=3.74e-12
+  mcrdlm4d_ca_w_0_300_s_0_800=1.18e-05 mcrdlm4d_cc_w_0_300_s_0_800=6.11e-11 mcrdlm4d_cf_w_0_300_s_0_800=4.77e-12
+  mcrdlm4d_ca_w_0_300_s_1_000=1.18e-05 mcrdlm4d_cc_w_0_300_s_1_000=5.30e-11 mcrdlm4d_cf_w_0_300_s_1_000=5.86e-12
+  mcrdlm4d_ca_w_0_300_s_1_200=1.18e-05 mcrdlm4d_cc_w_0_300_s_1_200=4.70e-11 mcrdlm4d_cf_w_0_300_s_1_200=6.93e-12
+  mcrdlm4d_ca_w_0_300_s_2_100=1.18e-05 mcrdlm4d_cc_w_0_300_s_2_100=3.09e-11 mcrdlm4d_cf_w_0_300_s_2_100=1.16e-11
+  mcrdlm4d_ca_w_0_300_s_3_300=1.18e-05 mcrdlm4d_cc_w_0_300_s_3_300=2.07e-11 mcrdlm4d_cf_w_0_300_s_3_300=1.62e-11
+  mcrdlm4d_ca_w_0_300_s_9_000=1.18e-05 mcrdlm4d_cc_w_0_300_s_9_000=4.33e-12 mcrdlm4d_cf_w_0_300_s_9_000=2.78e-11
+  mcrdlm4d_ca_w_2_400_s_0_300=1.18e-05 mcrdlm4d_cc_w_2_400_s_0_300=1.21e-10 mcrdlm4d_cf_w_2_400_s_0_300=1.97e-12
+  mcrdlm4d_ca_w_2_400_s_0_360=1.18e-05 mcrdlm4d_cc_w_2_400_s_0_360=1.13e-10 mcrdlm4d_cf_w_2_400_s_0_360=2.32e-12
+  mcrdlm4d_ca_w_2_400_s_0_450=1.18e-05 mcrdlm4d_cc_w_2_400_s_0_450=1.04e-10 mcrdlm4d_cf_w_2_400_s_0_450=2.84e-12
+  mcrdlm4d_ca_w_2_400_s_0_600=1.18e-05 mcrdlm4d_cc_w_2_400_s_0_600=9.11e-11 mcrdlm4d_cf_w_2_400_s_0_600=3.69e-12
+  mcrdlm4d_ca_w_2_400_s_0_800=1.18e-05 mcrdlm4d_cc_w_2_400_s_0_800=7.78e-11 mcrdlm4d_cf_w_2_400_s_0_800=4.82e-12
+  mcrdlm4d_ca_w_2_400_s_1_000=1.18e-05 mcrdlm4d_cc_w_2_400_s_1_000=6.79e-11 mcrdlm4d_cf_w_2_400_s_1_000=5.92e-12
+  mcrdlm4d_ca_w_2_400_s_1_200=1.18e-05 mcrdlm4d_cc_w_2_400_s_1_200=6.02e-11 mcrdlm4d_cf_w_2_400_s_1_200=7.01e-12
+  mcrdlm4d_ca_w_2_400_s_2_100=1.18e-05 mcrdlm4d_cc_w_2_400_s_2_100=4.00e-11 mcrdlm4d_cf_w_2_400_s_2_100=1.16e-11
+  mcrdlm4d_ca_w_2_400_s_3_300=1.18e-05 mcrdlm4d_cc_w_2_400_s_3_300=2.66e-11 mcrdlm4d_cf_w_2_400_s_3_300=1.68e-11
+  mcrdlm4d_ca_w_2_400_s_9_000=1.18e-05 mcrdlm4d_cc_w_2_400_s_9_000=5.79e-12 mcrdlm4d_cf_w_2_400_s_9_000=3.07e-11
+  mcrdlm4p1_ca_w_0_300_s_0_300=1.23e-05 mcrdlm4p1_cc_w_0_300_s_0_300=9.56e-11 mcrdlm4p1_cf_w_0_300_s_0_300=2.03e-12
+  mcrdlm4p1_ca_w_0_300_s_0_360=1.23e-05 mcrdlm4p1_cc_w_0_300_s_0_360=8.97e-11 mcrdlm4p1_cf_w_0_300_s_0_360=2.40e-12
+  mcrdlm4p1_ca_w_0_300_s_0_450=1.23e-05 mcrdlm4p1_cc_w_0_300_s_0_450=8.17e-11 mcrdlm4p1_cf_w_0_300_s_0_450=2.97e-12
+  mcrdlm4p1_ca_w_0_300_s_0_600=1.23e-05 mcrdlm4p1_cc_w_0_300_s_0_600=7.12e-11 mcrdlm4p1_cf_w_0_300_s_0_600=3.90e-12
+  mcrdlm4p1_ca_w_0_300_s_0_800=1.23e-05 mcrdlm4p1_cc_w_0_300_s_0_800=6.08e-11 mcrdlm4p1_cf_w_0_300_s_0_800=4.98e-12
+  mcrdlm4p1_ca_w_0_300_s_1_000=1.23e-05 mcrdlm4p1_cc_w_0_300_s_1_000=5.28e-11 mcrdlm4p1_cf_w_0_300_s_1_000=6.10e-12
+  mcrdlm4p1_ca_w_0_300_s_1_200=1.23e-05 mcrdlm4p1_cc_w_0_300_s_1_200=4.67e-11 mcrdlm4p1_cf_w_0_300_s_1_200=7.21e-12
+  mcrdlm4p1_ca_w_0_300_s_2_100=1.23e-05 mcrdlm4p1_cc_w_0_300_s_2_100=3.06e-11 mcrdlm4p1_cf_w_0_300_s_2_100=1.20e-11
+  mcrdlm4p1_ca_w_0_300_s_3_300=1.23e-05 mcrdlm4p1_cc_w_0_300_s_3_300=2.02e-11 mcrdlm4p1_cf_w_0_300_s_3_300=1.68e-11
+  mcrdlm4p1_ca_w_0_300_s_9_000=1.23e-05 mcrdlm4p1_cc_w_0_300_s_9_000=4.09e-12 mcrdlm4p1_cf_w_0_300_s_9_000=2.85e-11
+  mcrdlm4p1_ca_w_2_400_s_0_300=1.23e-05 mcrdlm4p1_cc_w_2_400_s_0_300=1.20e-10 mcrdlm4p1_cf_w_2_400_s_0_300=2.07e-12
+  mcrdlm4p1_ca_w_2_400_s_0_360=1.23e-05 mcrdlm4p1_cc_w_2_400_s_0_360=1.13e-10 mcrdlm4p1_cf_w_2_400_s_0_360=2.43e-12
+  mcrdlm4p1_ca_w_2_400_s_0_450=1.23e-05 mcrdlm4p1_cc_w_2_400_s_0_450=1.03e-10 mcrdlm4p1_cf_w_2_400_s_0_450=2.97e-12
+  mcrdlm4p1_ca_w_2_400_s_0_600=1.23e-05 mcrdlm4p1_cc_w_2_400_s_0_600=9.05e-11 mcrdlm4p1_cf_w_2_400_s_0_600=3.86e-12
+  mcrdlm4p1_ca_w_2_400_s_0_800=1.23e-05 mcrdlm4p1_cc_w_2_400_s_0_800=7.73e-11 mcrdlm4p1_cf_w_2_400_s_0_800=5.04e-12
+  mcrdlm4p1_ca_w_2_400_s_1_000=1.23e-05 mcrdlm4p1_cc_w_2_400_s_1_000=6.74e-11 mcrdlm4p1_cf_w_2_400_s_1_000=6.18e-12
+  mcrdlm4p1_ca_w_2_400_s_1_200=1.23e-05 mcrdlm4p1_cc_w_2_400_s_1_200=5.97e-11 mcrdlm4p1_cf_w_2_400_s_1_200=7.31e-12
+  mcrdlm4p1_ca_w_2_400_s_2_100=1.23e-05 mcrdlm4p1_cc_w_2_400_s_2_100=3.94e-11 mcrdlm4p1_cf_w_2_400_s_2_100=1.20e-11
+  mcrdlm4p1_ca_w_2_400_s_3_300=1.23e-05 mcrdlm4p1_cc_w_2_400_s_3_300=2.60e-11 mcrdlm4p1_cf_w_2_400_s_3_300=1.74e-11
+  mcrdlm4p1_ca_w_2_400_s_9_000=1.23e-05 mcrdlm4p1_cc_w_2_400_s_9_000=5.51e-12 mcrdlm4p1_cf_w_2_400_s_9_000=3.13e-11
+  mcrdlm4l1_ca_w_0_300_s_0_300=1.39e-05 mcrdlm4l1_cc_w_0_300_s_0_300=9.52e-11 mcrdlm4l1_cf_w_0_300_s_0_300=2.28e-12
+  mcrdlm4l1_ca_w_0_300_s_0_360=1.39e-05 mcrdlm4l1_cc_w_0_300_s_0_360=8.93e-11 mcrdlm4l1_cf_w_0_300_s_0_360=2.69e-12
+  mcrdlm4l1_ca_w_0_300_s_0_450=1.39e-05 mcrdlm4l1_cc_w_0_300_s_0_450=8.13e-11 mcrdlm4l1_cf_w_0_300_s_0_450=3.32e-12
+  mcrdlm4l1_ca_w_0_300_s_0_600=1.39e-05 mcrdlm4l1_cc_w_0_300_s_0_600=7.06e-11 mcrdlm4l1_cf_w_0_300_s_0_600=4.36e-12
+  mcrdlm4l1_ca_w_0_300_s_0_800=1.39e-05 mcrdlm4l1_cc_w_0_300_s_0_800=6.02e-11 mcrdlm4l1_cf_w_0_300_s_0_800=5.56e-12
+  mcrdlm4l1_ca_w_0_300_s_1_000=1.39e-05 mcrdlm4l1_cc_w_0_300_s_1_000=5.20e-11 mcrdlm4l1_cf_w_0_300_s_1_000=6.81e-12
+  mcrdlm4l1_ca_w_0_300_s_1_200=1.39e-05 mcrdlm4l1_cc_w_0_300_s_1_200=4.58e-11 mcrdlm4l1_cf_w_0_300_s_1_200=8.02e-12
+  mcrdlm4l1_ca_w_0_300_s_2_100=1.39e-05 mcrdlm4l1_cc_w_0_300_s_2_100=2.96e-11 mcrdlm4l1_cf_w_0_300_s_2_100=1.32e-11
+  mcrdlm4l1_ca_w_0_300_s_3_300=1.39e-05 mcrdlm4l1_cc_w_0_300_s_3_300=1.91e-11 mcrdlm4l1_cf_w_0_300_s_3_300=1.84e-11
+  mcrdlm4l1_ca_w_0_300_s_9_000=1.39e-05 mcrdlm4l1_cc_w_0_300_s_9_000=3.53e-12 mcrdlm4l1_cf_w_0_300_s_9_000=3.00e-11
+  mcrdlm4l1_ca_w_2_400_s_0_300=1.39e-05 mcrdlm4l1_cc_w_2_400_s_0_300=1.19e-10 mcrdlm4l1_cf_w_2_400_s_0_300=2.30e-12
+  mcrdlm4l1_ca_w_2_400_s_0_360=1.39e-05 mcrdlm4l1_cc_w_2_400_s_0_360=1.12e-10 mcrdlm4l1_cf_w_2_400_s_0_360=2.71e-12
+  mcrdlm4l1_ca_w_2_400_s_0_450=1.39e-05 mcrdlm4l1_cc_w_2_400_s_0_450=1.02e-10 mcrdlm4l1_cf_w_2_400_s_0_450=3.31e-12
+  mcrdlm4l1_ca_w_2_400_s_0_600=1.39e-05 mcrdlm4l1_cc_w_2_400_s_0_600=8.92e-11 mcrdlm4l1_cf_w_2_400_s_0_600=4.31e-12
+  mcrdlm4l1_ca_w_2_400_s_0_800=1.39e-05 mcrdlm4l1_cc_w_2_400_s_0_800=7.59e-11 mcrdlm4l1_cf_w_2_400_s_0_800=5.61e-12
+  mcrdlm4l1_ca_w_2_400_s_1_000=1.39e-05 mcrdlm4l1_cc_w_2_400_s_1_000=6.59e-11 mcrdlm4l1_cf_w_2_400_s_1_000=6.88e-12
+  mcrdlm4l1_ca_w_2_400_s_1_200=1.39e-05 mcrdlm4l1_cc_w_2_400_s_1_200=5.82e-11 mcrdlm4l1_cf_w_2_400_s_1_200=8.13e-12
+  mcrdlm4l1_ca_w_2_400_s_2_100=1.39e-05 mcrdlm4l1_cc_w_2_400_s_2_100=3.79e-11 mcrdlm4l1_cf_w_2_400_s_2_100=1.33e-11
+  mcrdlm4l1_ca_w_2_400_s_3_300=1.39e-05 mcrdlm4l1_cc_w_2_400_s_3_300=2.46e-11 mcrdlm4l1_cf_w_2_400_s_3_300=1.91e-11
+  mcrdlm4l1_ca_w_2_400_s_9_000=1.39e-05 mcrdlm4l1_cc_w_2_400_s_9_000=4.75e-12 mcrdlm4l1_cf_w_2_400_s_9_000=3.31e-11
+  mcrdlm4m1_ca_w_0_300_s_0_300=1.68e-05 mcrdlm4m1_cc_w_0_300_s_0_300=9.45e-11 mcrdlm4m1_cf_w_0_300_s_0_300=2.75e-12
+  mcrdlm4m1_ca_w_0_300_s_0_360=1.68e-05 mcrdlm4m1_cc_w_0_300_s_0_360=8.85e-11 mcrdlm4m1_cf_w_0_300_s_0_360=3.24e-12
+  mcrdlm4m1_ca_w_0_300_s_0_450=1.68e-05 mcrdlm4m1_cc_w_0_300_s_0_450=8.04e-11 mcrdlm4m1_cf_w_0_300_s_0_450=4.00e-12
+  mcrdlm4m1_ca_w_0_300_s_0_600=1.68e-05 mcrdlm4m1_cc_w_0_300_s_0_600=6.96e-11 mcrdlm4m1_cf_w_0_300_s_0_600=5.23e-12
+  mcrdlm4m1_ca_w_0_300_s_0_800=1.68e-05 mcrdlm4m1_cc_w_0_300_s_0_800=5.90e-11 mcrdlm4m1_cf_w_0_300_s_0_800=6.68e-12
+  mcrdlm4m1_ca_w_0_300_s_1_000=1.68e-05 mcrdlm4m1_cc_w_0_300_s_1_000=5.07e-11 mcrdlm4m1_cf_w_0_300_s_1_000=8.13e-12
+  mcrdlm4m1_ca_w_0_300_s_1_200=1.68e-05 mcrdlm4m1_cc_w_0_300_s_1_200=4.45e-11 mcrdlm4m1_cf_w_0_300_s_1_200=9.59e-12
+  mcrdlm4m1_ca_w_0_300_s_2_100=1.68e-05 mcrdlm4m1_cc_w_0_300_s_2_100=2.78e-11 mcrdlm4m1_cf_w_0_300_s_2_100=1.56e-11
+  mcrdlm4m1_ca_w_0_300_s_3_300=1.68e-05 mcrdlm4m1_cc_w_0_300_s_3_300=1.73e-11 mcrdlm4m1_cf_w_0_300_s_3_300=2.12e-11
+  mcrdlm4m1_ca_w_0_300_s_9_000=1.68e-05 mcrdlm4m1_cc_w_0_300_s_9_000=2.73e-12 mcrdlm4m1_cf_w_0_300_s_9_000=3.27e-11
+  mcrdlm4m1_ca_w_2_400_s_0_300=1.68e-05 mcrdlm4m1_cc_w_2_400_s_0_300=1.17e-10 mcrdlm4m1_cf_w_2_400_s_0_300=2.77e-12
+  mcrdlm4m1_ca_w_2_400_s_0_360=1.68e-05 mcrdlm4m1_cc_w_2_400_s_0_360=1.10e-10 mcrdlm4m1_cf_w_2_400_s_0_360=3.25e-12
+  mcrdlm4m1_ca_w_2_400_s_0_450=1.68e-05 mcrdlm4m1_cc_w_2_400_s_0_450=9.97e-11 mcrdlm4m1_cf_w_2_400_s_0_450=3.98e-12
+  mcrdlm4m1_ca_w_2_400_s_0_600=1.68e-05 mcrdlm4m1_cc_w_2_400_s_0_600=8.68e-11 mcrdlm4m1_cf_w_2_400_s_0_600=5.17e-12
+  mcrdlm4m1_ca_w_2_400_s_0_800=1.68e-05 mcrdlm4m1_cc_w_2_400_s_0_800=7.35e-11 mcrdlm4m1_cf_w_2_400_s_0_800=6.73e-12
+  mcrdlm4m1_ca_w_2_400_s_1_000=1.68e-05 mcrdlm4m1_cc_w_2_400_s_1_000=6.35e-11 mcrdlm4m1_cf_w_2_400_s_1_000=8.24e-12
+  mcrdlm4m1_ca_w_2_400_s_1_200=1.68e-05 mcrdlm4m1_cc_w_2_400_s_1_200=5.57e-11 mcrdlm4m1_cf_w_2_400_s_1_200=9.70e-12
+  mcrdlm4m1_ca_w_2_400_s_2_100=1.68e-05 mcrdlm4m1_cc_w_2_400_s_2_100=3.54e-11 mcrdlm4m1_cf_w_2_400_s_2_100=1.57e-11
+  mcrdlm4m1_ca_w_2_400_s_3_300=1.68e-05 mcrdlm4m1_cc_w_2_400_s_3_300=2.23e-11 mcrdlm4m1_cf_w_2_400_s_3_300=2.21e-11
+  mcrdlm4m1_ca_w_2_400_s_9_000=1.68e-05 mcrdlm4m1_cc_w_2_400_s_9_000=3.74e-12 mcrdlm4m1_cf_w_2_400_s_9_000=3.60e-11
+  mcrdlm4m2_ca_w_0_300_s_0_300=2.20e-05 mcrdlm4m2_cc_w_0_300_s_0_300=9.32e-11 mcrdlm4m2_cf_w_0_300_s_0_300=3.58e-12
+  mcrdlm4m2_ca_w_0_300_s_0_360=2.20e-05 mcrdlm4m2_cc_w_0_300_s_0_360=8.70e-11 mcrdlm4m2_cf_w_0_300_s_0_360=4.21e-12
+  mcrdlm4m2_ca_w_0_300_s_0_450=2.20e-05 mcrdlm4m2_cc_w_0_300_s_0_450=7.89e-11 mcrdlm4m2_cf_w_0_300_s_0_450=5.17e-12
+  mcrdlm4m2_ca_w_0_300_s_0_600=2.20e-05 mcrdlm4m2_cc_w_0_300_s_0_600=6.78e-11 mcrdlm4m2_cf_w_0_300_s_0_600=6.73e-12
+  mcrdlm4m2_ca_w_0_300_s_0_800=2.20e-05 mcrdlm4m2_cc_w_0_300_s_0_800=5.71e-11 mcrdlm4m2_cf_w_0_300_s_0_800=8.59e-12
+  mcrdlm4m2_ca_w_0_300_s_1_000=2.20e-05 mcrdlm4m2_cc_w_0_300_s_1_000=4.85e-11 mcrdlm4m2_cf_w_0_300_s_1_000=1.04e-11
+  mcrdlm4m2_ca_w_0_300_s_1_200=2.20e-05 mcrdlm4m2_cc_w_0_300_s_1_200=4.22e-11 mcrdlm4m2_cf_w_0_300_s_1_200=1.22e-11
+  mcrdlm4m2_ca_w_0_300_s_2_100=2.20e-05 mcrdlm4m2_cc_w_0_300_s_2_100=2.52e-11 mcrdlm4m2_cf_w_0_300_s_2_100=1.93e-11
+  mcrdlm4m2_ca_w_0_300_s_3_300=2.20e-05 mcrdlm4m2_cc_w_0_300_s_3_300=1.49e-11 mcrdlm4m2_cf_w_0_300_s_3_300=2.56e-11
+  mcrdlm4m2_ca_w_0_300_s_9_000=2.20e-05 mcrdlm4m2_cc_w_0_300_s_9_000=1.97e-12 mcrdlm4m2_cf_w_0_300_s_9_000=3.64e-11
+  mcrdlm4m2_ca_w_2_400_s_0_300=2.20e-05 mcrdlm4m2_cc_w_2_400_s_0_300=1.13e-10 mcrdlm4m2_cf_w_2_400_s_0_300=3.60e-12
+  mcrdlm4m2_ca_w_2_400_s_0_360=2.20e-05 mcrdlm4m2_cc_w_2_400_s_0_360=1.06e-10 mcrdlm4m2_cf_w_2_400_s_0_360=4.22e-12
+  mcrdlm4m2_ca_w_2_400_s_0_450=2.20e-05 mcrdlm4m2_cc_w_2_400_s_0_450=9.65e-11 mcrdlm4m2_cf_w_2_400_s_0_450=5.17e-12
+  mcrdlm4m2_ca_w_2_400_s_0_600=2.20e-05 mcrdlm4m2_cc_w_2_400_s_0_600=8.34e-11 mcrdlm4m2_cf_w_2_400_s_0_600=6.68e-12
+  mcrdlm4m2_ca_w_2_400_s_0_800=2.20e-05 mcrdlm4m2_cc_w_2_400_s_0_800=7.02e-11 mcrdlm4m2_cf_w_2_400_s_0_800=8.65e-12
+  mcrdlm4m2_ca_w_2_400_s_1_000=2.20e-05 mcrdlm4m2_cc_w_2_400_s_1_000=6.01e-11 mcrdlm4m2_cf_w_2_400_s_1_000=1.05e-11
+  mcrdlm4m2_ca_w_2_400_s_1_200=2.20e-05 mcrdlm4m2_cc_w_2_400_s_1_200=5.23e-11 mcrdlm4m2_cf_w_2_400_s_1_200=1.24e-11
+  mcrdlm4m2_ca_w_2_400_s_2_100=2.20e-05 mcrdlm4m2_cc_w_2_400_s_2_100=3.22e-11 mcrdlm4m2_cf_w_2_400_s_2_100=1.95e-11
+  mcrdlm4m2_ca_w_2_400_s_3_300=2.20e-05 mcrdlm4m2_cc_w_2_400_s_3_300=1.94e-11 mcrdlm4m2_cf_w_2_400_s_3_300=2.67e-11
+  mcrdlm4m2_ca_w_2_400_s_9_000=2.20e-05 mcrdlm4m2_cc_w_2_400_s_9_000=2.78e-12 mcrdlm4m2_cf_w_2_400_s_9_000=4.01e-11
+  mcrdlm4m3_ca_w_0_300_s_0_300=6.78e-05 mcrdlm4m3_cc_w_0_300_s_0_300=8.45e-11 mcrdlm4m3_cf_w_0_300_s_0_300=1.03e-11
+  mcrdlm4m3_ca_w_0_300_s_0_360=6.78e-05 mcrdlm4m3_cc_w_0_300_s_0_360=7.82e-11 mcrdlm4m3_cf_w_0_300_s_0_360=1.20e-11
+  mcrdlm4m3_ca_w_0_300_s_0_450=6.78e-05 mcrdlm4m3_cc_w_0_300_s_0_450=6.95e-11 mcrdlm4m3_cf_w_0_300_s_0_450=1.44e-11
+  mcrdlm4m3_ca_w_0_300_s_0_600=6.78e-05 mcrdlm4m3_cc_w_0_300_s_0_600=5.79e-11 mcrdlm4m3_cf_w_0_300_s_0_600=1.81e-11
+  mcrdlm4m3_ca_w_0_300_s_0_800=6.78e-05 mcrdlm4m3_cc_w_0_300_s_0_800=4.67e-11 mcrdlm4m3_cf_w_0_300_s_0_800=2.24e-11
+  mcrdlm4m3_ca_w_0_300_s_1_000=6.78e-05 mcrdlm4m3_cc_w_0_300_s_1_000=3.82e-11 mcrdlm4m3_cf_w_0_300_s_1_000=2.62e-11
+  mcrdlm4m3_ca_w_0_300_s_1_200=6.78e-05 mcrdlm4m3_cc_w_0_300_s_1_200=3.17e-11 mcrdlm4m3_cf_w_0_300_s_1_200=2.95e-11
+  mcrdlm4m3_ca_w_0_300_s_2_100=6.78e-05 mcrdlm4m3_cc_w_0_300_s_2_100=1.57e-11 mcrdlm4m3_cf_w_0_300_s_2_100=4.01e-11
+  mcrdlm4m3_ca_w_0_300_s_3_300=6.78e-05 mcrdlm4m3_cc_w_0_300_s_3_300=7.87e-12 mcrdlm4m3_cf_w_0_300_s_3_300=4.68e-11
+  mcrdlm4m3_ca_w_0_300_s_9_000=6.78e-05 mcrdlm4m3_cc_w_0_300_s_9_000=6.61e-13 mcrdlm4m3_cf_w_0_300_s_9_000=5.35e-11
+  mcrdlm4m3_ca_w_2_400_s_0_300=6.78e-05 mcrdlm4m3_cc_w_2_400_s_0_300=9.99e-11 mcrdlm4m3_cf_w_2_400_s_0_300=1.04e-11
+  mcrdlm4m3_ca_w_2_400_s_0_360=6.78e-05 mcrdlm4m3_cc_w_2_400_s_0_360=9.27e-11 mcrdlm4m3_cf_w_2_400_s_0_360=1.20e-11
+  mcrdlm4m3_ca_w_2_400_s_0_450=6.78e-05 mcrdlm4m3_cc_w_2_400_s_0_450=8.32e-11 mcrdlm4m3_cf_w_2_400_s_0_450=1.44e-11
+  mcrdlm4m3_ca_w_2_400_s_0_600=6.78e-05 mcrdlm4m3_cc_w_2_400_s_0_600=7.03e-11 mcrdlm4m3_cf_w_2_400_s_0_600=1.81e-11
+  mcrdlm4m3_ca_w_2_400_s_0_800=6.78e-05 mcrdlm4m3_cc_w_2_400_s_0_800=5.73e-11 mcrdlm4m3_cf_w_2_400_s_0_800=2.25e-11
+  mcrdlm4m3_ca_w_2_400_s_1_000=6.78e-05 mcrdlm4m3_cc_w_2_400_s_1_000=4.77e-11 mcrdlm4m3_cf_w_2_400_s_1_000=2.63e-11
+  mcrdlm4m3_ca_w_2_400_s_1_200=6.78e-05 mcrdlm4m3_cc_w_2_400_s_1_200=4.03e-11 mcrdlm4m3_cf_w_2_400_s_1_200=2.97e-11
+  mcrdlm4m3_ca_w_2_400_s_2_100=6.78e-05 mcrdlm4m3_cc_w_2_400_s_2_100=2.21e-11 mcrdlm4m3_cf_w_2_400_s_2_100=4.06e-11
+  mcrdlm4m3_ca_w_2_400_s_3_300=6.78e-05 mcrdlm4m3_cc_w_2_400_s_3_300=1.18e-11 mcrdlm4m3_cf_w_2_400_s_3_300=4.87e-11
+  mcrdlm4m3_ca_w_2_400_s_9_000=6.78e-05 mcrdlm4m3_cc_w_2_400_s_9_000=1.13e-12 mcrdlm4m3_cf_w_2_400_s_9_000=5.85e-11
+  mcrdlm5f_ca_w_1_600_s_1_600=1.04e-05 mcrdlm5f_cc_w_1_600_s_1_600=6.16e-11 mcrdlm5f_cf_w_1_600_s_1_600=8.33e-12
+  mcrdlm5f_ca_w_1_600_s_1_700=1.04e-05 mcrdlm5f_cc_w_1_600_s_1_700=5.84e-11 mcrdlm5f_cf_w_1_600_s_1_700=8.79e-12
+  mcrdlm5f_ca_w_1_600_s_1_900=1.04e-05 mcrdlm5f_cc_w_1_600_s_1_900=5.29e-11 mcrdlm5f_cf_w_1_600_s_1_900=9.71e-12
+  mcrdlm5f_ca_w_1_600_s_2_000=1.04e-05 mcrdlm5f_cc_w_1_600_s_2_000=5.06e-11 mcrdlm5f_cf_w_1_600_s_2_000=1.02e-11
+  mcrdlm5f_ca_w_1_600_s_2_400=1.04e-05 mcrdlm5f_cc_w_1_600_s_2_400=4.29e-11 mcrdlm5f_cf_w_1_600_s_2_400=1.19e-11
+  mcrdlm5f_ca_w_1_600_s_2_800=1.04e-05 mcrdlm5f_cc_w_1_600_s_2_800=3.71e-11 mcrdlm5f_cf_w_1_600_s_2_800=1.36e-11
+  mcrdlm5f_ca_w_1_600_s_3_200=1.04e-05 mcrdlm5f_cc_w_1_600_s_3_200=3.24e-11 mcrdlm5f_cf_w_1_600_s_3_200=1.52e-11
+  mcrdlm5f_ca_w_1_600_s_4_800=1.04e-05 mcrdlm5f_cc_w_1_600_s_4_800=2.03e-11 mcrdlm5f_cf_w_1_600_s_4_800=2.09e-11
+  mcrdlm5f_ca_w_1_600_s_10_000=1.04e-05 mcrdlm5f_cc_w_1_600_s_10_000=5.58e-12 mcrdlm5f_cf_w_1_600_s_10_000=3.13e-11
+  mcrdlm5f_ca_w_1_600_s_12_000=1.04e-05 mcrdlm5f_cc_w_1_600_s_12_000=3.48e-12 mcrdlm5f_cf_w_1_600_s_12_000=3.31e-11
+  mcrdlm5f_ca_w_4_000_s_1_600=1.04e-05 mcrdlm5f_cc_w_4_000_s_1_600=6.53e-11 mcrdlm5f_cf_w_4_000_s_1_600=8.33e-12
+  mcrdlm5f_ca_w_4_000_s_1_700=1.04e-05 mcrdlm5f_cc_w_4_000_s_1_700=6.21e-11 mcrdlm5f_cf_w_4_000_s_1_700=8.80e-12
+  mcrdlm5f_ca_w_4_000_s_1_900=1.04e-05 mcrdlm5f_cc_w_4_000_s_1_900=5.63e-11 mcrdlm5f_cf_w_4_000_s_1_900=9.73e-12
+  mcrdlm5f_ca_w_4_000_s_2_000=1.04e-05 mcrdlm5f_cc_w_4_000_s_2_000=5.38e-11 mcrdlm5f_cf_w_4_000_s_2_000=1.02e-11
+  mcrdlm5f_ca_w_4_000_s_2_400=1.04e-05 mcrdlm5f_cc_w_4_000_s_2_400=4.57e-11 mcrdlm5f_cf_w_4_000_s_2_400=1.20e-11
+  mcrdlm5f_ca_w_4_000_s_2_800=1.04e-05 mcrdlm5f_cc_w_4_000_s_2_800=3.94e-11 mcrdlm5f_cf_w_4_000_s_2_800=1.37e-11
+  mcrdlm5f_ca_w_4_000_s_3_200=1.04e-05 mcrdlm5f_cc_w_4_000_s_3_200=3.45e-11 mcrdlm5f_cf_w_4_000_s_3_200=1.53e-11
+  mcrdlm5f_ca_w_4_000_s_4_800=1.04e-05 mcrdlm5f_cc_w_4_000_s_4_800=2.17e-11 mcrdlm5f_cf_w_4_000_s_4_800=2.11e-11
+  mcrdlm5f_ca_w_4_000_s_10_000=1.04e-05 mcrdlm5f_cc_w_4_000_s_10_000=6.03e-12 mcrdlm5f_cf_w_4_000_s_10_000=3.20e-11
+  mcrdlm5f_ca_w_4_000_s_12_000=1.04e-05 mcrdlm5f_cc_w_4_000_s_12_000=3.78e-12 mcrdlm5f_cf_w_4_000_s_12_000=3.40e-11
+  mcrdlm5d_ca_w_1_600_s_1_600=1.08e-05 mcrdlm5d_cc_w_1_600_s_1_600=6.11e-11 mcrdlm5d_cf_w_1_600_s_1_600=8.63e-12
+  mcrdlm5d_ca_w_1_600_s_1_700=1.08e-05 mcrdlm5d_cc_w_1_600_s_1_700=5.80e-11 mcrdlm5d_cf_w_1_600_s_1_700=9.12e-12
+  mcrdlm5d_ca_w_1_600_s_1_900=1.08e-05 mcrdlm5d_cc_w_1_600_s_1_900=5.24e-11 mcrdlm5d_cf_w_1_600_s_1_900=1.01e-11
+  mcrdlm5d_ca_w_1_600_s_2_000=1.08e-05 mcrdlm5d_cc_w_1_600_s_2_000=5.02e-11 mcrdlm5d_cf_w_1_600_s_2_000=1.05e-11
+  mcrdlm5d_ca_w_1_600_s_2_400=1.08e-05 mcrdlm5d_cc_w_1_600_s_2_400=4.25e-11 mcrdlm5d_cf_w_1_600_s_2_400=1.24e-11
+  mcrdlm5d_ca_w_1_600_s_2_800=1.08e-05 mcrdlm5d_cc_w_1_600_s_2_800=3.66e-11 mcrdlm5d_cf_w_1_600_s_2_800=1.41e-11
+  mcrdlm5d_ca_w_1_600_s_3_200=1.08e-05 mcrdlm5d_cc_w_1_600_s_3_200=3.19e-11 mcrdlm5d_cf_w_1_600_s_3_200=1.58e-11
+  mcrdlm5d_ca_w_1_600_s_4_800=1.08e-05 mcrdlm5d_cc_w_1_600_s_4_800=1.98e-11 mcrdlm5d_cf_w_1_600_s_4_800=2.15e-11
+  mcrdlm5d_ca_w_1_600_s_10_000=1.08e-05 mcrdlm5d_cc_w_1_600_s_10_000=5.24e-12 mcrdlm5d_cf_w_1_600_s_10_000=3.20e-11
+  mcrdlm5d_ca_w_1_600_s_12_000=1.08e-05 mcrdlm5d_cc_w_1_600_s_12_000=3.22e-12 mcrdlm5d_cf_w_1_600_s_12_000=3.38e-11
+  mcrdlm5d_ca_w_4_000_s_1_600=1.08e-05 mcrdlm5d_cc_w_4_000_s_1_600=6.47e-11 mcrdlm5d_cf_w_4_000_s_1_600=8.64e-12
+  mcrdlm5d_ca_w_4_000_s_1_700=1.08e-05 mcrdlm5d_cc_w_4_000_s_1_700=6.15e-11 mcrdlm5d_cf_w_4_000_s_1_700=9.13e-12
+  mcrdlm5d_ca_w_4_000_s_1_900=1.08e-05 mcrdlm5d_cc_w_4_000_s_1_900=5.57e-11 mcrdlm5d_cf_w_4_000_s_1_900=1.01e-11
+  mcrdlm5d_ca_w_4_000_s_2_000=1.08e-05 mcrdlm5d_cc_w_4_000_s_2_000=5.32e-11 mcrdlm5d_cf_w_4_000_s_2_000=1.06e-11
+  mcrdlm5d_ca_w_4_000_s_2_400=1.08e-05 mcrdlm5d_cc_w_4_000_s_2_400=4.50e-11 mcrdlm5d_cf_w_4_000_s_2_400=1.24e-11
+  mcrdlm5d_ca_w_4_000_s_2_800=1.08e-05 mcrdlm5d_cc_w_4_000_s_2_800=3.87e-11 mcrdlm5d_cf_w_4_000_s_2_800=1.42e-11
+  mcrdlm5d_ca_w_4_000_s_3_200=1.08e-05 mcrdlm5d_cc_w_4_000_s_3_200=3.39e-11 mcrdlm5d_cf_w_4_000_s_3_200=1.59e-11
+  mcrdlm5d_ca_w_4_000_s_4_800=1.08e-05 mcrdlm5d_cc_w_4_000_s_4_800=2.11e-11 mcrdlm5d_cf_w_4_000_s_4_800=2.17e-11
+  mcrdlm5d_ca_w_4_000_s_10_000=1.08e-05 mcrdlm5d_cc_w_4_000_s_10_000=5.66e-12 mcrdlm5d_cf_w_4_000_s_10_000=3.27e-11
+  mcrdlm5d_ca_w_4_000_s_12_000=1.08e-05 mcrdlm5d_cc_w_4_000_s_12_000=3.47e-12 mcrdlm5d_cf_w_4_000_s_12_000=3.46e-11
+  mcrdlm5p1_ca_w_1_600_s_1_600=1.11e-05 mcrdlm5p1_cc_w_1_600_s_1_600=6.07e-11 mcrdlm5p1_cf_w_1_600_s_1_600=8.87e-12
+  mcrdlm5p1_ca_w_1_600_s_1_700=1.11e-05 mcrdlm5p1_cc_w_1_600_s_1_700=5.76e-11 mcrdlm5p1_cf_w_1_600_s_1_700=9.37e-12
+  mcrdlm5p1_ca_w_1_600_s_1_900=1.11e-05 mcrdlm5p1_cc_w_1_600_s_1_900=5.21e-11 mcrdlm5p1_cf_w_1_600_s_1_900=1.03e-11
+  mcrdlm5p1_ca_w_1_600_s_2_000=1.11e-05 mcrdlm5p1_cc_w_1_600_s_2_000=4.99e-11 mcrdlm5p1_cf_w_1_600_s_2_000=1.08e-11
+  mcrdlm5p1_ca_w_1_600_s_2_400=1.11e-05 mcrdlm5p1_cc_w_1_600_s_2_400=4.20e-11 mcrdlm5p1_cf_w_1_600_s_2_400=1.27e-11
+  mcrdlm5p1_ca_w_1_600_s_2_800=1.11e-05 mcrdlm5p1_cc_w_1_600_s_2_800=3.62e-11 mcrdlm5p1_cf_w_1_600_s_2_800=1.45e-11
+  mcrdlm5p1_ca_w_1_600_s_3_200=1.11e-05 mcrdlm5p1_cc_w_1_600_s_3_200=3.15e-11 mcrdlm5p1_cf_w_1_600_s_3_200=1.62e-11
+  mcrdlm5p1_ca_w_1_600_s_4_800=1.11e-05 mcrdlm5p1_cc_w_1_600_s_4_800=1.95e-11 mcrdlm5p1_cf_w_1_600_s_4_800=2.20e-11
+  mcrdlm5p1_ca_w_1_600_s_10_000=1.11e-05 mcrdlm5p1_cc_w_1_600_s_10_000=5.02e-12 mcrdlm5p1_cf_w_1_600_s_10_000=3.24e-11
+  mcrdlm5p1_ca_w_1_600_s_12_000=1.11e-05 mcrdlm5p1_cc_w_1_600_s_12_000=3.05e-12 mcrdlm5p1_cf_w_1_600_s_12_000=3.42e-11
+  mcrdlm5p1_ca_w_4_000_s_1_600=1.11e-05 mcrdlm5p1_cc_w_4_000_s_1_600=6.43e-11 mcrdlm5p1_cf_w_4_000_s_1_600=8.86e-12
+  mcrdlm5p1_ca_w_4_000_s_1_700=1.11e-05 mcrdlm5p1_cc_w_4_000_s_1_700=6.09e-11 mcrdlm5p1_cf_w_4_000_s_1_700=9.34e-12
+  mcrdlm5p1_ca_w_4_000_s_1_900=1.11e-05 mcrdlm5p1_cc_w_4_000_s_1_900=5.53e-11 mcrdlm5p1_cf_w_4_000_s_1_900=1.03e-11
+  mcrdlm5p1_ca_w_4_000_s_2_000=1.11e-05 mcrdlm5p1_cc_w_4_000_s_2_000=5.28e-11 mcrdlm5p1_cf_w_4_000_s_2_000=1.08e-11
+  mcrdlm5p1_ca_w_4_000_s_2_400=1.11e-05 mcrdlm5p1_cc_w_4_000_s_2_400=4.46e-11 mcrdlm5p1_cf_w_4_000_s_2_400=1.27e-11
+  mcrdlm5p1_ca_w_4_000_s_2_800=1.11e-05 mcrdlm5p1_cc_w_4_000_s_2_800=3.84e-11 mcrdlm5p1_cf_w_4_000_s_2_800=1.45e-11
+  mcrdlm5p1_ca_w_4_000_s_3_200=1.11e-05 mcrdlm5p1_cc_w_4_000_s_3_200=3.34e-11 mcrdlm5p1_cf_w_4_000_s_3_200=1.62e-11
+  mcrdlm5p1_ca_w_4_000_s_4_800=1.11e-05 mcrdlm5p1_cc_w_4_000_s_4_800=2.07e-11 mcrdlm5p1_cf_w_4_000_s_4_800=2.22e-11
+  mcrdlm5p1_ca_w_4_000_s_10_000=1.11e-05 mcrdlm5p1_cc_w_4_000_s_10_000=5.40e-12 mcrdlm5p1_cf_w_4_000_s_10_000=3.32e-11
+  mcrdlm5p1_ca_w_4_000_s_12_000=1.11e-05 mcrdlm5p1_cc_w_4_000_s_12_000=3.30e-12 mcrdlm5p1_cf_w_4_000_s_12_000=3.51e-11
+  mcrdlm5l1_ca_w_1_600_s_1_600=1.19e-05 mcrdlm5l1_cc_w_1_600_s_1_600=6.01e-11 mcrdlm5l1_cf_w_1_600_s_1_600=9.45e-12
+  mcrdlm5l1_ca_w_1_600_s_1_700=1.19e-05 mcrdlm5l1_cc_w_1_600_s_1_700=5.68e-11 mcrdlm5l1_cf_w_1_600_s_1_700=9.99e-12
+  mcrdlm5l1_ca_w_1_600_s_1_900=1.19e-05 mcrdlm5l1_cc_w_1_600_s_1_900=5.13e-11 mcrdlm5l1_cf_w_1_600_s_1_900=1.10e-11
+  mcrdlm5l1_ca_w_1_600_s_2_000=1.19e-05 mcrdlm5l1_cc_w_1_600_s_2_000=4.90e-11 mcrdlm5l1_cf_w_1_600_s_2_000=1.15e-11
+  mcrdlm5l1_ca_w_1_600_s_2_400=1.19e-05 mcrdlm5l1_cc_w_1_600_s_2_400=4.11e-11 mcrdlm5l1_cf_w_1_600_s_2_400=1.35e-11
+  mcrdlm5l1_ca_w_1_600_s_2_800=1.19e-05 mcrdlm5l1_cc_w_1_600_s_2_800=3.53e-11 mcrdlm5l1_cf_w_1_600_s_2_800=1.54e-11
+  mcrdlm5l1_ca_w_1_600_s_3_200=1.19e-05 mcrdlm5l1_cc_w_1_600_s_3_200=3.06e-11 mcrdlm5l1_cf_w_1_600_s_3_200=1.72e-11
+  mcrdlm5l1_ca_w_1_600_s_4_800=1.19e-05 mcrdlm5l1_cc_w_1_600_s_4_800=1.86e-11 mcrdlm5l1_cf_w_1_600_s_4_800=2.32e-11
+  mcrdlm5l1_ca_w_1_600_s_10_000=1.19e-05 mcrdlm5l1_cc_w_1_600_s_10_000=4.49e-12 mcrdlm5l1_cf_w_1_600_s_10_000=3.36e-11
+  mcrdlm5l1_ca_w_1_600_s_12_000=1.19e-05 mcrdlm5l1_cc_w_1_600_s_12_000=2.65e-12 mcrdlm5l1_cf_w_1_600_s_12_000=3.53e-11
+  mcrdlm5l1_ca_w_4_000_s_1_600=1.19e-05 mcrdlm5l1_cc_w_4_000_s_1_600=6.32e-11 mcrdlm5l1_cf_w_4_000_s_1_600=9.45e-12
+  mcrdlm5l1_ca_w_4_000_s_1_700=1.19e-05 mcrdlm5l1_cc_w_4_000_s_1_700=5.98e-11 mcrdlm5l1_cf_w_4_000_s_1_700=9.98e-12
+  mcrdlm5l1_ca_w_4_000_s_1_900=1.19e-05 mcrdlm5l1_cc_w_4_000_s_1_900=5.42e-11 mcrdlm5l1_cf_w_4_000_s_1_900=1.10e-11
+  mcrdlm5l1_ca_w_4_000_s_2_000=1.19e-05 mcrdlm5l1_cc_w_4_000_s_2_000=5.16e-11 mcrdlm5l1_cf_w_4_000_s_2_000=1.15e-11
+  mcrdlm5l1_ca_w_4_000_s_2_400=1.19e-05 mcrdlm5l1_cc_w_4_000_s_2_400=4.34e-11 mcrdlm5l1_cf_w_4_000_s_2_400=1.35e-11
+  mcrdlm5l1_ca_w_4_000_s_2_800=1.19e-05 mcrdlm5l1_cc_w_4_000_s_2_800=3.73e-11 mcrdlm5l1_cf_w_4_000_s_2_800=1.54e-11
+  mcrdlm5l1_ca_w_4_000_s_3_200=1.19e-05 mcrdlm5l1_cc_w_4_000_s_3_200=3.23e-11 mcrdlm5l1_cf_w_4_000_s_3_200=1.72e-11
+  mcrdlm5l1_ca_w_4_000_s_4_800=1.19e-05 mcrdlm5l1_cc_w_4_000_s_4_800=1.96e-11 mcrdlm5l1_cf_w_4_000_s_4_800=2.35e-11
+  mcrdlm5l1_ca_w_4_000_s_10_000=1.19e-05 mcrdlm5l1_cc_w_4_000_s_10_000=4.82e-12 mcrdlm5l1_cf_w_4_000_s_10_000=3.44e-11
+  mcrdlm5l1_ca_w_4_000_s_12_000=1.19e-05 mcrdlm5l1_cc_w_4_000_s_12_000=2.83e-12 mcrdlm5l1_cf_w_4_000_s_12_000=3.62e-11
+  mcrdlm5m1_ca_w_1_600_s_1_600=1.32e-05 mcrdlm5m1_cc_w_1_600_s_1_600=5.88e-11 mcrdlm5m1_cf_w_1_600_s_1_600=1.05e-11
+  mcrdlm5m1_ca_w_1_600_s_1_700=1.32e-05 mcrdlm5m1_cc_w_1_600_s_1_700=5.54e-11 mcrdlm5m1_cf_w_1_600_s_1_700=1.10e-11
+  mcrdlm5m1_ca_w_1_600_s_1_900=1.32e-05 mcrdlm5m1_cc_w_1_600_s_1_900=4.99e-11 mcrdlm5m1_cf_w_1_600_s_1_900=1.22e-11
+  mcrdlm5m1_ca_w_1_600_s_2_000=1.32e-05 mcrdlm5m1_cc_w_1_600_s_2_000=4.76e-11 mcrdlm5m1_cf_w_1_600_s_2_000=1.27e-11
+  mcrdlm5m1_ca_w_1_600_s_2_400=1.32e-05 mcrdlm5m1_cc_w_1_600_s_2_400=3.97e-11 mcrdlm5m1_cf_w_1_600_s_2_400=1.49e-11
+  mcrdlm5m1_ca_w_1_600_s_2_800=1.32e-05 mcrdlm5m1_cc_w_1_600_s_2_800=3.39e-11 mcrdlm5m1_cf_w_1_600_s_2_800=1.69e-11
+  mcrdlm5m1_ca_w_1_600_s_3_200=1.32e-05 mcrdlm5m1_cc_w_1_600_s_3_200=2.91e-11 mcrdlm5m1_cf_w_1_600_s_3_200=1.88e-11
+  mcrdlm5m1_ca_w_1_600_s_4_800=1.32e-05 mcrdlm5m1_cc_w_1_600_s_4_800=1.71e-11 mcrdlm5m1_cf_w_1_600_s_4_800=2.52e-11
+  mcrdlm5m1_ca_w_1_600_s_10_000=1.32e-05 mcrdlm5m1_cc_w_1_600_s_10_000=3.76e-12 mcrdlm5m1_cf_w_1_600_s_10_000=3.56e-11
+  mcrdlm5m1_ca_w_1_600_s_12_000=1.32e-05 mcrdlm5m1_cc_w_1_600_s_12_000=2.13e-12 mcrdlm5m1_cf_w_1_600_s_12_000=3.71e-11
+  mcrdlm5m1_ca_w_4_000_s_1_600=1.32e-05 mcrdlm5m1_cc_w_4_000_s_1_600=6.15e-11 mcrdlm5m1_cf_w_4_000_s_1_600=1.05e-11
+  mcrdlm5m1_ca_w_4_000_s_1_700=1.32e-05 mcrdlm5m1_cc_w_4_000_s_1_700=5.82e-11 mcrdlm5m1_cf_w_4_000_s_1_700=1.10e-11
+  mcrdlm5m1_ca_w_4_000_s_1_900=1.32e-05 mcrdlm5m1_cc_w_4_000_s_1_900=5.24e-11 mcrdlm5m1_cf_w_4_000_s_1_900=1.22e-11
+  mcrdlm5m1_ca_w_4_000_s_2_000=1.32e-05 mcrdlm5m1_cc_w_4_000_s_2_000=5.00e-11 mcrdlm5m1_cf_w_4_000_s_2_000=1.27e-11
+  mcrdlm5m1_ca_w_4_000_s_2_400=1.32e-05 mcrdlm5m1_cc_w_4_000_s_2_400=4.18e-11 mcrdlm5m1_cf_w_4_000_s_2_400=1.49e-11
+  mcrdlm5m1_ca_w_4_000_s_2_800=1.32e-05 mcrdlm5m1_cc_w_4_000_s_2_800=3.55e-11 mcrdlm5m1_cf_w_4_000_s_2_800=1.70e-11
+  mcrdlm5m1_ca_w_4_000_s_3_200=1.32e-05 mcrdlm5m1_cc_w_4_000_s_3_200=3.06e-11 mcrdlm5m1_cf_w_4_000_s_3_200=1.89e-11
+  mcrdlm5m1_ca_w_4_000_s_4_800=1.32e-05 mcrdlm5m1_cc_w_4_000_s_4_800=1.81e-11 mcrdlm5m1_cf_w_4_000_s_4_800=2.55e-11
+  mcrdlm5m1_ca_w_4_000_s_10_000=1.32e-05 mcrdlm5m1_cc_w_4_000_s_10_000=3.99e-12 mcrdlm5m1_cf_w_4_000_s_10_000=3.62e-11
+  mcrdlm5m1_ca_w_4_000_s_12_000=1.32e-05 mcrdlm5m1_cc_w_4_000_s_12_000=2.28e-12 mcrdlm5m1_cf_w_4_000_s_12_000=3.79e-11
+  mcrdlm5m2_ca_w_1_600_s_1_600=1.51e-05 mcrdlm5m2_cc_w_1_600_s_1_600=5.70e-11 mcrdlm5m2_cf_w_1_600_s_1_600=1.18e-11
+  mcrdlm5m2_ca_w_1_600_s_1_700=1.51e-05 mcrdlm5m2_cc_w_1_600_s_1_700=5.37e-11 mcrdlm5m2_cf_w_1_600_s_1_700=1.25e-11
+  mcrdlm5m2_ca_w_1_600_s_1_900=1.51e-05 mcrdlm5m2_cc_w_1_600_s_1_900=4.82e-11 mcrdlm5m2_cf_w_1_600_s_1_900=1.38e-11
+  mcrdlm5m2_ca_w_1_600_s_2_000=1.51e-05 mcrdlm5m2_cc_w_1_600_s_2_000=4.59e-11 mcrdlm5m2_cf_w_1_600_s_2_000=1.44e-11
+  mcrdlm5m2_ca_w_1_600_s_2_400=1.51e-05 mcrdlm5m2_cc_w_1_600_s_2_400=3.81e-11 mcrdlm5m2_cf_w_1_600_s_2_400=1.68e-11
+  mcrdlm5m2_ca_w_1_600_s_2_800=1.51e-05 mcrdlm5m2_cc_w_1_600_s_2_800=3.21e-11 mcrdlm5m2_cf_w_1_600_s_2_800=1.90e-11
+  mcrdlm5m2_ca_w_1_600_s_3_200=1.51e-05 mcrdlm5m2_cc_w_1_600_s_3_200=2.74e-11 mcrdlm5m2_cf_w_1_600_s_3_200=2.11e-11
+  mcrdlm5m2_ca_w_1_600_s_4_800=1.51e-05 mcrdlm5m2_cc_w_1_600_s_4_800=1.55e-11 mcrdlm5m2_cf_w_1_600_s_4_800=2.79e-11
+  mcrdlm5m2_ca_w_1_600_s_10_000=1.51e-05 mcrdlm5m2_cc_w_1_600_s_10_000=3.02e-12 mcrdlm5m2_cf_w_1_600_s_10_000=3.79e-11
+  mcrdlm5m2_ca_w_1_600_s_12_000=1.51e-05 mcrdlm5m2_cc_w_1_600_s_12_000=1.65e-12 mcrdlm5m2_cf_w_1_600_s_12_000=3.92e-11
+  mcrdlm5m2_ca_w_4_000_s_1_600=1.51e-05 mcrdlm5m2_cc_w_4_000_s_1_600=5.95e-11 mcrdlm5m2_cf_w_4_000_s_1_600=1.18e-11
+  mcrdlm5m2_ca_w_4_000_s_1_700=1.51e-05 mcrdlm5m2_cc_w_4_000_s_1_700=5.62e-11 mcrdlm5m2_cf_w_4_000_s_1_700=1.25e-11
+  mcrdlm5m2_ca_w_4_000_s_1_900=1.51e-05 mcrdlm5m2_cc_w_4_000_s_1_900=5.04e-11 mcrdlm5m2_cf_w_4_000_s_1_900=1.38e-11
+  mcrdlm5m2_ca_w_4_000_s_2_000=1.51e-05 mcrdlm5m2_cc_w_4_000_s_2_000=4.79e-11 mcrdlm5m2_cf_w_4_000_s_2_000=1.44e-11
+  mcrdlm5m2_ca_w_4_000_s_2_400=1.51e-05 mcrdlm5m2_cc_w_4_000_s_2_400=3.97e-11 mcrdlm5m2_cf_w_4_000_s_2_400=1.68e-11
+  mcrdlm5m2_ca_w_4_000_s_2_800=1.51e-05 mcrdlm5m2_cc_w_4_000_s_2_800=3.35e-11 mcrdlm5m2_cf_w_4_000_s_2_800=1.91e-11
+  mcrdlm5m2_ca_w_4_000_s_3_200=1.51e-05 mcrdlm5m2_cc_w_4_000_s_3_200=2.87e-11 mcrdlm5m2_cf_w_4_000_s_3_200=2.12e-11
+  mcrdlm5m2_ca_w_4_000_s_4_800=1.51e-05 mcrdlm5m2_cc_w_4_000_s_4_800=1.64e-11 mcrdlm5m2_cf_w_4_000_s_4_800=2.81e-11
+  mcrdlm5m2_ca_w_4_000_s_10_000=1.51e-05 mcrdlm5m2_cc_w_4_000_s_10_000=3.22e-12 mcrdlm5m2_cf_w_4_000_s_10_000=3.86e-11
+  mcrdlm5m2_ca_w_4_000_s_12_000=1.51e-05 mcrdlm5m2_cc_w_4_000_s_12_000=1.72e-12 mcrdlm5m2_cf_w_4_000_s_12_000=4.00e-11
+  mcrdlm5m3_ca_w_1_600_s_1_600=2.21e-05 mcrdlm5m3_cc_w_1_600_s_1_600=5.20e-11 mcrdlm5m3_cf_w_1_600_s_1_600=1.68e-11
+  mcrdlm5m3_ca_w_1_600_s_1_700=2.21e-05 mcrdlm5m3_cc_w_1_600_s_1_700=4.87e-11 mcrdlm5m3_cf_w_1_600_s_1_700=1.76e-11
+  mcrdlm5m3_ca_w_1_600_s_1_900=2.21e-05 mcrdlm5m3_cc_w_1_600_s_1_900=4.32e-11 mcrdlm5m3_cf_w_1_600_s_1_900=1.93e-11
+  mcrdlm5m3_ca_w_1_600_s_2_000=2.21e-05 mcrdlm5m3_cc_w_1_600_s_2_000=4.09e-11 mcrdlm5m3_cf_w_1_600_s_2_000=2.01e-11
+  mcrdlm5m3_ca_w_1_600_s_2_400=2.21e-05 mcrdlm5m3_cc_w_1_600_s_2_400=3.31e-11 mcrdlm5m3_cf_w_1_600_s_2_400=2.32e-11
+  mcrdlm5m3_ca_w_1_600_s_2_800=2.21e-05 mcrdlm5m3_cc_w_1_600_s_2_800=2.72e-11 mcrdlm5m3_cf_w_1_600_s_2_800=2.60e-11
+  mcrdlm5m3_ca_w_1_600_s_3_200=2.21e-05 mcrdlm5m3_cc_w_1_600_s_3_200=2.26e-11 mcrdlm5m3_cf_w_1_600_s_3_200=2.85e-11
+  mcrdlm5m3_ca_w_1_600_s_4_800=2.21e-05 mcrdlm5m3_cc_w_1_600_s_4_800=1.16e-11 mcrdlm5m3_cf_w_1_600_s_4_800=3.61e-11
+  mcrdlm5m3_ca_w_1_600_s_10_000=2.21e-05 mcrdlm5m3_cc_w_1_600_s_10_000=1.67e-12 mcrdlm5m3_cf_w_1_600_s_10_000=4.47e-11
+  mcrdlm5m3_ca_w_1_600_s_12_000=2.21e-05 mcrdlm5m3_cc_w_1_600_s_12_000=8.20e-13 mcrdlm5m3_cf_w_1_600_s_12_000=4.55e-11
+  mcrdlm5m3_ca_w_4_000_s_1_600=2.21e-05 mcrdlm5m3_cc_w_4_000_s_1_600=5.40e-11 mcrdlm5m3_cf_w_4_000_s_1_600=1.68e-11
+  mcrdlm5m3_ca_w_4_000_s_1_700=2.21e-05 mcrdlm5m3_cc_w_4_000_s_1_700=5.07e-11 mcrdlm5m3_cf_w_4_000_s_1_700=1.76e-11
+  mcrdlm5m3_ca_w_4_000_s_1_900=2.21e-05 mcrdlm5m3_cc_w_4_000_s_1_900=4.49e-11 mcrdlm5m3_cf_w_4_000_s_1_900=1.93e-11
+  mcrdlm5m3_ca_w_4_000_s_2_000=2.21e-05 mcrdlm5m3_cc_w_4_000_s_2_000=4.25e-11 mcrdlm5m3_cf_w_4_000_s_2_000=2.01e-11
+  mcrdlm5m3_ca_w_4_000_s_2_400=2.21e-05 mcrdlm5m3_cc_w_4_000_s_2_400=3.44e-11 mcrdlm5m3_cf_w_4_000_s_2_400=2.33e-11
+  mcrdlm5m3_ca_w_4_000_s_2_800=2.21e-05 mcrdlm5m3_cc_w_4_000_s_2_800=2.84e-11 mcrdlm5m3_cf_w_4_000_s_2_800=2.61e-11
+  mcrdlm5m3_ca_w_4_000_s_3_200=2.21e-05 mcrdlm5m3_cc_w_4_000_s_3_200=2.37e-11 mcrdlm5m3_cf_w_4_000_s_3_200=2.86e-11
+  mcrdlm5m3_ca_w_4_000_s_4_800=2.21e-05 mcrdlm5m3_cc_w_4_000_s_4_800=1.23e-11 mcrdlm5m3_cf_w_4_000_s_4_800=3.63e-11
+  mcrdlm5m3_ca_w_4_000_s_10_000=2.21e-05 mcrdlm5m3_cc_w_4_000_s_10_000=1.79e-12 mcrdlm5m3_cf_w_4_000_s_10_000=4.54e-11
+  mcrdlm5m3_ca_w_4_000_s_12_000=2.21e-05 mcrdlm5m3_cc_w_4_000_s_12_000=9.05e-13 mcrdlm5m3_cf_w_4_000_s_12_000=4.63e-11
+  mcrdlm5m4_ca_w_1_600_s_1_600=5.76e-05 mcrdlm5m4_cc_w_1_600_s_1_600=4.07e-11 mcrdlm5m4_cf_w_1_600_s_1_600=3.61e-11
+  mcrdlm5m4_ca_w_1_600_s_1_700=5.76e-05 mcrdlm5m4_cc_w_1_600_s_1_700=3.76e-11 mcrdlm5m4_cf_w_1_600_s_1_700=3.75e-11
+  mcrdlm5m4_ca_w_1_600_s_1_900=5.76e-05 mcrdlm5m4_cc_w_1_600_s_1_900=3.23e-11 mcrdlm5m4_cf_w_1_600_s_1_900=4.02e-11
+  mcrdlm5m4_ca_w_1_600_s_2_000=5.76e-05 mcrdlm5m4_cc_w_1_600_s_2_000=3.01e-11 mcrdlm5m4_cf_w_1_600_s_2_000=4.14e-11
+  mcrdlm5m4_ca_w_1_600_s_2_400=5.76e-05 mcrdlm5m4_cc_w_1_600_s_2_400=2.30e-11 mcrdlm5m4_cf_w_1_600_s_2_400=4.57e-11
+  mcrdlm5m4_ca_w_1_600_s_2_800=5.76e-05 mcrdlm5m4_cc_w_1_600_s_2_800=1.79e-11 mcrdlm5m4_cf_w_1_600_s_2_800=4.93e-11
+  mcrdlm5m4_ca_w_1_600_s_3_200=5.76e-05 mcrdlm5m4_cc_w_1_600_s_3_200=1.42e-11 mcrdlm5m4_cf_w_1_600_s_3_200=5.21e-11
+  mcrdlm5m4_ca_w_1_600_s_4_800=5.76e-05 mcrdlm5m4_cc_w_1_600_s_4_800=6.02e-12 mcrdlm5m4_cf_w_1_600_s_4_800=5.89e-11
+  mcrdlm5m4_ca_w_1_600_s_10_000=5.76e-05 mcrdlm5m4_cc_w_1_600_s_10_000=6.15e-13 mcrdlm5m4_cf_w_1_600_s_10_000=6.41e-11
+  mcrdlm5m4_ca_w_1_600_s_12_000=5.76e-05 mcrdlm5m4_cc_w_1_600_s_12_000=3.05e-13 mcrdlm5m4_cf_w_1_600_s_12_000=6.44e-11
+  mcrdlm5m4_ca_w_4_000_s_1_600=5.76e-05 mcrdlm5m4_cc_w_4_000_s_1_600=4.25e-11 mcrdlm5m4_cf_w_4_000_s_1_600=3.61e-11
+  mcrdlm5m4_ca_w_4_000_s_1_700=5.76e-05 mcrdlm5m4_cc_w_4_000_s_1_700=3.94e-11 mcrdlm5m4_cf_w_4_000_s_1_700=3.75e-11
+  mcrdlm5m4_ca_w_4_000_s_1_900=5.76e-05 mcrdlm5m4_cc_w_4_000_s_1_900=3.40e-11 mcrdlm5m4_cf_w_4_000_s_1_900=4.02e-11
+  mcrdlm5m4_ca_w_4_000_s_2_000=5.76e-05 mcrdlm5m4_cc_w_4_000_s_2_000=3.16e-11 mcrdlm5m4_cf_w_4_000_s_2_000=4.14e-11
+  mcrdlm5m4_ca_w_4_000_s_2_400=5.76e-05 mcrdlm5m4_cc_w_4_000_s_2_400=2.43e-11 mcrdlm5m4_cf_w_4_000_s_2_400=4.58e-11
+  mcrdlm5m4_ca_w_4_000_s_2_800=5.76e-05 mcrdlm5m4_cc_w_4_000_s_2_800=1.91e-11 mcrdlm5m4_cf_w_4_000_s_2_800=4.93e-11
+  mcrdlm5m4_ca_w_4_000_s_3_200=5.76e-05 mcrdlm5m4_cc_w_4_000_s_3_200=1.52e-11 mcrdlm5m4_cf_w_4_000_s_3_200=5.22e-11
+  mcrdlm5m4_ca_w_4_000_s_4_800=5.76e-05 mcrdlm5m4_cc_w_4_000_s_4_800=6.66e-12 mcrdlm5m4_cf_w_4_000_s_4_800=5.93e-11
+  mcrdlm5m4_ca_w_4_000_s_10_000=5.76e-05 mcrdlm5m4_cc_w_4_000_s_10_000=7.25e-13 mcrdlm5m4_cf_w_4_000_s_10_000=6.50e-11
+  mcrdlm5m4_ca_w_4_000_s_12_000=5.76e-05 mcrdlm5m4_cc_w_4_000_s_12_000=3.55e-13 mcrdlm5m4_cf_w_4_000_s_12_000=6.54e-11
+  cp1f=8.67e-05 cp1fsw=7.73e-11
+  cl1f=3.12e-05 cl1fsw=7.23e-11
+  cl1d=4.77e-05 cl1dsw=7.16e-11
+  cl1p1=7.09e-05 cl1p1sw=7.10e-11
+  cm1f=2.17e-05 cm1fsw=9.36e-11
+  cm1d=2.86e-05 cm1dsw=9.34e-11
+  cm1p1=3.55e-05 cm1p1sw=9.31e-11
+  cm1l1=8.73e-05 cm1l1sw=9.20e-11
+  cm2f=1.49e-05 cm2fsw=9.39e-11
+  cm2d=1.79e-05 cm2dsw=9.38e-11
+  cm2p1=2.04e-05 cm2p1sw=9.37e-11
+  cm2l1=3.10e-05 cm2l1sw=9.35e-11
+  cm2m1=9.04e-05 cm2m1sw=9.20e-11
+  cm3f=1.08e-05 cm3fsw=9.74e-11
+  cm3d=1.23e-05 cm3dsw=9.72e-11
+  cm3p1=1.35e-05 cm3p1sw=9.72e-11
+  cm3l1=1.74e-05 cm3l1sw=9.68e-11
+  cm3m1=2.75e-05 cm3m1sw=9.60e-11
+  cm3m2=6.49e-05 cm3m2sw=9.45e-11
+  cm4f=7.66e-06 cm4fsw=9.80e-11
+  cm4d=8.37e-06 cm4dsw=9.80e-11
+  cm4p1=8.88e-06 cm4p1sw=9.78e-11
+  cm4l1=1.04e-05 cm4l1sw=9.77e-11
+  cm4m1=1.34e-05 cm4m1sw=9.74e-11
+  cm4m2=1.86e-05 cm4m2sw=9.69e-11
+  cm4m3=6.43e-05 cm4m3sw=9.50e-11
+  cm5f=5.81e-06 cm5fsw=7.20e-11
+  cm5d=6.21e-06 cm5dsw=7.19e-11
+  cm5p1=6.49e-06 cm5p1sw=7.18e-11
+  cm5l1=7.27e-06 cm5l1sw=7.15e-11
+  cm5m1=8.59e-06 cm5m1sw=7.12e-11
+  cm5m2=1.05e-05 cm5m2sw=7.09e-11
+  cm5m3=1.75e-05 cm5m3sw=7.09e-11
+  cm5m4=5.30e-05 cm5m4sw=7.88e-11
+  crdlf=2.26e-06 crdlfsw=4.99e-11
+  crdld=2.32e-06 crdldsw=4.98e-11
+  crdlp1=2.36e-06 crdlp1sw=4.98e-11
+  crdll1=2.45e-06 crdll1sw=4.97e-11
+  crdlm1=2.58e-06 crdlm1sw=4.95e-11
+  crdlm2=2.73e-06 crdlm2sw=4.94e-11
+  crdlm3=3.06e-06 crdlm3sw=4.92e-11
+  crdlm4=3.47e-06 crdlm4sw=4.91e-11
+  crdlm5=4.58e-06 crdlm5sw=4.93e-11
+  cl1p1f=1.58e-04 cl1p1fsw=7.50e-11
+  cm1p1f=1.22e-04 cm1p1fsw=7.61e-11
+  cm2p1f=1.07e-04 cm2p1fsw=7.67e-11
+  cm3p1f=1.00e-04 cm3p1fsw=7.70e-11
+  cm4p1f=9.56e-05 cm4p1fsw=7.72e-11
+  cm5p1f=9.32e-05 cm5p1fsw=7.72e-11
+  crdlp1f=8.90e-05 crdlp1fsw=7.73e-11
+  cm1l1f=1.19e-04 cm1l1fsw=6.95e-11
+  cm1l1d=1.35e-04 cm1l1dsw=6.88e-11
+  cm1l1p1=1.59e-04 cm1l1p1sw=6.81e-11
+  cm2l1f=6.22e-05 cm2l1fsw=7.12e-11
+  cm2l1d=7.87e-05 cm2l1dsw=7.04e-11
+  cm2l1p1=1.02e-04 cm2l1p1sw=6.97e-11
+  cm3l1f=4.86e-05 cm3l1fsw=7.18e-11
+  cm3l1d=6.51e-05 cm3l1dsw=7.10e-11
+  cm3l1p1=8.83e-05 cm3l1p1sw=7.05e-11
+  cm4l1f=4.16e-05 cm4l1fsw=7.21e-11
+  cm4l1d=5.81e-05 cm4l1dsw=7.13e-11
+  cm4l1p1=8.13e-05 cm4l1p1sw=7.07e-11
+  cm5l1f=3.85e-05 cm5l1fsw=7.22e-11
+  cm5l1d=5.50e-05 cm5l1dsw=7.14e-11
+  cm5l1p1=7.81e-05 cm5l1p1sw=7.08e-11
+  crdll1f=3.36e-05 crdll1fsw=7.22e-11
+  crdll1d=5.02e-05 crdll1dsw=7.16e-11
+  crdll1p1=7.33e-05 crdll1p1sw=7.10e-11
+  cm2m1f=1.12e-04 cm2m1fsw=9.09e-11
+  cm2m1d=1.19e-04 cm2m1dsw=9.10e-11
+  cm2m1p1=1.26e-04 cm2m1p1sw=9.07e-11
+  cm2m1l1=1.78e-04 cm2m1l1sw=8.90e-11
+  cm3m1f=4.93e-05 cm3m1fsw=9.27e-11
+  cm3m1d=5.62e-05 cm3m1dsw=9.25e-11
+  cm3m1p1=6.31e-05 cm3m1p1sw=9.23e-11
+  cm3m1l1=1.15e-04 cm3m1l1sw=9.02e-11
+  cm4m1f=3.51e-05 cm4m1fsw=9.35e-11
+  cm4m1d=4.20e-05 cm4m1dsw=9.33e-11
+  cm4m1p1=4.90e-05 cm4m1p1sw=9.31e-11
+  cm4m1l1=1.01e-04 cm4m1l1sw=9.13e-11
+  cm5m1f=3.03e-05 cm5m1fsw=9.38e-11
+  cm5m1d=3.72e-05 cm5m1dsw=9.35e-11
+  cm5m1p1=4.42e-05 cm5m1p1sw=9.32e-11
+  cm5m1l1=9.59e-05 cm5m1l1sw=9.16e-11
+  crdlm1f=2.43e-05 crdlm1fsw=9.40e-11
+  crdlm1d=3.12e-05 crdlm1dsw=9.37e-11
+  crdlm1p1=3.81e-05 crdlm1p1sw=9.34e-11
+  crdlm1l1=8.99e-05 crdlm1l1sw=9.19e-11
+  cm3m2f=7.98e-05 cm3m2fsw=9.15e-11
+  cm3m2d=8.28e-05 cm3m2dsw=9.18e-11
+  cm3m2p1=8.53e-05 cm3m2p1sw=9.13e-11
+  cm3m2l1=9.58e-05 cm3m2l1sw=9.16e-11
+  cm3m2m1=1.55e-04 cm3m2m1sw=8.94e-11
+  cm4m2f=3.35e-05 cm4m2fsw=9.35e-11
+  cm4m2d=3.65e-05 cm4m2dsw=9.33e-11
+  cm4m2p1=3.90e-05 cm4m2p1sw=9.32e-11
+  cm4m2l1=4.95e-05 cm4m2l1sw=9.29e-11
+  cm4m2m1=1.09e-04 cm4m2m1sw=9.06e-11
+  cm5m2f=2.54e-05 cm5m2fsw=9.39e-11
+  cm5m2d=2.84e-05 cm5m2dsw=9.38e-11
+  cm5m2p1=3.09e-05 cm5m2p1sw=9.37e-11
+  cm5m2l1=4.14e-05 cm5m2l1sw=9.33e-11
+  cm5m2m1=1.01e-04 cm5m2m1sw=9.11e-11
+  crdlm2f=1.77e-05 crdlm2fsw=9.42e-11
+  crdlm2d=2.07e-05 crdlm2dsw=9.41e-11
+  crdlm2p1=2.32e-05 crdlm2p1sw=9.39e-11
+  crdlm2l1=3.37e-05 crdlm2l1sw=9.36e-11
+  crdlm2m1=9.32e-05 crdlm2m1sw=9.17e-11
+  cm4m3f=7.52e-05 cm4m3fsw=9.40e-11
+  cm4m3d=7.67e-05 cm4m3dsw=9.38e-11
+  cm4m3p1=7.78e-05 cm4m3p1sw=9.37e-11
+  cm4m3l1=8.17e-05 cm4m3l1sw=9.30e-11
+  cm4m3m1=9.19e-05 cm4m3m1sw=9.26e-11
+  cm4m3m2=1.29e-04 cm4m3m2sw=9.12e-11
+  cm5m3f=2.83e-05 cm5m3fsw=9.57e-11
+  cm5m3d=2.98e-05 cm5m3dsw=9.56e-11
+  cm5m3p1=3.10e-05 cm5m3p1sw=9.55e-11
+  cm5m3l1=3.48e-05 cm5m3l1sw=9.52e-11
+  cm5m3m1=4.50e-05 cm5m3m1sw=9.44e-11
+  cm5m3m2=8.23e-05 cm5m3m2sw=9.31e-11
+  crdlm3f=1.39e-05 crdlm3fsw=9.72e-11
+  crdlm3d=1.54e-05 crdlm3dsw=9.72e-11
+  crdlm3p1=1.65e-05 crdlm3p1sw=9.71e-11
+  crdlm3l1=2.04e-05 crdlm3l1sw=9.67e-11
+  crdlm3m1=3.06e-05 crdlm3m1sw=9.60e-11
+  crdlm3m2=6.79e-05 crdlm3m2sw=9.48e-11
+  cm5m4f=6.06e-05 cm5m4fsw=9.42e-11
+  cm5m4d=6.13e-05 cm5m4dsw=9.42e-11
+  cm5m4p1=6.19e-05 cm5m4p1sw=9.41e-11
+  cm5m4l1=6.34e-05 cm5m4l1sw=9.40e-11
+  cm5m4m1=6.64e-05 cm5m4m1sw=9.37e-11
+  cm5m4m2=7.15e-05 cm5m4m2sw=9.33e-11
+  cm5m4m3=1.17e-04 cm5m4m3sw=9.14e-11
+  crdlm4f=1.11e-05 crdlm4fsw=9.77e-11
+  crdlm4d=1.18e-05 crdlm4dsw=9.76e-11
+  crdlm4p1=1.23e-05 crdlm4p1sw=9.76e-11
+  crdlm4l1=1.39e-05 crdlm4l1sw=9.75e-11
+  crdlm4m1=1.68e-05 crdlm4m1sw=9.72e-11
+  crdlm4m2=2.20e-05 crdlm4m2sw=9.68e-11
+  crdlm4m3=6.78e-05 crdlm4m3sw=9.49e-11
+  crdlm5f=1.04e-05 crdlm5fsw=6.99e-11
+  crdlm5d=1.08e-05 crdlm5dsw=6.97e-11
+  crdlm5p1=1.11e-05 crdlm5p1sw=6.96e-11
+  crdlm5l1=1.19e-05 crdlm5l1sw=6.95e-11
+  crdlm5m1=1.32e-05 crdlm5m1sw=6.92e-11
+  crdlm5m2=1.51e-05 crdlm5m2sw=6.88e-11
+  crdlm5m3=2.21e-05 crdlm5m3sw=6.87e-11
+  crdlm5m4=5.76e-05 crdlm5m4sw=7.67e-11
