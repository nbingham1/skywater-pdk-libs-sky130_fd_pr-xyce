* SKY130 Spice File.
* Number of bins: 1
* 9 parameters
.param
+  sky130_fd_bs_flash__special_sonosfet_original__tox_mult=1.0
+  sky130_fd_bs_flash__special_sonosfet_original__ajunction_mult=1.0
+  sky130_fd_bs_flash__special_sonosfet_original__pjunction_mult=1.0
+  sky130_fd_bs_flash__special_sonosfet_original__overlap_mult=1.0
+  sky130_fd_bs_flash__special_sonosfet_original__lint_diff=0.0
+  sky130_fd_bs_flash__special_sonosfet_original__wint_diff=0.0
+  sky130_fd_bs_flash__special_sonosfet_original__dlc_diff=0.0
+  sky130_fd_bs_flash__special_sonosfet_original__dwc_diff=0.0
*
* sky130_fd_bs_flash__special_sonosfet_original, Bin 000, W = 0.45, L = 0.22
* ------------------------------------
+  sky130_fd_bs_flash__special_sonosfet_original__rdsw_diff_0=0.0
+  sky130_fd_bs_flash__special_sonosfet_original__vth0_diff_0=-2.1028
+  sky130_fd_bs_flash__special_sonosfet_original__u0_diff_0=6.2558e-4
+  sky130_fd_bs_flash__special_sonosfet_original__vsat_diff_0=0.0
+  sky130_fd_bs_flash__special_sonosfet_original__voff_diff_0=0.0
+  sky130_fd_bs_flash__special_sonosfet_original__k2_diff_0=0.0
+  sky130_fd_bs_flash__special_sonosfet_original__nfactor_diff_0=0.0
+  sky130_fd_bs_flash__special_sonosfet_original__kt1_diff_0=-3.2289e-1
