* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 8
.param
+  sky130_fd_pr__esd_pfet_g5v0d10v5__toxe_mult=1.042
+  sky130_fd_pr__esd_pfet_g5v0d10v5__rshp_mult=1.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__overlap_mult=1.1981e+0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__ajunction_mult=1.0559e+0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__pjunction_mult=1.0542e+0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__lint_diff=-1.21275e-8
+  sky130_fd_pr__esd_pfet_g5v0d10v5__wint_diff=2.252e-8
+  sky130_fd_pr__esd_pfet_g5v0d10v5__dlc_diff=-1.21275e-8
+  sky130_fd_pr__esd_pfet_g5v0d10v5__dwc_diff=2.252e-8
*
* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 000, W = 14.5, L = 0.55
* -----------------------------------
+  sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_0=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_0=0.0066792
+  sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_0=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_0=0.0055732
+  sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_0=57405.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_0=-0.039836
+  sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_0=-0.84048
+  sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_0=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_0=1.8175e-9
+  sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_0=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_0=-4.3477e-19
+  sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_0=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_0=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_0=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_0=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_0=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_0=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_0=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_0=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_0=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_0=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_0=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_0=-0.032489
*
* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 001, W = 15.5, L = 0.55
* -----------------------------------
+  sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_1=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_1=0.11937
+  sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_1=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_1=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_1=0.013842
+  sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_1=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_1=-0.0048548
+  sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_1=11004.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_1=0.050578
+  sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_1=9.3332e-11
+  sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_1=0.59173
+  sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_1=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_1=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_1=-2.2152e-18
+  sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_1=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_1=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_1=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_1=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_1=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_1=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_1=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_1=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_1=0.0
*
* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 002, W = 16.5, L = 0.55
* -----------------------------------
+  sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_2=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_2=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_2=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_2=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_2=5.2299e-2
+  sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_2=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_2=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_2=9.1344e-3
+  sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_2=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_2=-4.0166e-4
+  sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_2=-1.2687e-2
+  sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_2=2.4782e-11
+  sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_2=3.6143e+4
+  sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_2=4.0028e-1
+  sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_2=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_2=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_2=1.3690e-19
+  sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_2=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_2=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_2=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_2=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_2=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_2=0.0
*
* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 003, W = 17.5, L = 0.55
* -----------------------------------
+  sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_3=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_3=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_3=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_3=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_3=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_3=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_3=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_3=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_3=2.0000e-2
+  sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_3=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_3=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_3=6.1506e-3
+  sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_3=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_3=5.9152e-3
+  sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_3=-4.2250e-2
+  sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_3=1.8174e-9
+  sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_3=2.3364e+4
+  sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_3=4.0000e-6
+  sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_3=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_3=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_3=-5.2157e-19
+  sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_3=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_3=0.0
*
* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 004, W = 19.5, L = 0.55
* -----------------------------------
+  sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_4=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_4=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_4=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_4=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_4=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_4=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_4=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_4=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_4=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_4=-0.049006
+  sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_4=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_4=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_4=0.0067633
+  sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_4=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_4=0.0052948
+  sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_4=-0.042196
+  sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_4=1.782e-9
+  sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_4=47926.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_4=-1.0053
+  sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_4=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_4=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_4=-4.6278e-19
+  sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_4=0.0
*
* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 005, W = 21.5, L = 0.55
* -----------------------------------
+  sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_5=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_5=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_5=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_5=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_5=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_5=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_5=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_5=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_5=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_5=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_5=0.13767
+  sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_5=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_5=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_5=0.014733
+  sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_5=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_5=-0.0063472
+  sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_5=0.06743
+  sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_5=-2.5905e-12
+  sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_5=15839.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_5=0.62815
+  sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_5=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_5=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_5=-2.734e-18
*
* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 006, W = 23.5, L = 0.55
* -----------------------------------
+  sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_6=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_6=-2.9719e-18
+  sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_6=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_6=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_6=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_6=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_6=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_6=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_6=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_6=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_6=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_6=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_6=0.15175
+  sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_6=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_6=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_6=0.014735
+  sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_6=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_6=-0.0073782
+  sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_6=0.086313
+  sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_6=-6.8974e-11
+  sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_6=27158.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_6=0.57872
+  sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_6=0.0
*
* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 007, W = 26.5, L = 0.55
* -----------------------------------
+  sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_7=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_7=-1.8438e-18
+  sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_7=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_7=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_7=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_7=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_7=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_7=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_7=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_7=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_7=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_7=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_7=0.10854
+  sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_7=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_7=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_7=0.013897
+  sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_7=0.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_7=-0.0041489
+  sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_7=0.035699
+  sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_7=1.8882e-10
+  sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_7=12478.0
+  sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_7=0.60147
+  sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_7=0.0
.include "sky130_fd_pr__esd_pfet_g5v0d10v5.pm3.spice"
