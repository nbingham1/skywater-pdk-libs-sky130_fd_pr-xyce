* SKY130 Spice File.
* Number of bins: 1
* 9 parameters
.param
+  sky130_fd_bs_flash__special_sonosfet_star__tox_mult=1.0
+  sky130_fd_bs_flash__special_sonosfet_star__ajunction_mult=1.0
+  sky130_fd_bs_flash__special_sonosfet_star__pjunction_mult=1.0
+  sky130_fd_bs_flash__special_sonosfet_star__overlap_mult=1.0
+  sky130_fd_bs_flash__special_sonosfet_star__lint_diff=0.0
+  sky130_fd_bs_flash__special_sonosfet_star__wint_diff=0.0
+  sky130_fd_bs_flash__special_sonosfet_star__dlc_diff=0.0
+  sky130_fd_bs_flash__special_sonosfet_star__dwc_diff=0.0
*
* sky130_fd_bs_flash__special_sonosfet_star, Bin 000, W = 0.45, L = 0.22
* ------------------------------------
+  sky130_fd_bs_flash__special_sonosfet_star__k2_diff_0=0.0
+  sky130_fd_bs_flash__special_sonosfet_star__vth0_diff_0=5.0690e-1
+  sky130_fd_bs_flash__special_sonosfet_star__u0_diff_0=-2.1647e-3
+  sky130_fd_bs_flash__special_sonosfet_star__vsat_diff_0=0.0
+  sky130_fd_bs_flash__special_sonosfet_star__kt1_diff_0=-4.2963e-1
+  sky130_fd_bs_flash__special_sonosfet_star__nfactor_diff_0=0.0
+  sky130_fd_bs_flash__special_sonosfet_star__rdsw_diff_0=0.0
+  sky130_fd_bs_flash__special_sonosfet_star__voff_diff_0=0.0
*
* sky130_fd_bs_flash__special_sonosfet_star, Bin 001, W = 1.00, L = 0.50
* ------------------------------------
+  sky130_fd_bs_flash__special_sonosfet_star__k2_diff_1=0.0
+  sky130_fd_bs_flash__special_sonosfet_star__vth0_diff_1=1.3855
+  sky130_fd_bs_flash__special_sonosfet_star__vsat_diff_1=0.0
+  sky130_fd_bs_flash__special_sonosfet_star__kt1_diff_1=-3.2807e-1
+  sky130_fd_bs_flash__special_sonosfet_star__u0_diff_1=-5.0631e-3
+  sky130_fd_bs_flash__special_sonosfet_star__nfactor_diff_1=0.0
+  sky130_fd_bs_flash__special_sonosfet_star__rdsw_diff_1=0.0
+  sky130_fd_bs_flash__special_sonosfet_star__voff_diff_1=0.0
*
* sky130_fd_bs_flash__special_sonosfet_star, Bin 002, W = 0.35, L = 0.15
* ------------------------------------
+  sky130_fd_bs_flash__special_sonosfet_star__k2_diff_2=0.0
+  sky130_fd_bs_flash__special_sonosfet_star__vth0_diff_2=2.7494e-1
+  sky130_fd_bs_flash__special_sonosfet_star__u0_diff_2=-8.1788e-3
+  sky130_fd_bs_flash__special_sonosfet_star__vsat_diff_2=0.0
+  sky130_fd_bs_flash__special_sonosfet_star__kt1_diff_2=-6.7944e-1
+  sky130_fd_bs_flash__special_sonosfet_star__nfactor_diff_2=0.0
+  sky130_fd_bs_flash__special_sonosfet_star__rdsw_diff_2=0.0
+  sky130_fd_bs_flash__special_sonosfet_star__voff_diff_2=0.0
